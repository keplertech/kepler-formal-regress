module ibex_core (alert_major_o,
    alert_minor_o,
    clk_i,
    core_sleep_o,
    data_err_i,
    data_gnt_i,
    data_req_o,
    data_rvalid_i,
    data_we_o,
    debug_req_i,
    fetch_enable_i,
    instr_err_i,
    instr_gnt_i,
    instr_req_o,
    instr_rvalid_i,
    irq_external_i,
    irq_nm_i,
    irq_software_i,
    irq_timer_i,
    rst_ni,
    test_en_i,
    boot_addr_i,
    data_addr_o,
    data_be_o,
    data_rdata_i,
    data_wdata_o,
    hart_id_i,
    instr_addr_o,
    instr_rdata_i,
    irq_fast_i);
 output alert_major_o;
 output alert_minor_o;
 input clk_i;
 output core_sleep_o;
 input data_err_i;
 input data_gnt_i;
 output data_req_o;
 input data_rvalid_i;
 output data_we_o;
 input debug_req_i;
 input fetch_enable_i;
 input instr_err_i;
 input instr_gnt_i;
 output instr_req_o;
 input instr_rvalid_i;
 input irq_external_i;
 input irq_nm_i;
 input irq_software_i;
 input irq_timer_i;
 input rst_ni;
 input test_en_i;
 input [31:0] boot_addr_i;
 output [31:0] data_addr_o;
 output [3:0] data_be_o;
 input [31:0] data_rdata_i;
 output [31:0] data_wdata_o;
 input [31:0] hart_id_i;
 output [31:0] instr_addr_o;
 input [31:0] instr_rdata_i;
 input [14:0] irq_fast_i;

 wire net_8;
 wire net_7;
 wire net_6;
 wire net_5;
 wire net_4;
 wire net_3;
 wire net_2;
 wire net_1;
 wire net;
 wire \alu_adder_result_ex[0] ;
 wire \alu_adder_result_ex[1] ;
 wire net460;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net461;
 wire net462;
 wire _03652_;
 wire _03659_;
 wire _03665_;
 wire _03671_;
 wire _03677_;
 wire _03682_;
 wire _03687_;
 wire _03692_;
 wire _03697_;
 wire _03702_;
 wire _03707_;
 wire _03712_;
 wire _03717_;
 wire _03722_;
 wire _03727_;
 wire _03732_;
 wire _03737_;
 wire _03742_;
 wire _03747_;
 wire _03752_;
 wire _03757_;
 wire _03762_;
 wire _03767_;
 wire _03772_;
 wire _03777_;
 wire _03782_;
 wire _03787_;
 wire _03792_;
 wire _03798_;
 wire _03803_;
 wire _03808_;
 wire _03814_;
 wire _08254_;
 wire _09346_;
 wire _10414_;
 wire _11205_;
 wire _12286_;
 wire _13402_;
 wire _14300_;
 wire _15132_;
 wire _15569_;
 wire _02071_;
 wire _02146_;
 wire _02213_;
 wire _02289_;
 wire _02368_;
 wire _02445_;
 wire _02509_;
 wire _02555_;
 wire _02622_;
 wire _02687_;
 wire _02752_;
 wire _02824_;
 wire _02890_;
 wire _02957_;
 wire _03024_;
 wire _03091_;
 wire _03165_;
 wire _03230_;
 wire _03301_;
 wire _03373_;
 wire _03442_;
 wire _03511_;
 wire _03581_;
 wire _03632_;
 wire _00078_;
 wire _00089_;
 wire _00100_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00010_;
 wire _00021_;
 wire _00032_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00044_;
 wire _00055_;
 wire _00066_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _03895_;
 wire _06507_;
 wire _03960_;
 wire _04001_;
 wire _04076_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06519_;
 wire _06520_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06528_;
 wire _06530_;
 wire _06534_;
 wire _06537_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06545_;
 wire _06549_;
 wire _06551_;
 wire _06559_;
 wire _06562_;
 wire _03832_;
 wire _03844_;
 wire _03865_;
 wire _03896_;
 wire _03930_;
 wire _03961_;
 wire _04003_;
 wire _04077_;
 wire _04141_;
 wire _04211_;
 wire _04288_;
 wire _04364_;
 wire _04443_;
 wire _04524_;
 wire _04604_;
 wire _04705_;
 wire _04831_;
 wire _04949_;
 wire _05051_;
 wire _05172_;
 wire _05275_;
 wire _05417_;
 wire _05527_;
 wire _05631_;
 wire _05741_;
 wire _05861_;
 wire _05955_;
 wire _06064_;
 wire _06141_;
 wire _06234_;
 wire _06322_;
 wire _06407_;
 wire _06463_;
 wire _06506_;
 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04002_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06508_;
 wire _06512_;
 wire _06517_;
 wire _06518_;
 wire _06521_;
 wire _06522_;
 wire _06527_;
 wire _06529_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06535_;
 wire _06536_;
 wire _06538_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06550_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06560_;
 wire _06561_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire _10563_;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire _10582_;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire _10602_;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire _10609_;
 wire _10610_;
 wire _10611_;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire _10618_;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire _10632_;
 wire _10633_;
 wire _10634_;
 wire _10635_;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire _10652_;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire _10671_;
 wire _10672_;
 wire _10673_;
 wire _10674_;
 wire _10675_;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire _10689_;
 wire _10690_;
 wire _10691_;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10727_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire _10740_;
 wire _10741_;
 wire _10742_;
 wire _10743_;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10751_;
 wire _10752_;
 wire _10753_;
 wire _10754_;
 wire _10755_;
 wire _10756_;
 wire _10757_;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10771_;
 wire _10772_;
 wire _10773_;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire _10781_;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire _10785_;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire _10795_;
 wire _10796_;
 wire _10797_;
 wire _10798_;
 wire _10799_;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire _10807_;
 wire _10808_;
 wire _10809_;
 wire _10810_;
 wire _10811_;
 wire _10812_;
 wire _10813_;
 wire _10814_;
 wire _10815_;
 wire _10816_;
 wire _10817_;
 wire _10818_;
 wire _10819_;
 wire _10820_;
 wire _10821_;
 wire _10822_;
 wire _10823_;
 wire _10824_;
 wire _10825_;
 wire _10826_;
 wire _10827_;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire _10831_;
 wire _10832_;
 wire _10833_;
 wire _10834_;
 wire _10835_;
 wire _10836_;
 wire _10837_;
 wire _10838_;
 wire _10839_;
 wire _10840_;
 wire _10841_;
 wire _10842_;
 wire _10843_;
 wire _10844_;
 wire _10845_;
 wire _10846_;
 wire _10847_;
 wire _10848_;
 wire _10849_;
 wire _10850_;
 wire _10851_;
 wire _10852_;
 wire _10853_;
 wire _10854_;
 wire _10855_;
 wire _10856_;
 wire _10857_;
 wire _10858_;
 wire _10859_;
 wire _10860_;
 wire _10861_;
 wire _10862_;
 wire _10863_;
 wire _10864_;
 wire _10865_;
 wire _10866_;
 wire _10867_;
 wire _10868_;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire _10872_;
 wire _10873_;
 wire _10874_;
 wire _10875_;
 wire _10876_;
 wire _10877_;
 wire _10878_;
 wire _10879_;
 wire _10880_;
 wire _10881_;
 wire _10882_;
 wire _10883_;
 wire _10884_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire _10889_;
 wire _10890_;
 wire _10891_;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire _10903_;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire _10907_;
 wire _10908_;
 wire _10909_;
 wire _10910_;
 wire _10911_;
 wire _10912_;
 wire _10913_;
 wire _10914_;
 wire _10915_;
 wire _10916_;
 wire _10917_;
 wire _10918_;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10922_;
 wire _10923_;
 wire _10924_;
 wire _10925_;
 wire _10926_;
 wire _10927_;
 wire _10928_;
 wire _10929_;
 wire _10930_;
 wire _10931_;
 wire _10932_;
 wire _10933_;
 wire _10934_;
 wire _10935_;
 wire _10936_;
 wire _10937_;
 wire _10938_;
 wire _10939_;
 wire _10940_;
 wire _10941_;
 wire _10942_;
 wire _10943_;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire _10947_;
 wire _10948_;
 wire _10949_;
 wire _10950_;
 wire _10951_;
 wire _10952_;
 wire _10953_;
 wire _10954_;
 wire _10955_;
 wire _10956_;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire _10960_;
 wire _10961_;
 wire _10962_;
 wire _10963_;
 wire _10964_;
 wire _10965_;
 wire _10966_;
 wire _10967_;
 wire _10968_;
 wire _10969_;
 wire _10970_;
 wire _10971_;
 wire _10972_;
 wire _10973_;
 wire _10974_;
 wire _10975_;
 wire _10976_;
 wire _10977_;
 wire _10978_;
 wire _10979_;
 wire _10980_;
 wire _10981_;
 wire _10982_;
 wire _10983_;
 wire _10984_;
 wire _10985_;
 wire _10986_;
 wire _10987_;
 wire _10988_;
 wire _10989_;
 wire _10990_;
 wire _10991_;
 wire _10992_;
 wire _10993_;
 wire _10994_;
 wire _10995_;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire _10999_;
 wire _11000_;
 wire _11001_;
 wire _11002_;
 wire _11003_;
 wire _11004_;
 wire _11005_;
 wire _11006_;
 wire _11007_;
 wire _11008_;
 wire _11009_;
 wire _11010_;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire _11015_;
 wire _11016_;
 wire _11017_;
 wire _11018_;
 wire _11019_;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire _11025_;
 wire _11026_;
 wire _11027_;
 wire _11028_;
 wire _11029_;
 wire _11030_;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire _11034_;
 wire _11035_;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire _11043_;
 wire _11044_;
 wire _11045_;
 wire _11046_;
 wire _11047_;
 wire _11048_;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11052_;
 wire _11053_;
 wire _11054_;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire _11058_;
 wire _11059_;
 wire _11060_;
 wire _11061_;
 wire _11062_;
 wire _11063_;
 wire _11064_;
 wire _11065_;
 wire _11066_;
 wire _11067_;
 wire _11068_;
 wire _11069_;
 wire _11070_;
 wire _11071_;
 wire _11072_;
 wire _11073_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire _11077_;
 wire _11078_;
 wire _11079_;
 wire _11080_;
 wire _11081_;
 wire _11082_;
 wire _11083_;
 wire _11084_;
 wire _11085_;
 wire _11086_;
 wire _11087_;
 wire _11088_;
 wire _11089_;
 wire _11090_;
 wire _11091_;
 wire _11092_;
 wire _11093_;
 wire _11094_;
 wire _11095_;
 wire _11096_;
 wire _11097_;
 wire _11098_;
 wire _11099_;
 wire _11100_;
 wire _11101_;
 wire _11102_;
 wire _11103_;
 wire _11104_;
 wire _11105_;
 wire _11106_;
 wire _11107_;
 wire _11108_;
 wire _11109_;
 wire _11110_;
 wire _11111_;
 wire _11112_;
 wire _11113_;
 wire _11114_;
 wire _11115_;
 wire _11116_;
 wire _11117_;
 wire _11118_;
 wire _11119_;
 wire _11120_;
 wire _11121_;
 wire _11122_;
 wire _11123_;
 wire _11124_;
 wire _11125_;
 wire _11126_;
 wire _11127_;
 wire _11128_;
 wire _11129_;
 wire _11130_;
 wire _11131_;
 wire _11132_;
 wire _11133_;
 wire _11134_;
 wire _11135_;
 wire _11136_;
 wire _11137_;
 wire _11138_;
 wire _11139_;
 wire _11140_;
 wire _11141_;
 wire _11142_;
 wire _11143_;
 wire _11144_;
 wire _11145_;
 wire _11146_;
 wire _11147_;
 wire _11148_;
 wire _11149_;
 wire _11150_;
 wire _11151_;
 wire _11152_;
 wire _11153_;
 wire _11154_;
 wire _11155_;
 wire _11156_;
 wire _11157_;
 wire _11158_;
 wire _11159_;
 wire _11160_;
 wire _11161_;
 wire _11162_;
 wire _11163_;
 wire _11164_;
 wire _11165_;
 wire _11166_;
 wire _11167_;
 wire _11168_;
 wire _11169_;
 wire _11170_;
 wire _11171_;
 wire _11172_;
 wire _11173_;
 wire _11174_;
 wire _11175_;
 wire _11176_;
 wire _11177_;
 wire _11178_;
 wire _11179_;
 wire _11180_;
 wire _11181_;
 wire _11182_;
 wire _11183_;
 wire _11184_;
 wire _11185_;
 wire _11186_;
 wire _11187_;
 wire _11188_;
 wire _11189_;
 wire _11190_;
 wire _11191_;
 wire _11192_;
 wire _11193_;
 wire _11194_;
 wire _11195_;
 wire _11196_;
 wire _11197_;
 wire _11198_;
 wire _11199_;
 wire _11200_;
 wire _11201_;
 wire _11202_;
 wire _11203_;
 wire _11204_;
 wire _11206_;
 wire _11207_;
 wire _11208_;
 wire _11209_;
 wire _11210_;
 wire _11211_;
 wire _11212_;
 wire _11213_;
 wire _11214_;
 wire _11215_;
 wire _11216_;
 wire _11217_;
 wire _11218_;
 wire _11219_;
 wire _11220_;
 wire _11221_;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire _11225_;
 wire _11226_;
 wire _11227_;
 wire _11228_;
 wire _11229_;
 wire _11230_;
 wire _11231_;
 wire _11232_;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11237_;
 wire _11238_;
 wire _11239_;
 wire _11240_;
 wire _11241_;
 wire _11242_;
 wire _11243_;
 wire _11244_;
 wire _11245_;
 wire _11246_;
 wire _11247_;
 wire _11248_;
 wire _11249_;
 wire _11250_;
 wire _11251_;
 wire _11252_;
 wire _11253_;
 wire _11254_;
 wire _11255_;
 wire _11256_;
 wire _11257_;
 wire _11258_;
 wire _11259_;
 wire _11260_;
 wire _11261_;
 wire _11262_;
 wire _11263_;
 wire _11264_;
 wire _11265_;
 wire _11266_;
 wire _11267_;
 wire _11268_;
 wire _11269_;
 wire _11270_;
 wire _11271_;
 wire _11272_;
 wire _11273_;
 wire _11274_;
 wire _11275_;
 wire _11276_;
 wire _11277_;
 wire _11278_;
 wire _11279_;
 wire _11280_;
 wire _11281_;
 wire _11282_;
 wire _11283_;
 wire _11284_;
 wire _11285_;
 wire _11286_;
 wire _11287_;
 wire _11288_;
 wire _11289_;
 wire _11290_;
 wire _11291_;
 wire _11292_;
 wire _11293_;
 wire _11294_;
 wire _11295_;
 wire _11296_;
 wire _11297_;
 wire _11298_;
 wire _11299_;
 wire _11300_;
 wire _11301_;
 wire _11302_;
 wire _11303_;
 wire _11304_;
 wire _11305_;
 wire _11306_;
 wire _11307_;
 wire _11308_;
 wire _11309_;
 wire _11310_;
 wire _11311_;
 wire _11312_;
 wire _11313_;
 wire _11314_;
 wire _11315_;
 wire _11316_;
 wire _11317_;
 wire _11318_;
 wire _11319_;
 wire _11320_;
 wire _11321_;
 wire _11322_;
 wire _11323_;
 wire _11324_;
 wire _11325_;
 wire _11326_;
 wire _11327_;
 wire _11328_;
 wire _11329_;
 wire _11330_;
 wire _11331_;
 wire _11332_;
 wire _11333_;
 wire _11334_;
 wire _11335_;
 wire _11336_;
 wire _11337_;
 wire _11338_;
 wire _11339_;
 wire _11340_;
 wire _11341_;
 wire _11342_;
 wire _11343_;
 wire _11344_;
 wire _11345_;
 wire _11346_;
 wire _11347_;
 wire _11348_;
 wire _11349_;
 wire _11350_;
 wire _11351_;
 wire _11352_;
 wire _11353_;
 wire _11354_;
 wire _11355_;
 wire _11356_;
 wire _11357_;
 wire _11358_;
 wire _11359_;
 wire _11360_;
 wire _11361_;
 wire _11362_;
 wire _11363_;
 wire _11364_;
 wire _11365_;
 wire _11366_;
 wire _11367_;
 wire _11368_;
 wire _11369_;
 wire _11370_;
 wire _11371_;
 wire _11372_;
 wire _11373_;
 wire _11374_;
 wire _11375_;
 wire _11376_;
 wire _11377_;
 wire _11378_;
 wire _11379_;
 wire _11380_;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire _11384_;
 wire _11385_;
 wire _11386_;
 wire _11387_;
 wire _11388_;
 wire _11389_;
 wire _11390_;
 wire _11391_;
 wire _11392_;
 wire _11393_;
 wire _11394_;
 wire _11395_;
 wire _11396_;
 wire _11397_;
 wire _11398_;
 wire _11399_;
 wire _11400_;
 wire _11401_;
 wire _11402_;
 wire _11403_;
 wire _11404_;
 wire _11405_;
 wire _11406_;
 wire _11407_;
 wire _11408_;
 wire _11409_;
 wire _11410_;
 wire _11411_;
 wire _11412_;
 wire _11413_;
 wire _11414_;
 wire _11415_;
 wire _11416_;
 wire _11417_;
 wire _11418_;
 wire _11419_;
 wire _11420_;
 wire _11421_;
 wire _11422_;
 wire _11423_;
 wire _11424_;
 wire _11425_;
 wire _11426_;
 wire _11427_;
 wire _11428_;
 wire _11429_;
 wire _11430_;
 wire _11431_;
 wire _11432_;
 wire _11433_;
 wire _11434_;
 wire _11435_;
 wire _11436_;
 wire _11437_;
 wire _11438_;
 wire _11439_;
 wire _11440_;
 wire _11441_;
 wire _11442_;
 wire _11443_;
 wire _11444_;
 wire _11445_;
 wire _11446_;
 wire _11447_;
 wire _11448_;
 wire _11449_;
 wire _11450_;
 wire _11451_;
 wire _11452_;
 wire _11453_;
 wire _11454_;
 wire _11455_;
 wire _11456_;
 wire _11457_;
 wire _11458_;
 wire _11459_;
 wire _11460_;
 wire _11461_;
 wire _11462_;
 wire _11463_;
 wire _11464_;
 wire _11465_;
 wire _11466_;
 wire _11467_;
 wire _11468_;
 wire _11469_;
 wire _11470_;
 wire _11471_;
 wire _11472_;
 wire _11473_;
 wire _11474_;
 wire _11475_;
 wire _11476_;
 wire _11477_;
 wire _11478_;
 wire _11479_;
 wire _11480_;
 wire _11481_;
 wire _11482_;
 wire _11483_;
 wire _11484_;
 wire _11485_;
 wire _11486_;
 wire _11487_;
 wire _11488_;
 wire _11489_;
 wire _11490_;
 wire _11491_;
 wire _11492_;
 wire _11493_;
 wire _11494_;
 wire _11495_;
 wire _11496_;
 wire _11497_;
 wire _11498_;
 wire _11499_;
 wire _11500_;
 wire _11501_;
 wire _11502_;
 wire _11503_;
 wire _11504_;
 wire _11505_;
 wire _11506_;
 wire _11507_;
 wire _11508_;
 wire _11509_;
 wire _11510_;
 wire _11511_;
 wire _11512_;
 wire _11513_;
 wire _11514_;
 wire _11515_;
 wire _11516_;
 wire _11517_;
 wire _11518_;
 wire _11519_;
 wire _11520_;
 wire _11521_;
 wire _11522_;
 wire _11523_;
 wire _11524_;
 wire _11525_;
 wire _11526_;
 wire _11527_;
 wire _11528_;
 wire _11529_;
 wire _11530_;
 wire _11531_;
 wire _11532_;
 wire _11533_;
 wire _11534_;
 wire _11535_;
 wire _11536_;
 wire _11537_;
 wire _11538_;
 wire _11539_;
 wire _11540_;
 wire _11541_;
 wire _11542_;
 wire _11543_;
 wire _11544_;
 wire _11545_;
 wire _11546_;
 wire _11547_;
 wire _11548_;
 wire _11549_;
 wire _11550_;
 wire _11551_;
 wire _11552_;
 wire _11553_;
 wire _11554_;
 wire _11555_;
 wire _11556_;
 wire _11557_;
 wire _11558_;
 wire _11559_;
 wire _11560_;
 wire _11561_;
 wire _11562_;
 wire _11563_;
 wire _11564_;
 wire _11565_;
 wire _11566_;
 wire _11567_;
 wire _11568_;
 wire _11569_;
 wire _11570_;
 wire _11571_;
 wire _11572_;
 wire _11573_;
 wire _11574_;
 wire _11575_;
 wire _11576_;
 wire _11577_;
 wire _11578_;
 wire _11579_;
 wire _11580_;
 wire _11581_;
 wire _11582_;
 wire _11583_;
 wire _11584_;
 wire _11585_;
 wire _11586_;
 wire _11587_;
 wire _11588_;
 wire _11589_;
 wire _11590_;
 wire _11591_;
 wire _11592_;
 wire _11593_;
 wire _11594_;
 wire _11595_;
 wire _11596_;
 wire _11597_;
 wire _11598_;
 wire _11599_;
 wire _11600_;
 wire _11601_;
 wire _11602_;
 wire _11603_;
 wire _11604_;
 wire _11605_;
 wire _11606_;
 wire _11607_;
 wire _11608_;
 wire _11609_;
 wire _11610_;
 wire _11611_;
 wire _11612_;
 wire _11613_;
 wire _11614_;
 wire _11615_;
 wire _11616_;
 wire _11617_;
 wire _11618_;
 wire _11619_;
 wire _11620_;
 wire _11621_;
 wire _11622_;
 wire _11623_;
 wire _11624_;
 wire _11625_;
 wire _11626_;
 wire _11627_;
 wire _11628_;
 wire _11629_;
 wire _11630_;
 wire _11631_;
 wire _11632_;
 wire _11633_;
 wire _11634_;
 wire _11635_;
 wire _11636_;
 wire _11637_;
 wire _11638_;
 wire _11639_;
 wire _11640_;
 wire _11641_;
 wire _11642_;
 wire _11643_;
 wire _11644_;
 wire _11645_;
 wire _11646_;
 wire _11647_;
 wire _11648_;
 wire _11649_;
 wire _11650_;
 wire _11651_;
 wire _11652_;
 wire _11653_;
 wire _11654_;
 wire _11655_;
 wire _11656_;
 wire _11657_;
 wire _11658_;
 wire _11659_;
 wire _11660_;
 wire _11661_;
 wire _11662_;
 wire _11663_;
 wire _11664_;
 wire _11665_;
 wire _11666_;
 wire _11667_;
 wire _11668_;
 wire _11669_;
 wire _11670_;
 wire _11671_;
 wire _11672_;
 wire _11673_;
 wire _11674_;
 wire _11675_;
 wire _11676_;
 wire _11677_;
 wire _11678_;
 wire _11679_;
 wire _11680_;
 wire _11681_;
 wire _11682_;
 wire _11683_;
 wire _11684_;
 wire _11685_;
 wire _11686_;
 wire _11687_;
 wire _11688_;
 wire _11689_;
 wire _11690_;
 wire _11691_;
 wire _11692_;
 wire _11693_;
 wire _11694_;
 wire _11695_;
 wire _11696_;
 wire _11697_;
 wire _11698_;
 wire _11699_;
 wire _11700_;
 wire _11701_;
 wire _11702_;
 wire _11703_;
 wire _11704_;
 wire _11705_;
 wire _11706_;
 wire _11707_;
 wire _11708_;
 wire _11709_;
 wire _11710_;
 wire _11711_;
 wire _11712_;
 wire _11713_;
 wire _11714_;
 wire _11715_;
 wire _11716_;
 wire _11717_;
 wire _11718_;
 wire _11719_;
 wire _11720_;
 wire _11721_;
 wire _11722_;
 wire _11723_;
 wire _11724_;
 wire _11725_;
 wire _11726_;
 wire _11727_;
 wire _11728_;
 wire _11729_;
 wire _11730_;
 wire _11731_;
 wire _11732_;
 wire _11733_;
 wire _11734_;
 wire _11735_;
 wire _11736_;
 wire _11737_;
 wire _11738_;
 wire _11739_;
 wire _11740_;
 wire _11741_;
 wire _11742_;
 wire _11743_;
 wire _11744_;
 wire _11745_;
 wire _11746_;
 wire _11747_;
 wire _11748_;
 wire _11749_;
 wire _11750_;
 wire _11751_;
 wire _11752_;
 wire _11753_;
 wire _11754_;
 wire _11755_;
 wire _11756_;
 wire _11757_;
 wire _11758_;
 wire _11759_;
 wire _11760_;
 wire _11761_;
 wire _11762_;
 wire _11763_;
 wire _11764_;
 wire _11765_;
 wire _11766_;
 wire _11767_;
 wire _11768_;
 wire _11769_;
 wire _11770_;
 wire _11771_;
 wire _11772_;
 wire _11773_;
 wire _11774_;
 wire _11775_;
 wire _11776_;
 wire _11777_;
 wire _11778_;
 wire _11779_;
 wire _11780_;
 wire _11781_;
 wire _11782_;
 wire _11783_;
 wire _11784_;
 wire _11785_;
 wire _11786_;
 wire _11787_;
 wire _11788_;
 wire _11789_;
 wire _11790_;
 wire _11791_;
 wire _11792_;
 wire _11793_;
 wire _11794_;
 wire _11795_;
 wire _11796_;
 wire _11797_;
 wire _11798_;
 wire _11799_;
 wire _11800_;
 wire _11801_;
 wire _11802_;
 wire _11803_;
 wire _11804_;
 wire _11805_;
 wire _11806_;
 wire _11807_;
 wire _11808_;
 wire _11809_;
 wire _11810_;
 wire _11811_;
 wire _11812_;
 wire _11813_;
 wire _11814_;
 wire _11815_;
 wire _11816_;
 wire _11817_;
 wire _11818_;
 wire _11819_;
 wire _11820_;
 wire _11821_;
 wire _11822_;
 wire _11823_;
 wire _11824_;
 wire _11825_;
 wire _11826_;
 wire _11827_;
 wire _11828_;
 wire _11829_;
 wire _11830_;
 wire _11831_;
 wire _11832_;
 wire _11833_;
 wire _11834_;
 wire _11835_;
 wire _11836_;
 wire _11837_;
 wire _11838_;
 wire _11839_;
 wire _11840_;
 wire _11841_;
 wire _11842_;
 wire _11843_;
 wire _11844_;
 wire _11845_;
 wire _11846_;
 wire _11847_;
 wire _11848_;
 wire _11849_;
 wire _11850_;
 wire _11851_;
 wire _11852_;
 wire _11853_;
 wire _11854_;
 wire _11855_;
 wire _11856_;
 wire _11857_;
 wire _11858_;
 wire _11859_;
 wire _11860_;
 wire _11861_;
 wire _11862_;
 wire _11863_;
 wire _11864_;
 wire _11865_;
 wire _11866_;
 wire _11867_;
 wire _11868_;
 wire _11869_;
 wire _11870_;
 wire _11871_;
 wire _11872_;
 wire _11873_;
 wire _11874_;
 wire _11875_;
 wire _11876_;
 wire _11877_;
 wire _11878_;
 wire _11879_;
 wire _11880_;
 wire _11881_;
 wire _11882_;
 wire _11883_;
 wire _11884_;
 wire _11885_;
 wire _11886_;
 wire _11887_;
 wire _11888_;
 wire _11889_;
 wire _11890_;
 wire _11891_;
 wire _11892_;
 wire _11893_;
 wire _11894_;
 wire _11895_;
 wire _11896_;
 wire _11897_;
 wire _11898_;
 wire _11899_;
 wire _11900_;
 wire _11901_;
 wire _11902_;
 wire _11903_;
 wire _11904_;
 wire _11905_;
 wire _11906_;
 wire _11907_;
 wire _11908_;
 wire _11909_;
 wire _11910_;
 wire _11911_;
 wire _11912_;
 wire _11913_;
 wire _11914_;
 wire _11915_;
 wire _11916_;
 wire _11917_;
 wire _11918_;
 wire _11919_;
 wire _11920_;
 wire _11921_;
 wire _11922_;
 wire _11923_;
 wire _11924_;
 wire _11925_;
 wire _11926_;
 wire _11927_;
 wire _11928_;
 wire _11929_;
 wire _11930_;
 wire _11931_;
 wire _11932_;
 wire _11933_;
 wire _11934_;
 wire _11935_;
 wire _11936_;
 wire _11937_;
 wire _11938_;
 wire _11939_;
 wire _11940_;
 wire _11941_;
 wire _11942_;
 wire _11943_;
 wire _11944_;
 wire _11945_;
 wire _11946_;
 wire _11947_;
 wire _11948_;
 wire _11949_;
 wire _11950_;
 wire _11951_;
 wire _11952_;
 wire _11953_;
 wire _11954_;
 wire _11955_;
 wire _11956_;
 wire _11957_;
 wire _11958_;
 wire _11959_;
 wire _11960_;
 wire _11961_;
 wire _11962_;
 wire _11963_;
 wire _11964_;
 wire _11965_;
 wire _11966_;
 wire _11967_;
 wire _11968_;
 wire _11969_;
 wire _11970_;
 wire _11971_;
 wire _11972_;
 wire _11973_;
 wire _11974_;
 wire _11975_;
 wire _11976_;
 wire _11977_;
 wire _11978_;
 wire _11979_;
 wire _11980_;
 wire _11981_;
 wire _11982_;
 wire _11983_;
 wire _11984_;
 wire _11985_;
 wire _11986_;
 wire _11987_;
 wire _11988_;
 wire _11989_;
 wire _11990_;
 wire _11991_;
 wire _11992_;
 wire _11993_;
 wire _11994_;
 wire _11995_;
 wire _11996_;
 wire _11997_;
 wire _11998_;
 wire _11999_;
 wire _12000_;
 wire _12001_;
 wire _12002_;
 wire _12003_;
 wire _12004_;
 wire _12005_;
 wire _12006_;
 wire _12007_;
 wire _12008_;
 wire _12009_;
 wire _12010_;
 wire _12011_;
 wire _12012_;
 wire _12013_;
 wire _12014_;
 wire _12015_;
 wire _12016_;
 wire _12017_;
 wire _12018_;
 wire _12019_;
 wire _12020_;
 wire _12021_;
 wire _12022_;
 wire _12023_;
 wire _12024_;
 wire _12025_;
 wire _12026_;
 wire _12027_;
 wire _12028_;
 wire _12029_;
 wire _12030_;
 wire _12031_;
 wire _12032_;
 wire _12033_;
 wire _12034_;
 wire _12035_;
 wire _12036_;
 wire _12037_;
 wire _12038_;
 wire _12039_;
 wire _12040_;
 wire _12041_;
 wire _12042_;
 wire _12043_;
 wire _12044_;
 wire _12045_;
 wire _12046_;
 wire _12047_;
 wire _12048_;
 wire _12049_;
 wire _12050_;
 wire _12051_;
 wire _12052_;
 wire _12053_;
 wire _12054_;
 wire _12055_;
 wire _12056_;
 wire _12057_;
 wire _12058_;
 wire _12059_;
 wire _12060_;
 wire _12061_;
 wire _12062_;
 wire _12063_;
 wire _12064_;
 wire _12065_;
 wire _12066_;
 wire _12067_;
 wire _12068_;
 wire _12069_;
 wire _12070_;
 wire _12071_;
 wire _12072_;
 wire _12073_;
 wire _12074_;
 wire _12075_;
 wire _12076_;
 wire _12077_;
 wire _12078_;
 wire _12079_;
 wire _12080_;
 wire _12081_;
 wire _12082_;
 wire _12083_;
 wire _12084_;
 wire _12085_;
 wire _12086_;
 wire _12087_;
 wire _12088_;
 wire _12089_;
 wire _12090_;
 wire _12091_;
 wire _12092_;
 wire _12093_;
 wire _12094_;
 wire _12095_;
 wire _12096_;
 wire _12097_;
 wire _12098_;
 wire _12099_;
 wire _12100_;
 wire _12101_;
 wire _12102_;
 wire _12103_;
 wire _12104_;
 wire _12105_;
 wire _12106_;
 wire _12107_;
 wire _12108_;
 wire _12109_;
 wire _12110_;
 wire _12111_;
 wire _12112_;
 wire _12113_;
 wire _12114_;
 wire _12115_;
 wire _12116_;
 wire _12117_;
 wire _12118_;
 wire _12119_;
 wire _12120_;
 wire _12121_;
 wire _12122_;
 wire _12123_;
 wire _12124_;
 wire _12125_;
 wire _12126_;
 wire _12127_;
 wire _12128_;
 wire _12129_;
 wire _12130_;
 wire _12131_;
 wire _12132_;
 wire _12133_;
 wire _12134_;
 wire _12135_;
 wire _12136_;
 wire _12137_;
 wire _12138_;
 wire _12139_;
 wire _12140_;
 wire _12141_;
 wire _12142_;
 wire _12143_;
 wire _12144_;
 wire _12145_;
 wire _12146_;
 wire _12147_;
 wire _12148_;
 wire _12149_;
 wire _12150_;
 wire _12151_;
 wire _12152_;
 wire _12153_;
 wire _12154_;
 wire _12155_;
 wire _12156_;
 wire _12157_;
 wire _12158_;
 wire _12159_;
 wire _12160_;
 wire _12161_;
 wire _12162_;
 wire _12163_;
 wire _12164_;
 wire _12165_;
 wire _12166_;
 wire _12167_;
 wire _12168_;
 wire _12169_;
 wire _12170_;
 wire _12171_;
 wire _12172_;
 wire _12173_;
 wire _12174_;
 wire _12175_;
 wire _12176_;
 wire _12177_;
 wire _12178_;
 wire _12179_;
 wire _12180_;
 wire _12181_;
 wire _12182_;
 wire _12183_;
 wire _12184_;
 wire _12185_;
 wire _12186_;
 wire _12187_;
 wire _12188_;
 wire _12189_;
 wire _12190_;
 wire _12191_;
 wire _12192_;
 wire _12193_;
 wire _12194_;
 wire _12195_;
 wire _12196_;
 wire _12197_;
 wire _12198_;
 wire _12199_;
 wire _12200_;
 wire _12201_;
 wire _12202_;
 wire _12203_;
 wire _12204_;
 wire _12205_;
 wire _12206_;
 wire _12207_;
 wire _12208_;
 wire _12209_;
 wire _12210_;
 wire _12211_;
 wire _12212_;
 wire _12213_;
 wire _12214_;
 wire _12215_;
 wire _12216_;
 wire _12217_;
 wire _12218_;
 wire _12219_;
 wire _12220_;
 wire _12221_;
 wire _12222_;
 wire _12223_;
 wire _12224_;
 wire _12225_;
 wire _12226_;
 wire _12227_;
 wire _12228_;
 wire _12229_;
 wire _12230_;
 wire _12231_;
 wire _12232_;
 wire _12233_;
 wire _12234_;
 wire _12235_;
 wire _12236_;
 wire _12237_;
 wire _12238_;
 wire _12239_;
 wire _12240_;
 wire _12241_;
 wire _12242_;
 wire _12243_;
 wire _12244_;
 wire _12245_;
 wire _12246_;
 wire _12247_;
 wire _12248_;
 wire _12249_;
 wire _12250_;
 wire _12251_;
 wire _12252_;
 wire _12253_;
 wire _12254_;
 wire _12255_;
 wire _12256_;
 wire _12257_;
 wire _12258_;
 wire _12259_;
 wire _12260_;
 wire _12261_;
 wire _12262_;
 wire _12263_;
 wire _12264_;
 wire _12265_;
 wire _12266_;
 wire _12267_;
 wire _12268_;
 wire _12269_;
 wire _12270_;
 wire _12271_;
 wire _12272_;
 wire _12273_;
 wire _12274_;
 wire _12275_;
 wire _12276_;
 wire _12277_;
 wire _12278_;
 wire _12279_;
 wire _12280_;
 wire _12281_;
 wire _12282_;
 wire _12283_;
 wire _12284_;
 wire _12285_;
 wire _12287_;
 wire _12288_;
 wire _12289_;
 wire _12290_;
 wire _12291_;
 wire _12292_;
 wire _12293_;
 wire _12294_;
 wire _12295_;
 wire _12296_;
 wire _12297_;
 wire _12298_;
 wire _12299_;
 wire _12300_;
 wire _12301_;
 wire _12302_;
 wire _12303_;
 wire _12304_;
 wire _12305_;
 wire _12306_;
 wire _12307_;
 wire _12308_;
 wire _12309_;
 wire _12310_;
 wire _12311_;
 wire _12312_;
 wire _12313_;
 wire _12314_;
 wire _12315_;
 wire _12316_;
 wire _12317_;
 wire _12318_;
 wire _12319_;
 wire _12320_;
 wire _12321_;
 wire _12322_;
 wire _12323_;
 wire _12324_;
 wire _12325_;
 wire _12326_;
 wire _12327_;
 wire _12328_;
 wire _12329_;
 wire _12330_;
 wire _12331_;
 wire _12332_;
 wire _12333_;
 wire _12334_;
 wire _12335_;
 wire _12336_;
 wire _12337_;
 wire _12338_;
 wire _12339_;
 wire _12340_;
 wire _12341_;
 wire _12342_;
 wire _12343_;
 wire _12344_;
 wire _12345_;
 wire _12346_;
 wire _12347_;
 wire _12348_;
 wire _12349_;
 wire _12350_;
 wire _12351_;
 wire _12352_;
 wire _12353_;
 wire _12354_;
 wire _12355_;
 wire _12356_;
 wire _12357_;
 wire _12358_;
 wire _12359_;
 wire _12360_;
 wire _12361_;
 wire _12362_;
 wire _12363_;
 wire _12364_;
 wire _12365_;
 wire _12366_;
 wire _12367_;
 wire _12368_;
 wire _12369_;
 wire _12370_;
 wire _12371_;
 wire _12372_;
 wire _12373_;
 wire _12374_;
 wire _12375_;
 wire _12376_;
 wire _12377_;
 wire _12378_;
 wire _12379_;
 wire _12380_;
 wire _12381_;
 wire _12382_;
 wire _12383_;
 wire _12384_;
 wire _12385_;
 wire _12386_;
 wire _12387_;
 wire _12388_;
 wire _12389_;
 wire _12390_;
 wire _12391_;
 wire _12392_;
 wire _12393_;
 wire _12394_;
 wire _12395_;
 wire _12396_;
 wire _12397_;
 wire _12398_;
 wire _12399_;
 wire _12400_;
 wire _12401_;
 wire _12402_;
 wire _12403_;
 wire _12404_;
 wire _12405_;
 wire _12406_;
 wire _12407_;
 wire _12408_;
 wire _12409_;
 wire _12410_;
 wire _12411_;
 wire _12412_;
 wire _12413_;
 wire _12414_;
 wire _12415_;
 wire _12416_;
 wire _12417_;
 wire _12418_;
 wire _12419_;
 wire _12420_;
 wire _12421_;
 wire _12422_;
 wire _12423_;
 wire _12424_;
 wire _12425_;
 wire _12426_;
 wire _12427_;
 wire _12428_;
 wire _12429_;
 wire _12430_;
 wire _12431_;
 wire _12432_;
 wire _12433_;
 wire _12434_;
 wire _12435_;
 wire _12436_;
 wire _12437_;
 wire _12438_;
 wire _12439_;
 wire _12440_;
 wire _12441_;
 wire _12442_;
 wire _12443_;
 wire _12444_;
 wire _12445_;
 wire _12446_;
 wire _12447_;
 wire _12448_;
 wire _12449_;
 wire _12450_;
 wire _12451_;
 wire _12452_;
 wire _12453_;
 wire _12454_;
 wire _12455_;
 wire _12456_;
 wire _12457_;
 wire _12458_;
 wire _12459_;
 wire _12460_;
 wire _12461_;
 wire _12462_;
 wire _12463_;
 wire _12464_;
 wire _12465_;
 wire _12466_;
 wire _12467_;
 wire _12468_;
 wire _12469_;
 wire _12470_;
 wire _12471_;
 wire _12472_;
 wire _12473_;
 wire _12474_;
 wire _12475_;
 wire _12476_;
 wire _12477_;
 wire _12478_;
 wire _12479_;
 wire _12480_;
 wire _12481_;
 wire _12482_;
 wire _12483_;
 wire _12484_;
 wire _12485_;
 wire _12486_;
 wire _12487_;
 wire _12488_;
 wire _12489_;
 wire _12490_;
 wire _12491_;
 wire _12492_;
 wire _12493_;
 wire _12494_;
 wire _12495_;
 wire _12496_;
 wire _12497_;
 wire _12498_;
 wire _12499_;
 wire _12500_;
 wire _12501_;
 wire _12502_;
 wire _12503_;
 wire _12504_;
 wire _12505_;
 wire _12506_;
 wire _12507_;
 wire _12508_;
 wire _12509_;
 wire _12510_;
 wire _12511_;
 wire _12512_;
 wire _12513_;
 wire _12514_;
 wire _12515_;
 wire _12516_;
 wire _12517_;
 wire _12518_;
 wire _12519_;
 wire _12520_;
 wire _12521_;
 wire _12522_;
 wire _12523_;
 wire _12524_;
 wire _12525_;
 wire _12526_;
 wire _12527_;
 wire _12528_;
 wire _12529_;
 wire _12530_;
 wire _12531_;
 wire _12532_;
 wire _12533_;
 wire _12534_;
 wire _12535_;
 wire _12536_;
 wire _12537_;
 wire _12538_;
 wire _12539_;
 wire _12540_;
 wire _12541_;
 wire _12542_;
 wire _12543_;
 wire _12544_;
 wire _12545_;
 wire _12546_;
 wire _12547_;
 wire _12548_;
 wire _12549_;
 wire _12550_;
 wire _12551_;
 wire _12552_;
 wire _12553_;
 wire _12554_;
 wire _12555_;
 wire _12556_;
 wire _12557_;
 wire _12558_;
 wire _12559_;
 wire _12560_;
 wire _12561_;
 wire _12562_;
 wire _12563_;
 wire _12564_;
 wire _12565_;
 wire _12566_;
 wire _12567_;
 wire _12568_;
 wire _12569_;
 wire _12570_;
 wire _12571_;
 wire _12572_;
 wire _12573_;
 wire _12574_;
 wire _12575_;
 wire _12576_;
 wire _12577_;
 wire _12578_;
 wire _12579_;
 wire _12580_;
 wire _12581_;
 wire _12582_;
 wire _12583_;
 wire _12584_;
 wire _12585_;
 wire _12586_;
 wire _12587_;
 wire _12588_;
 wire _12589_;
 wire _12590_;
 wire _12591_;
 wire _12592_;
 wire _12593_;
 wire _12594_;
 wire _12595_;
 wire _12596_;
 wire _12597_;
 wire _12598_;
 wire _12599_;
 wire _12600_;
 wire _12601_;
 wire _12602_;
 wire _12603_;
 wire _12604_;
 wire _12605_;
 wire _12606_;
 wire _12607_;
 wire _12608_;
 wire _12609_;
 wire _12610_;
 wire _12611_;
 wire _12612_;
 wire _12613_;
 wire _12614_;
 wire _12615_;
 wire _12616_;
 wire _12617_;
 wire _12618_;
 wire _12619_;
 wire _12620_;
 wire _12621_;
 wire _12622_;
 wire _12623_;
 wire _12624_;
 wire _12625_;
 wire _12626_;
 wire _12627_;
 wire _12628_;
 wire _12629_;
 wire _12630_;
 wire _12631_;
 wire _12632_;
 wire _12633_;
 wire _12634_;
 wire _12635_;
 wire _12636_;
 wire _12637_;
 wire _12638_;
 wire _12639_;
 wire _12640_;
 wire _12641_;
 wire _12642_;
 wire _12643_;
 wire _12644_;
 wire _12645_;
 wire _12646_;
 wire _12647_;
 wire _12648_;
 wire _12649_;
 wire _12650_;
 wire _12651_;
 wire _12652_;
 wire _12653_;
 wire _12654_;
 wire _12655_;
 wire _12656_;
 wire _12657_;
 wire _12658_;
 wire _12659_;
 wire _12660_;
 wire _12661_;
 wire _12662_;
 wire _12663_;
 wire _12664_;
 wire _12665_;
 wire _12666_;
 wire _12667_;
 wire _12668_;
 wire _12669_;
 wire _12670_;
 wire _12671_;
 wire _12672_;
 wire _12673_;
 wire _12674_;
 wire _12675_;
 wire _12676_;
 wire _12677_;
 wire _12678_;
 wire _12679_;
 wire _12680_;
 wire _12681_;
 wire _12682_;
 wire _12683_;
 wire _12684_;
 wire _12685_;
 wire _12686_;
 wire _12687_;
 wire _12688_;
 wire _12689_;
 wire _12690_;
 wire _12691_;
 wire _12692_;
 wire _12693_;
 wire _12694_;
 wire _12695_;
 wire _12696_;
 wire _12697_;
 wire _12698_;
 wire _12699_;
 wire _12700_;
 wire _12701_;
 wire _12702_;
 wire _12703_;
 wire _12704_;
 wire _12705_;
 wire _12706_;
 wire _12707_;
 wire _12708_;
 wire _12709_;
 wire _12710_;
 wire _12711_;
 wire _12712_;
 wire _12713_;
 wire _12714_;
 wire _12715_;
 wire _12716_;
 wire _12717_;
 wire _12718_;
 wire _12719_;
 wire _12720_;
 wire _12721_;
 wire _12722_;
 wire _12723_;
 wire _12724_;
 wire _12725_;
 wire _12726_;
 wire _12727_;
 wire _12728_;
 wire _12729_;
 wire _12730_;
 wire _12731_;
 wire _12732_;
 wire _12733_;
 wire _12734_;
 wire _12735_;
 wire _12736_;
 wire _12737_;
 wire _12738_;
 wire _12739_;
 wire _12740_;
 wire _12741_;
 wire _12742_;
 wire _12743_;
 wire _12744_;
 wire _12745_;
 wire _12746_;
 wire _12747_;
 wire _12748_;
 wire _12749_;
 wire _12750_;
 wire _12751_;
 wire _12752_;
 wire _12753_;
 wire _12754_;
 wire _12755_;
 wire _12756_;
 wire _12757_;
 wire _12758_;
 wire _12759_;
 wire _12760_;
 wire _12761_;
 wire _12762_;
 wire _12763_;
 wire _12764_;
 wire _12765_;
 wire _12766_;
 wire _12767_;
 wire _12768_;
 wire _12769_;
 wire _12770_;
 wire _12771_;
 wire _12772_;
 wire _12773_;
 wire _12774_;
 wire _12775_;
 wire _12776_;
 wire _12777_;
 wire _12778_;
 wire _12779_;
 wire _12780_;
 wire _12781_;
 wire _12782_;
 wire _12783_;
 wire _12784_;
 wire _12785_;
 wire _12786_;
 wire _12787_;
 wire _12788_;
 wire _12789_;
 wire _12790_;
 wire _12791_;
 wire _12792_;
 wire _12793_;
 wire _12794_;
 wire _12795_;
 wire _12796_;
 wire _12797_;
 wire _12798_;
 wire _12799_;
 wire _12800_;
 wire _12801_;
 wire _12802_;
 wire _12803_;
 wire _12804_;
 wire _12805_;
 wire _12806_;
 wire _12807_;
 wire _12808_;
 wire _12809_;
 wire _12810_;
 wire _12811_;
 wire _12812_;
 wire _12813_;
 wire _12814_;
 wire _12815_;
 wire _12816_;
 wire _12817_;
 wire _12818_;
 wire _12819_;
 wire _12820_;
 wire _12821_;
 wire _12822_;
 wire _12823_;
 wire _12824_;
 wire _12825_;
 wire _12826_;
 wire _12827_;
 wire _12828_;
 wire _12829_;
 wire _12830_;
 wire _12831_;
 wire _12832_;
 wire _12833_;
 wire _12834_;
 wire _12835_;
 wire _12836_;
 wire _12837_;
 wire _12838_;
 wire _12839_;
 wire _12840_;
 wire _12841_;
 wire _12842_;
 wire _12843_;
 wire _12844_;
 wire _12845_;
 wire _12846_;
 wire _12847_;
 wire _12848_;
 wire _12849_;
 wire _12850_;
 wire _12851_;
 wire _12852_;
 wire _12853_;
 wire _12854_;
 wire _12855_;
 wire _12856_;
 wire _12857_;
 wire _12858_;
 wire _12859_;
 wire _12860_;
 wire _12861_;
 wire _12862_;
 wire _12863_;
 wire _12864_;
 wire _12865_;
 wire _12866_;
 wire _12867_;
 wire _12868_;
 wire _12869_;
 wire _12870_;
 wire _12871_;
 wire _12872_;
 wire _12873_;
 wire _12874_;
 wire _12875_;
 wire _12876_;
 wire _12877_;
 wire _12878_;
 wire _12879_;
 wire _12880_;
 wire _12881_;
 wire _12882_;
 wire _12883_;
 wire _12884_;
 wire _12885_;
 wire _12886_;
 wire _12887_;
 wire _12888_;
 wire _12889_;
 wire _12890_;
 wire _12891_;
 wire _12892_;
 wire _12893_;
 wire _12894_;
 wire _12895_;
 wire _12896_;
 wire _12897_;
 wire _12898_;
 wire _12899_;
 wire _12900_;
 wire _12901_;
 wire _12902_;
 wire _12903_;
 wire _12904_;
 wire _12905_;
 wire _12906_;
 wire _12907_;
 wire _12908_;
 wire _12909_;
 wire _12910_;
 wire _12911_;
 wire _12912_;
 wire _12913_;
 wire _12914_;
 wire _12915_;
 wire _12916_;
 wire _12917_;
 wire _12918_;
 wire _12919_;
 wire _12920_;
 wire _12921_;
 wire _12922_;
 wire _12923_;
 wire _12924_;
 wire _12925_;
 wire _12926_;
 wire _12927_;
 wire _12928_;
 wire _12929_;
 wire _12930_;
 wire _12931_;
 wire _12932_;
 wire _12933_;
 wire _12934_;
 wire _12935_;
 wire _12936_;
 wire _12937_;
 wire _12938_;
 wire _12939_;
 wire _12940_;
 wire _12941_;
 wire _12942_;
 wire _12943_;
 wire _12944_;
 wire _12945_;
 wire _12946_;
 wire _12947_;
 wire _12948_;
 wire _12949_;
 wire _12950_;
 wire _12951_;
 wire _12952_;
 wire _12953_;
 wire _12954_;
 wire _12955_;
 wire _12956_;
 wire _12957_;
 wire _12958_;
 wire _12959_;
 wire _12960_;
 wire _12961_;
 wire _12962_;
 wire _12963_;
 wire _12964_;
 wire _12965_;
 wire _12966_;
 wire _12967_;
 wire _12968_;
 wire _12969_;
 wire _12970_;
 wire _12971_;
 wire _12972_;
 wire _12973_;
 wire _12974_;
 wire _12975_;
 wire _12976_;
 wire _12977_;
 wire _12978_;
 wire _12979_;
 wire _12980_;
 wire _12981_;
 wire _12982_;
 wire _12983_;
 wire _12984_;
 wire _12985_;
 wire _12986_;
 wire _12987_;
 wire _12988_;
 wire _12989_;
 wire _12990_;
 wire _12991_;
 wire _12992_;
 wire _12993_;
 wire _12994_;
 wire _12995_;
 wire _12996_;
 wire _12997_;
 wire _12998_;
 wire _12999_;
 wire _13000_;
 wire _13001_;
 wire _13002_;
 wire _13003_;
 wire _13004_;
 wire _13005_;
 wire _13006_;
 wire _13007_;
 wire _13008_;
 wire _13009_;
 wire _13010_;
 wire _13011_;
 wire _13012_;
 wire _13013_;
 wire _13014_;
 wire _13015_;
 wire _13016_;
 wire _13017_;
 wire _13018_;
 wire _13019_;
 wire _13020_;
 wire _13021_;
 wire _13022_;
 wire _13023_;
 wire _13024_;
 wire _13025_;
 wire _13026_;
 wire _13027_;
 wire _13028_;
 wire _13029_;
 wire _13030_;
 wire _13031_;
 wire _13032_;
 wire _13033_;
 wire _13034_;
 wire _13035_;
 wire _13036_;
 wire _13037_;
 wire _13038_;
 wire _13039_;
 wire _13040_;
 wire _13041_;
 wire _13042_;
 wire _13043_;
 wire _13044_;
 wire _13045_;
 wire _13046_;
 wire _13047_;
 wire _13048_;
 wire _13049_;
 wire _13050_;
 wire _13051_;
 wire _13052_;
 wire _13053_;
 wire _13054_;
 wire _13055_;
 wire _13056_;
 wire _13057_;
 wire _13058_;
 wire _13059_;
 wire _13060_;
 wire _13061_;
 wire _13062_;
 wire _13063_;
 wire _13064_;
 wire _13065_;
 wire _13066_;
 wire _13067_;
 wire _13068_;
 wire _13069_;
 wire _13070_;
 wire _13071_;
 wire _13072_;
 wire _13073_;
 wire _13074_;
 wire _13075_;
 wire _13076_;
 wire _13077_;
 wire _13078_;
 wire _13079_;
 wire _13080_;
 wire _13081_;
 wire _13082_;
 wire _13083_;
 wire _13084_;
 wire _13085_;
 wire _13086_;
 wire _13087_;
 wire _13088_;
 wire _13089_;
 wire _13090_;
 wire _13091_;
 wire _13092_;
 wire _13093_;
 wire _13094_;
 wire _13095_;
 wire _13096_;
 wire _13097_;
 wire _13098_;
 wire _13099_;
 wire _13100_;
 wire _13101_;
 wire _13102_;
 wire _13103_;
 wire _13104_;
 wire _13105_;
 wire _13106_;
 wire _13107_;
 wire _13108_;
 wire _13109_;
 wire _13110_;
 wire _13111_;
 wire _13112_;
 wire _13113_;
 wire _13114_;
 wire _13115_;
 wire _13116_;
 wire _13117_;
 wire _13118_;
 wire _13119_;
 wire _13120_;
 wire _13121_;
 wire _13122_;
 wire _13123_;
 wire _13124_;
 wire _13125_;
 wire _13126_;
 wire _13127_;
 wire _13128_;
 wire _13129_;
 wire _13130_;
 wire _13131_;
 wire _13132_;
 wire _13133_;
 wire _13134_;
 wire _13135_;
 wire _13136_;
 wire _13137_;
 wire _13138_;
 wire _13139_;
 wire _13140_;
 wire _13141_;
 wire _13142_;
 wire _13143_;
 wire _13144_;
 wire _13145_;
 wire _13146_;
 wire _13147_;
 wire _13148_;
 wire _13149_;
 wire _13150_;
 wire _13151_;
 wire _13152_;
 wire _13153_;
 wire _13154_;
 wire _13155_;
 wire _13156_;
 wire _13157_;
 wire _13158_;
 wire _13159_;
 wire _13160_;
 wire _13161_;
 wire _13162_;
 wire _13163_;
 wire _13164_;
 wire _13165_;
 wire _13166_;
 wire _13167_;
 wire _13168_;
 wire _13169_;
 wire _13170_;
 wire _13171_;
 wire _13172_;
 wire _13173_;
 wire _13174_;
 wire _13175_;
 wire _13176_;
 wire _13177_;
 wire _13178_;
 wire _13179_;
 wire _13180_;
 wire _13181_;
 wire _13182_;
 wire _13183_;
 wire _13184_;
 wire _13185_;
 wire _13186_;
 wire _13187_;
 wire _13188_;
 wire _13189_;
 wire _13190_;
 wire _13191_;
 wire _13192_;
 wire _13193_;
 wire _13194_;
 wire _13195_;
 wire _13196_;
 wire _13197_;
 wire _13198_;
 wire _13199_;
 wire _13200_;
 wire _13201_;
 wire _13202_;
 wire _13203_;
 wire _13204_;
 wire _13205_;
 wire _13206_;
 wire _13207_;
 wire _13208_;
 wire _13209_;
 wire _13210_;
 wire _13211_;
 wire _13212_;
 wire _13213_;
 wire _13214_;
 wire _13215_;
 wire _13216_;
 wire _13217_;
 wire _13218_;
 wire _13219_;
 wire _13220_;
 wire _13221_;
 wire _13222_;
 wire _13223_;
 wire _13224_;
 wire _13225_;
 wire _13226_;
 wire _13227_;
 wire _13228_;
 wire _13229_;
 wire _13230_;
 wire _13231_;
 wire _13232_;
 wire _13233_;
 wire _13234_;
 wire _13235_;
 wire _13236_;
 wire _13237_;
 wire _13238_;
 wire _13239_;
 wire _13240_;
 wire _13241_;
 wire _13242_;
 wire _13243_;
 wire _13244_;
 wire _13245_;
 wire _13246_;
 wire _13247_;
 wire _13248_;
 wire _13249_;
 wire _13250_;
 wire _13251_;
 wire _13252_;
 wire _13253_;
 wire _13254_;
 wire _13255_;
 wire _13256_;
 wire _13257_;
 wire _13258_;
 wire _13259_;
 wire _13260_;
 wire _13261_;
 wire _13262_;
 wire _13263_;
 wire _13264_;
 wire _13265_;
 wire _13266_;
 wire _13267_;
 wire _13268_;
 wire _13269_;
 wire _13270_;
 wire _13271_;
 wire _13272_;
 wire _13273_;
 wire _13274_;
 wire _13275_;
 wire _13276_;
 wire _13277_;
 wire _13278_;
 wire _13279_;
 wire _13280_;
 wire _13281_;
 wire _13282_;
 wire _13283_;
 wire _13284_;
 wire _13285_;
 wire _13286_;
 wire _13287_;
 wire _13288_;
 wire _13289_;
 wire _13290_;
 wire _13291_;
 wire _13292_;
 wire _13293_;
 wire _13294_;
 wire _13295_;
 wire _13296_;
 wire _13297_;
 wire _13298_;
 wire _13299_;
 wire _13300_;
 wire _13301_;
 wire _13302_;
 wire _13303_;
 wire _13304_;
 wire _13305_;
 wire _13306_;
 wire _13307_;
 wire _13308_;
 wire _13309_;
 wire _13310_;
 wire _13311_;
 wire _13312_;
 wire _13313_;
 wire _13314_;
 wire _13315_;
 wire _13316_;
 wire _13317_;
 wire _13318_;
 wire _13319_;
 wire _13320_;
 wire _13321_;
 wire _13322_;
 wire _13323_;
 wire _13324_;
 wire _13325_;
 wire _13326_;
 wire _13327_;
 wire _13328_;
 wire _13329_;
 wire _13330_;
 wire _13331_;
 wire _13332_;
 wire _13333_;
 wire _13334_;
 wire _13335_;
 wire _13336_;
 wire _13337_;
 wire _13338_;
 wire _13339_;
 wire _13340_;
 wire _13341_;
 wire _13342_;
 wire _13343_;
 wire _13344_;
 wire _13345_;
 wire _13346_;
 wire _13347_;
 wire _13348_;
 wire _13349_;
 wire _13350_;
 wire _13351_;
 wire _13352_;
 wire _13353_;
 wire _13354_;
 wire _13355_;
 wire _13356_;
 wire _13357_;
 wire _13358_;
 wire _13359_;
 wire _13360_;
 wire _13361_;
 wire _13362_;
 wire _13363_;
 wire _13364_;
 wire _13365_;
 wire _13366_;
 wire _13367_;
 wire _13368_;
 wire _13369_;
 wire _13370_;
 wire _13371_;
 wire _13372_;
 wire _13373_;
 wire _13374_;
 wire _13375_;
 wire _13376_;
 wire _13377_;
 wire _13378_;
 wire _13379_;
 wire _13380_;
 wire _13381_;
 wire _13382_;
 wire _13383_;
 wire _13384_;
 wire _13385_;
 wire _13386_;
 wire _13387_;
 wire _13388_;
 wire _13389_;
 wire _13390_;
 wire _13391_;
 wire _13392_;
 wire _13393_;
 wire _13394_;
 wire _13395_;
 wire _13396_;
 wire _13397_;
 wire _13398_;
 wire _13399_;
 wire _13400_;
 wire _13401_;
 wire _13403_;
 wire _13404_;
 wire _13405_;
 wire _13406_;
 wire _13407_;
 wire _13408_;
 wire _13409_;
 wire _13410_;
 wire _13411_;
 wire _13412_;
 wire _13413_;
 wire _13414_;
 wire _13415_;
 wire _13416_;
 wire _13417_;
 wire _13418_;
 wire _13419_;
 wire _13420_;
 wire _13421_;
 wire _13422_;
 wire _13423_;
 wire _13424_;
 wire _13425_;
 wire _13426_;
 wire _13427_;
 wire _13428_;
 wire _13429_;
 wire _13430_;
 wire _13431_;
 wire _13432_;
 wire _13433_;
 wire _13434_;
 wire _13435_;
 wire _13436_;
 wire _13437_;
 wire _13438_;
 wire _13439_;
 wire _13440_;
 wire _13441_;
 wire _13442_;
 wire _13443_;
 wire _13444_;
 wire _13445_;
 wire _13446_;
 wire _13447_;
 wire _13448_;
 wire _13449_;
 wire _13450_;
 wire _13451_;
 wire _13452_;
 wire _13453_;
 wire _13454_;
 wire _13455_;
 wire _13456_;
 wire _13457_;
 wire _13458_;
 wire _13459_;
 wire _13460_;
 wire _13461_;
 wire _13462_;
 wire _13463_;
 wire _13464_;
 wire _13465_;
 wire _13466_;
 wire _13467_;
 wire _13468_;
 wire _13469_;
 wire _13470_;
 wire _13471_;
 wire _13472_;
 wire _13473_;
 wire _13474_;
 wire _13475_;
 wire _13476_;
 wire _13477_;
 wire _13478_;
 wire _13479_;
 wire _13480_;
 wire _13481_;
 wire _13482_;
 wire _13483_;
 wire _13484_;
 wire _13485_;
 wire _13486_;
 wire _13487_;
 wire _13488_;
 wire _13489_;
 wire _13490_;
 wire _13491_;
 wire _13492_;
 wire _13493_;
 wire _13494_;
 wire _13495_;
 wire _13496_;
 wire _13497_;
 wire _13498_;
 wire _13499_;
 wire _13500_;
 wire _13501_;
 wire _13502_;
 wire _13503_;
 wire _13504_;
 wire _13505_;
 wire _13506_;
 wire _13507_;
 wire _13508_;
 wire _13509_;
 wire _13510_;
 wire _13511_;
 wire _13512_;
 wire _13513_;
 wire _13514_;
 wire _13515_;
 wire _13516_;
 wire _13517_;
 wire _13518_;
 wire _13519_;
 wire _13520_;
 wire _13521_;
 wire _13522_;
 wire _13523_;
 wire _13524_;
 wire _13525_;
 wire _13526_;
 wire _13527_;
 wire _13528_;
 wire _13529_;
 wire _13530_;
 wire _13531_;
 wire _13532_;
 wire _13533_;
 wire _13534_;
 wire _13535_;
 wire _13536_;
 wire _13537_;
 wire _13538_;
 wire _13539_;
 wire _13540_;
 wire _13541_;
 wire _13542_;
 wire _13543_;
 wire _13544_;
 wire _13545_;
 wire _13546_;
 wire _13547_;
 wire _13548_;
 wire _13549_;
 wire _13550_;
 wire _13551_;
 wire _13552_;
 wire _13553_;
 wire _13554_;
 wire _13555_;
 wire _13556_;
 wire _13557_;
 wire _13558_;
 wire _13559_;
 wire _13560_;
 wire _13561_;
 wire _13562_;
 wire _13563_;
 wire _13564_;
 wire _13565_;
 wire _13566_;
 wire _13567_;
 wire _13568_;
 wire _13569_;
 wire _13570_;
 wire _13571_;
 wire _13572_;
 wire _13573_;
 wire _13574_;
 wire _13575_;
 wire _13576_;
 wire _13577_;
 wire _13578_;
 wire _13579_;
 wire _13580_;
 wire _13581_;
 wire _13582_;
 wire _13583_;
 wire _13584_;
 wire _13585_;
 wire _13586_;
 wire _13587_;
 wire _13588_;
 wire _13589_;
 wire _13590_;
 wire _13591_;
 wire _13592_;
 wire _13593_;
 wire _13594_;
 wire _13595_;
 wire _13596_;
 wire _13597_;
 wire _13598_;
 wire _13599_;
 wire _13600_;
 wire _13601_;
 wire _13602_;
 wire _13603_;
 wire _13604_;
 wire _13605_;
 wire _13606_;
 wire _13607_;
 wire _13608_;
 wire _13609_;
 wire _13610_;
 wire _13611_;
 wire _13612_;
 wire _13613_;
 wire _13614_;
 wire _13615_;
 wire _13616_;
 wire _13617_;
 wire _13618_;
 wire _13619_;
 wire _13620_;
 wire _13621_;
 wire _13622_;
 wire _13623_;
 wire _13624_;
 wire _13625_;
 wire _13626_;
 wire _13627_;
 wire _13628_;
 wire _13629_;
 wire _13630_;
 wire _13631_;
 wire _13632_;
 wire _13633_;
 wire _13634_;
 wire _13635_;
 wire _13636_;
 wire _13637_;
 wire _13638_;
 wire _13639_;
 wire _13640_;
 wire _13641_;
 wire _13642_;
 wire _13643_;
 wire _13644_;
 wire _13645_;
 wire _13646_;
 wire _13647_;
 wire _13648_;
 wire _13649_;
 wire _13650_;
 wire _13651_;
 wire _13652_;
 wire _13653_;
 wire _13654_;
 wire _13655_;
 wire _13656_;
 wire _13657_;
 wire _13658_;
 wire _13659_;
 wire _13660_;
 wire _13661_;
 wire _13662_;
 wire _13663_;
 wire _13664_;
 wire _13665_;
 wire _13666_;
 wire _13667_;
 wire _13668_;
 wire _13669_;
 wire _13670_;
 wire _13671_;
 wire _13672_;
 wire _13673_;
 wire _13674_;
 wire _13675_;
 wire _13676_;
 wire _13677_;
 wire _13678_;
 wire _13679_;
 wire _13680_;
 wire _13681_;
 wire _13682_;
 wire _13683_;
 wire _13684_;
 wire _13685_;
 wire _13686_;
 wire _13687_;
 wire _13688_;
 wire _13689_;
 wire _13690_;
 wire _13691_;
 wire _13692_;
 wire _13693_;
 wire _13694_;
 wire _13695_;
 wire _13696_;
 wire _13697_;
 wire _13698_;
 wire _13699_;
 wire _13700_;
 wire _13701_;
 wire _13702_;
 wire _13703_;
 wire _13704_;
 wire _13705_;
 wire _13706_;
 wire _13707_;
 wire _13708_;
 wire _13709_;
 wire _13710_;
 wire _13711_;
 wire _13712_;
 wire _13713_;
 wire _13714_;
 wire _13715_;
 wire _13716_;
 wire _13717_;
 wire _13718_;
 wire _13719_;
 wire _13720_;
 wire _13721_;
 wire _13722_;
 wire _13723_;
 wire _13724_;
 wire _13725_;
 wire _13726_;
 wire _13727_;
 wire _13728_;
 wire _13729_;
 wire _13730_;
 wire _13731_;
 wire _13732_;
 wire _13733_;
 wire _13734_;
 wire _13735_;
 wire _13736_;
 wire _13737_;
 wire _13738_;
 wire _13739_;
 wire _13740_;
 wire _13741_;
 wire _13742_;
 wire _13743_;
 wire _13744_;
 wire _13745_;
 wire _13746_;
 wire _13747_;
 wire _13748_;
 wire _13749_;
 wire _13750_;
 wire _13751_;
 wire _13752_;
 wire _13753_;
 wire _13754_;
 wire _13755_;
 wire _13756_;
 wire _13757_;
 wire _13758_;
 wire _13759_;
 wire _13760_;
 wire _13761_;
 wire _13762_;
 wire _13763_;
 wire _13764_;
 wire _13765_;
 wire _13766_;
 wire _13767_;
 wire _13768_;
 wire _13769_;
 wire _13770_;
 wire _13771_;
 wire _13772_;
 wire _13773_;
 wire _13774_;
 wire _13775_;
 wire _13776_;
 wire _13777_;
 wire _13778_;
 wire _13779_;
 wire _13780_;
 wire _13781_;
 wire _13782_;
 wire _13783_;
 wire _13784_;
 wire _13785_;
 wire _13786_;
 wire _13787_;
 wire _13788_;
 wire _13789_;
 wire _13790_;
 wire _13791_;
 wire _13792_;
 wire _13793_;
 wire _13794_;
 wire _13795_;
 wire _13796_;
 wire _13797_;
 wire _13798_;
 wire _13799_;
 wire _13800_;
 wire _13801_;
 wire _13802_;
 wire _13803_;
 wire _13804_;
 wire _13805_;
 wire _13806_;
 wire _13807_;
 wire _13808_;
 wire _13809_;
 wire _13810_;
 wire _13811_;
 wire _13812_;
 wire _13813_;
 wire _13814_;
 wire _13815_;
 wire _13816_;
 wire _13817_;
 wire _13818_;
 wire _13819_;
 wire _13820_;
 wire _13821_;
 wire _13822_;
 wire _13823_;
 wire _13824_;
 wire _13825_;
 wire _13826_;
 wire _13827_;
 wire _13828_;
 wire _13829_;
 wire _13830_;
 wire _13831_;
 wire _13832_;
 wire _13833_;
 wire _13834_;
 wire _13835_;
 wire _13836_;
 wire _13837_;
 wire _13838_;
 wire _13839_;
 wire _13840_;
 wire _13841_;
 wire _13842_;
 wire _13843_;
 wire _13844_;
 wire _13845_;
 wire _13846_;
 wire _13847_;
 wire _13848_;
 wire _13849_;
 wire _13850_;
 wire _13851_;
 wire _13852_;
 wire _13853_;
 wire _13854_;
 wire _13855_;
 wire _13856_;
 wire _13857_;
 wire _13858_;
 wire _13859_;
 wire _13860_;
 wire _13861_;
 wire _13862_;
 wire _13863_;
 wire _13864_;
 wire _13865_;
 wire _13866_;
 wire _13867_;
 wire _13868_;
 wire _13869_;
 wire _13870_;
 wire _13871_;
 wire _13872_;
 wire _13873_;
 wire _13874_;
 wire _13875_;
 wire _13876_;
 wire _13877_;
 wire _13878_;
 wire _13879_;
 wire _13880_;
 wire _13881_;
 wire _13882_;
 wire _13883_;
 wire _13884_;
 wire _13885_;
 wire _13886_;
 wire _13887_;
 wire _13888_;
 wire _13889_;
 wire _13890_;
 wire _13891_;
 wire _13892_;
 wire _13893_;
 wire _13894_;
 wire _13895_;
 wire _13896_;
 wire _13897_;
 wire _13898_;
 wire _13899_;
 wire _13900_;
 wire _13901_;
 wire _13902_;
 wire _13903_;
 wire _13904_;
 wire _13905_;
 wire _13906_;
 wire _13907_;
 wire _13908_;
 wire _13909_;
 wire _13910_;
 wire _13911_;
 wire _13912_;
 wire _13913_;
 wire _13914_;
 wire _13915_;
 wire _13916_;
 wire _13917_;
 wire _13918_;
 wire _13919_;
 wire _13920_;
 wire _13921_;
 wire _13922_;
 wire _13923_;
 wire _13924_;
 wire _13925_;
 wire _13926_;
 wire _13927_;
 wire _13928_;
 wire _13929_;
 wire _13930_;
 wire _13931_;
 wire _13932_;
 wire _13933_;
 wire _13934_;
 wire _13935_;
 wire _13936_;
 wire _13937_;
 wire _13938_;
 wire _13939_;
 wire _13940_;
 wire _13941_;
 wire _13942_;
 wire _13943_;
 wire _13944_;
 wire _13945_;
 wire _13946_;
 wire _13947_;
 wire _13948_;
 wire _13949_;
 wire _13950_;
 wire _13951_;
 wire _13952_;
 wire _13953_;
 wire _13954_;
 wire _13955_;
 wire _13956_;
 wire _13957_;
 wire _13958_;
 wire _13959_;
 wire _13960_;
 wire _13961_;
 wire _13962_;
 wire _13963_;
 wire _13964_;
 wire _13965_;
 wire _13966_;
 wire _13967_;
 wire _13968_;
 wire _13969_;
 wire _13970_;
 wire _13971_;
 wire _13972_;
 wire _13973_;
 wire _13974_;
 wire _13975_;
 wire _13976_;
 wire _13977_;
 wire _13978_;
 wire _13979_;
 wire _13980_;
 wire _13981_;
 wire _13982_;
 wire _13983_;
 wire _13984_;
 wire _13985_;
 wire _13986_;
 wire _13987_;
 wire _13988_;
 wire _13989_;
 wire _13990_;
 wire _13991_;
 wire _13992_;
 wire _13993_;
 wire _13994_;
 wire _13995_;
 wire _13996_;
 wire _13997_;
 wire _13998_;
 wire _13999_;
 wire _14000_;
 wire _14001_;
 wire _14002_;
 wire _14003_;
 wire _14004_;
 wire _14005_;
 wire _14006_;
 wire _14007_;
 wire _14008_;
 wire _14009_;
 wire _14010_;
 wire _14011_;
 wire _14012_;
 wire _14013_;
 wire _14014_;
 wire _14015_;
 wire _14016_;
 wire _14017_;
 wire _14018_;
 wire _14019_;
 wire _14020_;
 wire _14021_;
 wire _14022_;
 wire _14023_;
 wire _14024_;
 wire _14025_;
 wire _14026_;
 wire _14027_;
 wire _14028_;
 wire _14029_;
 wire _14030_;
 wire _14031_;
 wire _14032_;
 wire _14033_;
 wire _14034_;
 wire _14035_;
 wire _14036_;
 wire _14037_;
 wire _14038_;
 wire _14039_;
 wire _14040_;
 wire _14041_;
 wire _14042_;
 wire _14043_;
 wire _14044_;
 wire _14045_;
 wire _14046_;
 wire _14047_;
 wire _14048_;
 wire _14049_;
 wire _14050_;
 wire _14051_;
 wire _14052_;
 wire _14053_;
 wire _14054_;
 wire _14055_;
 wire _14056_;
 wire _14057_;
 wire _14058_;
 wire _14059_;
 wire _14060_;
 wire _14061_;
 wire _14062_;
 wire _14063_;
 wire _14064_;
 wire _14065_;
 wire _14066_;
 wire _14067_;
 wire _14068_;
 wire _14069_;
 wire _14070_;
 wire _14071_;
 wire _14072_;
 wire _14073_;
 wire _14074_;
 wire _14075_;
 wire _14076_;
 wire _14077_;
 wire _14078_;
 wire _14079_;
 wire _14080_;
 wire _14081_;
 wire _14082_;
 wire _14083_;
 wire _14084_;
 wire _14085_;
 wire _14086_;
 wire _14087_;
 wire _14088_;
 wire _14089_;
 wire _14090_;
 wire _14091_;
 wire _14092_;
 wire _14093_;
 wire _14094_;
 wire _14095_;
 wire _14096_;
 wire _14097_;
 wire _14098_;
 wire _14099_;
 wire _14100_;
 wire _14101_;
 wire _14102_;
 wire _14103_;
 wire _14104_;
 wire _14105_;
 wire _14106_;
 wire _14107_;
 wire _14108_;
 wire _14109_;
 wire _14110_;
 wire _14111_;
 wire _14112_;
 wire _14113_;
 wire _14114_;
 wire _14115_;
 wire _14116_;
 wire _14117_;
 wire _14118_;
 wire _14119_;
 wire _14120_;
 wire _14121_;
 wire _14122_;
 wire _14123_;
 wire _14124_;
 wire _14125_;
 wire _14126_;
 wire _14127_;
 wire _14128_;
 wire _14129_;
 wire _14130_;
 wire _14131_;
 wire _14132_;
 wire _14133_;
 wire _14134_;
 wire _14135_;
 wire _14136_;
 wire _14137_;
 wire _14138_;
 wire _14139_;
 wire _14140_;
 wire _14141_;
 wire _14142_;
 wire _14143_;
 wire _14144_;
 wire _14145_;
 wire _14146_;
 wire _14147_;
 wire _14148_;
 wire _14149_;
 wire _14150_;
 wire _14151_;
 wire _14152_;
 wire _14153_;
 wire _14154_;
 wire _14155_;
 wire _14156_;
 wire _14157_;
 wire _14158_;
 wire _14159_;
 wire _14160_;
 wire _14161_;
 wire _14162_;
 wire _14163_;
 wire _14164_;
 wire _14165_;
 wire _14166_;
 wire _14167_;
 wire _14168_;
 wire _14169_;
 wire _14170_;
 wire _14171_;
 wire _14172_;
 wire _14173_;
 wire _14174_;
 wire _14175_;
 wire _14176_;
 wire _14177_;
 wire _14178_;
 wire _14179_;
 wire _14180_;
 wire _14181_;
 wire _14182_;
 wire _14183_;
 wire _14184_;
 wire _14185_;
 wire _14186_;
 wire _14187_;
 wire _14188_;
 wire _14189_;
 wire _14190_;
 wire _14191_;
 wire _14192_;
 wire _14193_;
 wire _14194_;
 wire _14195_;
 wire _14196_;
 wire _14197_;
 wire _14198_;
 wire _14199_;
 wire _14200_;
 wire _14201_;
 wire _14202_;
 wire _14203_;
 wire _14204_;
 wire _14205_;
 wire _14206_;
 wire _14207_;
 wire _14208_;
 wire _14209_;
 wire _14210_;
 wire _14211_;
 wire _14212_;
 wire _14213_;
 wire _14214_;
 wire _14215_;
 wire _14216_;
 wire _14217_;
 wire _14218_;
 wire _14219_;
 wire _14220_;
 wire _14221_;
 wire _14222_;
 wire _14223_;
 wire _14224_;
 wire _14225_;
 wire _14226_;
 wire _14227_;
 wire _14228_;
 wire _14229_;
 wire _14230_;
 wire _14231_;
 wire _14232_;
 wire _14233_;
 wire _14234_;
 wire _14235_;
 wire _14236_;
 wire _14237_;
 wire _14238_;
 wire _14239_;
 wire _14240_;
 wire _14241_;
 wire _14242_;
 wire _14243_;
 wire _14244_;
 wire _14245_;
 wire _14246_;
 wire _14247_;
 wire _14248_;
 wire _14249_;
 wire _14250_;
 wire _14251_;
 wire _14252_;
 wire _14253_;
 wire _14254_;
 wire _14255_;
 wire _14256_;
 wire _14257_;
 wire _14258_;
 wire _14259_;
 wire _14260_;
 wire _14261_;
 wire _14262_;
 wire _14263_;
 wire _14264_;
 wire _14265_;
 wire _14266_;
 wire _14267_;
 wire _14268_;
 wire _14269_;
 wire _14270_;
 wire _14271_;
 wire _14272_;
 wire _14273_;
 wire _14274_;
 wire _14275_;
 wire _14276_;
 wire _14277_;
 wire _14278_;
 wire _14279_;
 wire _14280_;
 wire _14281_;
 wire _14282_;
 wire _14283_;
 wire _14284_;
 wire _14285_;
 wire _14286_;
 wire _14287_;
 wire _14288_;
 wire _14289_;
 wire _14290_;
 wire _14291_;
 wire _14292_;
 wire _14293_;
 wire _14294_;
 wire _14295_;
 wire _14296_;
 wire _14297_;
 wire _14298_;
 wire _14299_;
 wire _14301_;
 wire _14302_;
 wire _14303_;
 wire _14304_;
 wire _14305_;
 wire _14306_;
 wire _14307_;
 wire _14308_;
 wire _14309_;
 wire _14310_;
 wire _14311_;
 wire _14312_;
 wire _14313_;
 wire _14314_;
 wire _14315_;
 wire _14316_;
 wire _14317_;
 wire _14318_;
 wire _14319_;
 wire _14320_;
 wire _14321_;
 wire _14322_;
 wire _14323_;
 wire _14324_;
 wire _14325_;
 wire _14326_;
 wire _14327_;
 wire _14328_;
 wire _14329_;
 wire _14330_;
 wire _14331_;
 wire _14332_;
 wire _14333_;
 wire _14334_;
 wire _14335_;
 wire _14336_;
 wire _14337_;
 wire _14338_;
 wire _14339_;
 wire _14340_;
 wire _14341_;
 wire _14342_;
 wire _14343_;
 wire _14344_;
 wire _14345_;
 wire _14346_;
 wire _14347_;
 wire _14348_;
 wire _14349_;
 wire _14350_;
 wire _14351_;
 wire _14352_;
 wire _14353_;
 wire _14354_;
 wire _14355_;
 wire _14356_;
 wire _14357_;
 wire _14358_;
 wire _14359_;
 wire _14360_;
 wire _14361_;
 wire _14362_;
 wire _14363_;
 wire _14364_;
 wire _14365_;
 wire _14366_;
 wire _14367_;
 wire _14368_;
 wire _14369_;
 wire _14370_;
 wire _14371_;
 wire _14372_;
 wire _14373_;
 wire _14374_;
 wire _14375_;
 wire _14376_;
 wire _14377_;
 wire _14378_;
 wire _14379_;
 wire _14380_;
 wire _14381_;
 wire _14382_;
 wire _14383_;
 wire _14384_;
 wire _14385_;
 wire _14386_;
 wire _14387_;
 wire _14388_;
 wire _14389_;
 wire _14390_;
 wire _14391_;
 wire _14392_;
 wire _14393_;
 wire _14394_;
 wire _14395_;
 wire _14396_;
 wire _14397_;
 wire _14398_;
 wire _14399_;
 wire _14400_;
 wire _14401_;
 wire _14402_;
 wire _14403_;
 wire _14404_;
 wire _14405_;
 wire _14406_;
 wire _14407_;
 wire _14408_;
 wire _14409_;
 wire _14410_;
 wire _14411_;
 wire _14412_;
 wire _14413_;
 wire _14414_;
 wire _14415_;
 wire _14416_;
 wire _14417_;
 wire _14418_;
 wire _14419_;
 wire _14420_;
 wire _14421_;
 wire _14422_;
 wire _14423_;
 wire _14424_;
 wire _14425_;
 wire _14426_;
 wire _14427_;
 wire _14428_;
 wire _14429_;
 wire _14430_;
 wire _14431_;
 wire _14432_;
 wire _14433_;
 wire _14434_;
 wire _14435_;
 wire _14436_;
 wire _14437_;
 wire _14438_;
 wire _14439_;
 wire _14440_;
 wire _14441_;
 wire _14442_;
 wire _14443_;
 wire _14444_;
 wire _14445_;
 wire _14446_;
 wire _14447_;
 wire _14448_;
 wire _14449_;
 wire _14450_;
 wire _14451_;
 wire _14452_;
 wire _14453_;
 wire _14454_;
 wire _14455_;
 wire _14456_;
 wire _14457_;
 wire _14458_;
 wire _14459_;
 wire _14460_;
 wire _14461_;
 wire _14462_;
 wire _14463_;
 wire _14464_;
 wire _14465_;
 wire _14466_;
 wire _14467_;
 wire _14468_;
 wire _14469_;
 wire _14470_;
 wire _14471_;
 wire _14472_;
 wire _14473_;
 wire _14474_;
 wire _14475_;
 wire _14476_;
 wire _14477_;
 wire _14478_;
 wire _14479_;
 wire _14480_;
 wire _14481_;
 wire _14482_;
 wire _14483_;
 wire _14484_;
 wire _14485_;
 wire _14486_;
 wire _14487_;
 wire _14488_;
 wire _14489_;
 wire _14490_;
 wire _14491_;
 wire _14492_;
 wire _14493_;
 wire _14494_;
 wire _14495_;
 wire _14496_;
 wire _14497_;
 wire _14498_;
 wire _14499_;
 wire _14500_;
 wire _14501_;
 wire _14502_;
 wire _14503_;
 wire _14504_;
 wire _14505_;
 wire _14506_;
 wire _14507_;
 wire _14508_;
 wire _14509_;
 wire _14510_;
 wire _14511_;
 wire _14512_;
 wire _14513_;
 wire _14514_;
 wire _14515_;
 wire _14516_;
 wire _14517_;
 wire _14518_;
 wire _14519_;
 wire _14520_;
 wire _14521_;
 wire _14522_;
 wire _14523_;
 wire _14524_;
 wire _14525_;
 wire _14526_;
 wire _14527_;
 wire _14528_;
 wire _14529_;
 wire _14530_;
 wire _14531_;
 wire _14532_;
 wire _14533_;
 wire _14534_;
 wire _14535_;
 wire _14536_;
 wire _14537_;
 wire _14538_;
 wire _14539_;
 wire _14540_;
 wire _14541_;
 wire _14542_;
 wire _14543_;
 wire _14544_;
 wire _14545_;
 wire _14546_;
 wire _14547_;
 wire _14548_;
 wire _14549_;
 wire _14550_;
 wire _14551_;
 wire _14552_;
 wire _14553_;
 wire _14554_;
 wire _14555_;
 wire _14556_;
 wire _14557_;
 wire _14558_;
 wire _14559_;
 wire _14560_;
 wire _14561_;
 wire _14562_;
 wire _14563_;
 wire _14564_;
 wire _14565_;
 wire _14566_;
 wire _14567_;
 wire _14568_;
 wire _14569_;
 wire _14570_;
 wire _14571_;
 wire _14572_;
 wire _14573_;
 wire _14574_;
 wire _14575_;
 wire _14576_;
 wire _14577_;
 wire _14578_;
 wire _14579_;
 wire _14580_;
 wire _14581_;
 wire _14582_;
 wire _14583_;
 wire _14584_;
 wire _14585_;
 wire _14586_;
 wire _14587_;
 wire _14588_;
 wire _14589_;
 wire _14590_;
 wire _14591_;
 wire _14592_;
 wire _14593_;
 wire _14594_;
 wire _14595_;
 wire _14596_;
 wire _14597_;
 wire _14598_;
 wire _14599_;
 wire _14600_;
 wire _14601_;
 wire _14602_;
 wire _14603_;
 wire _14604_;
 wire _14605_;
 wire _14606_;
 wire _14607_;
 wire _14608_;
 wire _14609_;
 wire _14610_;
 wire _14611_;
 wire _14612_;
 wire _14613_;
 wire _14614_;
 wire _14615_;
 wire _14616_;
 wire _14617_;
 wire _14618_;
 wire _14619_;
 wire _14620_;
 wire _14621_;
 wire _14622_;
 wire _14623_;
 wire _14624_;
 wire _14625_;
 wire _14626_;
 wire _14627_;
 wire _14628_;
 wire _14629_;
 wire _14630_;
 wire _14631_;
 wire _14632_;
 wire _14633_;
 wire _14634_;
 wire _14635_;
 wire _14636_;
 wire _14637_;
 wire _14638_;
 wire _14639_;
 wire _14640_;
 wire _14641_;
 wire _14642_;
 wire _14643_;
 wire _14644_;
 wire _14645_;
 wire _14646_;
 wire _14647_;
 wire _14648_;
 wire _14649_;
 wire _14650_;
 wire _14651_;
 wire _14652_;
 wire _14653_;
 wire _14654_;
 wire _14655_;
 wire _14656_;
 wire _14657_;
 wire _14658_;
 wire _14659_;
 wire _14660_;
 wire _14661_;
 wire _14662_;
 wire _14663_;
 wire _14664_;
 wire _14665_;
 wire _14666_;
 wire _14667_;
 wire _14668_;
 wire _14669_;
 wire _14670_;
 wire _14671_;
 wire _14672_;
 wire _14673_;
 wire _14674_;
 wire _14675_;
 wire _14676_;
 wire _14677_;
 wire _14678_;
 wire _14679_;
 wire _14680_;
 wire _14681_;
 wire _14682_;
 wire _14683_;
 wire _14684_;
 wire _14685_;
 wire _14686_;
 wire _14687_;
 wire _14688_;
 wire _14689_;
 wire _14690_;
 wire _14691_;
 wire _14692_;
 wire _14693_;
 wire _14694_;
 wire _14695_;
 wire _14696_;
 wire _14697_;
 wire _14698_;
 wire _14699_;
 wire _14700_;
 wire _14701_;
 wire _14702_;
 wire _14703_;
 wire _14704_;
 wire _14705_;
 wire _14706_;
 wire _14707_;
 wire _14708_;
 wire _14709_;
 wire _14710_;
 wire _14711_;
 wire _14712_;
 wire _14713_;
 wire _14714_;
 wire _14715_;
 wire _14716_;
 wire _14717_;
 wire _14718_;
 wire _14719_;
 wire _14720_;
 wire _14721_;
 wire _14722_;
 wire _14723_;
 wire _14724_;
 wire _14725_;
 wire _14726_;
 wire _14727_;
 wire _14728_;
 wire _14729_;
 wire _14730_;
 wire _14731_;
 wire _14732_;
 wire _14733_;
 wire _14734_;
 wire _14735_;
 wire _14736_;
 wire _14737_;
 wire _14738_;
 wire _14739_;
 wire _14740_;
 wire _14741_;
 wire _14742_;
 wire _14743_;
 wire _14744_;
 wire _14745_;
 wire _14746_;
 wire _14747_;
 wire _14748_;
 wire _14749_;
 wire _14750_;
 wire _14751_;
 wire _14752_;
 wire _14753_;
 wire _14754_;
 wire _14755_;
 wire _14756_;
 wire _14757_;
 wire _14758_;
 wire _14759_;
 wire _14760_;
 wire _14761_;
 wire _14762_;
 wire _14763_;
 wire _14764_;
 wire _14765_;
 wire _14766_;
 wire _14767_;
 wire _14768_;
 wire _14769_;
 wire _14770_;
 wire _14771_;
 wire _14772_;
 wire _14773_;
 wire _14774_;
 wire _14775_;
 wire _14776_;
 wire _14777_;
 wire _14778_;
 wire _14779_;
 wire _14780_;
 wire _14781_;
 wire _14782_;
 wire _14783_;
 wire _14784_;
 wire _14785_;
 wire _14786_;
 wire _14787_;
 wire _14788_;
 wire _14789_;
 wire _14790_;
 wire _14791_;
 wire _14792_;
 wire _14793_;
 wire _14794_;
 wire _14795_;
 wire _14796_;
 wire _14797_;
 wire _14798_;
 wire _14799_;
 wire _14800_;
 wire _14801_;
 wire _14802_;
 wire _14803_;
 wire _14804_;
 wire _14805_;
 wire _14806_;
 wire _14807_;
 wire _14808_;
 wire _14809_;
 wire _14810_;
 wire _14811_;
 wire _14812_;
 wire _14813_;
 wire _14814_;
 wire _14815_;
 wire _14816_;
 wire _14817_;
 wire _14818_;
 wire _14819_;
 wire _14820_;
 wire _14821_;
 wire _14822_;
 wire _14823_;
 wire _14824_;
 wire _14825_;
 wire _14826_;
 wire _14827_;
 wire _14828_;
 wire _14829_;
 wire _14830_;
 wire _14831_;
 wire _14832_;
 wire _14833_;
 wire _14834_;
 wire _14835_;
 wire _14836_;
 wire _14837_;
 wire _14838_;
 wire _14839_;
 wire _14840_;
 wire _14841_;
 wire _14842_;
 wire _14843_;
 wire _14844_;
 wire _14845_;
 wire _14846_;
 wire _14847_;
 wire _14848_;
 wire _14849_;
 wire _14850_;
 wire _14851_;
 wire _14852_;
 wire _14853_;
 wire _14854_;
 wire _14855_;
 wire _14856_;
 wire _14857_;
 wire _14858_;
 wire _14859_;
 wire _14860_;
 wire _14861_;
 wire _14862_;
 wire _14863_;
 wire _14864_;
 wire _14865_;
 wire _14866_;
 wire _14867_;
 wire _14868_;
 wire _14869_;
 wire _14870_;
 wire _14871_;
 wire _14872_;
 wire _14873_;
 wire _14874_;
 wire _14875_;
 wire _14876_;
 wire _14877_;
 wire _14878_;
 wire _14879_;
 wire _14880_;
 wire _14881_;
 wire _14882_;
 wire _14883_;
 wire _14884_;
 wire _14885_;
 wire _14886_;
 wire _14887_;
 wire _14888_;
 wire _14889_;
 wire _14890_;
 wire _14891_;
 wire _14892_;
 wire _14893_;
 wire _14894_;
 wire _14895_;
 wire _14896_;
 wire _14897_;
 wire _14898_;
 wire _14899_;
 wire _14900_;
 wire _14901_;
 wire _14902_;
 wire _14903_;
 wire _14904_;
 wire _14905_;
 wire _14906_;
 wire _14907_;
 wire _14908_;
 wire _14909_;
 wire _14910_;
 wire _14911_;
 wire _14912_;
 wire _14913_;
 wire _14914_;
 wire _14915_;
 wire _14916_;
 wire _14917_;
 wire _14918_;
 wire _14919_;
 wire _14920_;
 wire _14921_;
 wire _14922_;
 wire _14923_;
 wire _14924_;
 wire _14925_;
 wire _14926_;
 wire _14927_;
 wire _14928_;
 wire _14929_;
 wire _14930_;
 wire _14931_;
 wire _14932_;
 wire _14933_;
 wire _14934_;
 wire _14935_;
 wire _14936_;
 wire _14937_;
 wire _14938_;
 wire _14939_;
 wire _14940_;
 wire _14941_;
 wire _14942_;
 wire _14943_;
 wire _14944_;
 wire _14945_;
 wire _14946_;
 wire _14947_;
 wire _14948_;
 wire _14949_;
 wire _14950_;
 wire _14951_;
 wire _14952_;
 wire _14953_;
 wire _14954_;
 wire _14955_;
 wire _14956_;
 wire _14957_;
 wire _14958_;
 wire _14959_;
 wire _14960_;
 wire _14961_;
 wire _14962_;
 wire _14963_;
 wire _14964_;
 wire _14965_;
 wire _14966_;
 wire _14967_;
 wire _14968_;
 wire _14969_;
 wire _14970_;
 wire _14971_;
 wire _14972_;
 wire _14973_;
 wire _14974_;
 wire _14975_;
 wire _14976_;
 wire _14977_;
 wire _14978_;
 wire _14979_;
 wire _14980_;
 wire _14981_;
 wire _14982_;
 wire _14983_;
 wire _14984_;
 wire _14985_;
 wire _14986_;
 wire _14987_;
 wire _14988_;
 wire _14989_;
 wire _14990_;
 wire _14991_;
 wire _14992_;
 wire _14993_;
 wire _14994_;
 wire _14995_;
 wire _14996_;
 wire _14997_;
 wire _14998_;
 wire _14999_;
 wire _15000_;
 wire _15001_;
 wire _15002_;
 wire _15003_;
 wire _15004_;
 wire _15005_;
 wire _15006_;
 wire _15007_;
 wire _15008_;
 wire _15009_;
 wire _15010_;
 wire _15011_;
 wire _15012_;
 wire _15013_;
 wire _15014_;
 wire _15015_;
 wire _15016_;
 wire _15017_;
 wire _15018_;
 wire _15019_;
 wire _15020_;
 wire _15021_;
 wire _15022_;
 wire _15023_;
 wire _15024_;
 wire _15025_;
 wire _15026_;
 wire _15027_;
 wire _15028_;
 wire _15029_;
 wire _15030_;
 wire _15031_;
 wire _15032_;
 wire _15033_;
 wire _15034_;
 wire _15035_;
 wire _15036_;
 wire _15037_;
 wire _15038_;
 wire _15039_;
 wire _15040_;
 wire _15041_;
 wire _15042_;
 wire _15043_;
 wire _15044_;
 wire _15045_;
 wire _15046_;
 wire _15047_;
 wire _15048_;
 wire _15049_;
 wire _15050_;
 wire _15051_;
 wire _15052_;
 wire _15053_;
 wire _15054_;
 wire _15055_;
 wire _15056_;
 wire _15057_;
 wire _15058_;
 wire _15059_;
 wire _15060_;
 wire _15061_;
 wire _15062_;
 wire _15063_;
 wire _15064_;
 wire _15065_;
 wire _15066_;
 wire _15067_;
 wire _15068_;
 wire _15069_;
 wire _15070_;
 wire _15071_;
 wire _15072_;
 wire _15073_;
 wire _15074_;
 wire _15075_;
 wire _15076_;
 wire _15077_;
 wire _15078_;
 wire _15079_;
 wire _15080_;
 wire _15081_;
 wire _15082_;
 wire _15083_;
 wire _15084_;
 wire _15085_;
 wire _15086_;
 wire _15087_;
 wire _15088_;
 wire _15089_;
 wire _15090_;
 wire _15091_;
 wire _15092_;
 wire _15093_;
 wire _15094_;
 wire _15095_;
 wire _15096_;
 wire _15097_;
 wire _15098_;
 wire _15099_;
 wire _15100_;
 wire _15101_;
 wire _15102_;
 wire _15103_;
 wire _15104_;
 wire _15105_;
 wire _15106_;
 wire _15107_;
 wire _15108_;
 wire _15109_;
 wire _15110_;
 wire _15111_;
 wire _15112_;
 wire _15113_;
 wire _15114_;
 wire _15115_;
 wire _15116_;
 wire _15117_;
 wire _15118_;
 wire _15119_;
 wire _15120_;
 wire _15121_;
 wire _15122_;
 wire _15123_;
 wire _15124_;
 wire _15125_;
 wire _15126_;
 wire _15127_;
 wire _15128_;
 wire _15129_;
 wire _15130_;
 wire _15131_;
 wire _15133_;
 wire _15134_;
 wire _15135_;
 wire _15136_;
 wire _15137_;
 wire _15138_;
 wire _15139_;
 wire _15140_;
 wire _15141_;
 wire _15142_;
 wire _15143_;
 wire _15144_;
 wire _15145_;
 wire _15146_;
 wire _15147_;
 wire _15148_;
 wire _15149_;
 wire _15150_;
 wire _15151_;
 wire _15152_;
 wire _15153_;
 wire _15154_;
 wire _15155_;
 wire _15156_;
 wire _15157_;
 wire _15158_;
 wire _15159_;
 wire _15160_;
 wire _15161_;
 wire _15162_;
 wire _15163_;
 wire _15164_;
 wire _15165_;
 wire _15166_;
 wire _15167_;
 wire _15168_;
 wire _15169_;
 wire _15170_;
 wire _15171_;
 wire _15172_;
 wire _15173_;
 wire _15174_;
 wire _15175_;
 wire _15176_;
 wire _15177_;
 wire _15178_;
 wire _15179_;
 wire _15180_;
 wire _15181_;
 wire _15182_;
 wire _15183_;
 wire _15184_;
 wire _15185_;
 wire _15186_;
 wire _15187_;
 wire _15188_;
 wire _15189_;
 wire _15190_;
 wire _15191_;
 wire _15192_;
 wire _15193_;
 wire _15194_;
 wire _15195_;
 wire _15196_;
 wire _15197_;
 wire _15198_;
 wire _15199_;
 wire _15200_;
 wire _15201_;
 wire _15202_;
 wire _15203_;
 wire _15204_;
 wire _15205_;
 wire _15206_;
 wire _15207_;
 wire _15208_;
 wire _15209_;
 wire _15210_;
 wire _15211_;
 wire _15212_;
 wire _15213_;
 wire _15214_;
 wire _15215_;
 wire _15216_;
 wire _15217_;
 wire _15218_;
 wire _15219_;
 wire _15220_;
 wire _15221_;
 wire _15222_;
 wire _15223_;
 wire _15224_;
 wire _15225_;
 wire _15226_;
 wire _15227_;
 wire _15228_;
 wire _15229_;
 wire _15230_;
 wire _15231_;
 wire _15232_;
 wire _15233_;
 wire _15234_;
 wire _15235_;
 wire _15236_;
 wire _15237_;
 wire _15238_;
 wire _15239_;
 wire _15240_;
 wire _15241_;
 wire _15242_;
 wire _15243_;
 wire _15244_;
 wire _15245_;
 wire _15246_;
 wire _15247_;
 wire _15248_;
 wire _15249_;
 wire _15250_;
 wire _15251_;
 wire _15252_;
 wire _15253_;
 wire _15254_;
 wire _15255_;
 wire _15256_;
 wire _15257_;
 wire _15258_;
 wire _15259_;
 wire _15260_;
 wire _15261_;
 wire _15262_;
 wire _15263_;
 wire _15264_;
 wire _15265_;
 wire _15266_;
 wire _15267_;
 wire _15268_;
 wire _15269_;
 wire _15270_;
 wire _15271_;
 wire _15272_;
 wire _15273_;
 wire _15274_;
 wire _15275_;
 wire _15276_;
 wire _15277_;
 wire _15278_;
 wire _15279_;
 wire _15280_;
 wire _15281_;
 wire _15282_;
 wire _15283_;
 wire _15284_;
 wire _15285_;
 wire _15286_;
 wire _15287_;
 wire _15288_;
 wire _15289_;
 wire _15290_;
 wire _15291_;
 wire _15292_;
 wire _15293_;
 wire _15294_;
 wire _15295_;
 wire _15296_;
 wire _15297_;
 wire _15298_;
 wire _15299_;
 wire _15300_;
 wire _15301_;
 wire _15302_;
 wire _15303_;
 wire _15304_;
 wire _15305_;
 wire _15306_;
 wire _15307_;
 wire _15308_;
 wire _15309_;
 wire _15310_;
 wire _15311_;
 wire _15312_;
 wire _15313_;
 wire _15314_;
 wire _15315_;
 wire _15316_;
 wire _15317_;
 wire _15318_;
 wire _15319_;
 wire _15320_;
 wire _15321_;
 wire _15322_;
 wire _15323_;
 wire _15324_;
 wire _15325_;
 wire _15326_;
 wire _15327_;
 wire _15328_;
 wire _15329_;
 wire _15330_;
 wire _15331_;
 wire _15332_;
 wire _15333_;
 wire _15334_;
 wire _15335_;
 wire _15336_;
 wire _15337_;
 wire _15338_;
 wire _15339_;
 wire _15340_;
 wire _15341_;
 wire _15342_;
 wire _15343_;
 wire _15344_;
 wire _15345_;
 wire _15346_;
 wire _15347_;
 wire _15348_;
 wire _15349_;
 wire _15350_;
 wire _15351_;
 wire _15352_;
 wire _15353_;
 wire _15354_;
 wire _15355_;
 wire _15356_;
 wire _15357_;
 wire _15358_;
 wire _15359_;
 wire _15360_;
 wire _15361_;
 wire _15362_;
 wire _15363_;
 wire _15364_;
 wire _15365_;
 wire _15366_;
 wire _15367_;
 wire _15368_;
 wire _15369_;
 wire _15370_;
 wire _15371_;
 wire _15372_;
 wire _15373_;
 wire _15374_;
 wire _15375_;
 wire _15376_;
 wire _15377_;
 wire _15378_;
 wire _15379_;
 wire _15380_;
 wire _15381_;
 wire _15382_;
 wire _15383_;
 wire _15384_;
 wire _15385_;
 wire _15386_;
 wire _15387_;
 wire _15388_;
 wire _15389_;
 wire _15390_;
 wire _15391_;
 wire _15392_;
 wire _15393_;
 wire _15394_;
 wire _15395_;
 wire _15396_;
 wire _15397_;
 wire _15398_;
 wire _15399_;
 wire _15400_;
 wire _15401_;
 wire _15402_;
 wire _15403_;
 wire _15404_;
 wire _15405_;
 wire _15406_;
 wire _15407_;
 wire _15408_;
 wire _15409_;
 wire _15410_;
 wire _15411_;
 wire _15412_;
 wire _15413_;
 wire _15414_;
 wire _15415_;
 wire _15416_;
 wire _15417_;
 wire _15418_;
 wire _15419_;
 wire _15420_;
 wire _15421_;
 wire _15422_;
 wire _15423_;
 wire _15424_;
 wire _15425_;
 wire _15426_;
 wire _15427_;
 wire _15428_;
 wire _15429_;
 wire _15430_;
 wire _15431_;
 wire _15432_;
 wire _15433_;
 wire _15434_;
 wire _15435_;
 wire _15436_;
 wire _15437_;
 wire _15438_;
 wire _15439_;
 wire _15440_;
 wire _15441_;
 wire _15442_;
 wire _15443_;
 wire _15444_;
 wire _15445_;
 wire _15446_;
 wire _15447_;
 wire _15448_;
 wire _15449_;
 wire _15450_;
 wire _15451_;
 wire _15452_;
 wire _15453_;
 wire _15454_;
 wire _15455_;
 wire _15456_;
 wire _15457_;
 wire _15458_;
 wire _15459_;
 wire _15460_;
 wire _15461_;
 wire _15462_;
 wire _15463_;
 wire _15464_;
 wire _15465_;
 wire _15466_;
 wire _15467_;
 wire _15468_;
 wire _15469_;
 wire _15470_;
 wire _15471_;
 wire _15472_;
 wire _15473_;
 wire _15474_;
 wire _15475_;
 wire _15476_;
 wire _15477_;
 wire _15478_;
 wire _15479_;
 wire _15480_;
 wire _15481_;
 wire _15482_;
 wire _15483_;
 wire _15484_;
 wire _15485_;
 wire _15486_;
 wire _15487_;
 wire _15488_;
 wire _15489_;
 wire _15490_;
 wire _15491_;
 wire _15492_;
 wire _15493_;
 wire _15494_;
 wire _15495_;
 wire _15496_;
 wire _15497_;
 wire _15498_;
 wire _15499_;
 wire _15500_;
 wire _15501_;
 wire _15502_;
 wire _15503_;
 wire _15504_;
 wire _15505_;
 wire _15506_;
 wire _15507_;
 wire _15508_;
 wire _15509_;
 wire _15510_;
 wire _15511_;
 wire _15512_;
 wire _15513_;
 wire _15514_;
 wire _15515_;
 wire _15516_;
 wire _15517_;
 wire _15518_;
 wire _15519_;
 wire _15520_;
 wire _15521_;
 wire _15522_;
 wire _15523_;
 wire _15524_;
 wire _15525_;
 wire _15526_;
 wire _15527_;
 wire _15528_;
 wire _15529_;
 wire _15530_;
 wire _15531_;
 wire _15532_;
 wire _15533_;
 wire _15534_;
 wire _15535_;
 wire _15536_;
 wire _15537_;
 wire _15538_;
 wire _15539_;
 wire _15540_;
 wire _15541_;
 wire _15542_;
 wire _15543_;
 wire _15544_;
 wire _15545_;
 wire _15546_;
 wire _15547_;
 wire _15548_;
 wire _15549_;
 wire _15550_;
 wire _15551_;
 wire _15552_;
 wire _15553_;
 wire _15554_;
 wire _15555_;
 wire _15556_;
 wire _15557_;
 wire _15558_;
 wire _15559_;
 wire _15560_;
 wire _15561_;
 wire _15562_;
 wire _15563_;
 wire _15564_;
 wire _15565_;
 wire _15566_;
 wire _15567_;
 wire _15568_;
 wire _15570_;
 wire _15571_;
 wire _15572_;
 wire _15573_;
 wire _15574_;
 wire _15575_;
 wire _15576_;
 wire _15577_;
 wire _15578_;
 wire _15579_;
 wire _15580_;
 wire _15581_;
 wire _15582_;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire core_busy_q;
 wire \core_clock_gate_i.en_latch ;
 wire net439;
 wire \cs_registers_i.csr_mstatus_mie_o ;
 wire \cs_registers_i.csr_mstatus_tw_o ;
 wire \cs_registers_i.debug_ebreakm_o ;
 wire \cs_registers_i.debug_ebreaku_o ;
 wire \cs_registers_i.debug_mode_i ;
 wire \cs_registers_i.debug_single_step_o ;
 wire \cs_registers_i.nmi_mode_i ;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net474;
 wire net348;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net349;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.div_by_zero_q ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.div_valid ;
 wire net350;
 wire fetch_enable_q;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire \id_stage_i.branch_set ;
 wire \id_stage_i.controller_i.controller_run_o ;
 wire \id_stage_i.controller_i.exc_req_q ;
 wire \id_stage_i.controller_i.illegal_insn_q ;
 wire \id_stage_i.controller_i.instr_fetch_err_i ;
 wire \id_stage_i.controller_i.instr_fetch_err_plus2_i ;
 wire \id_stage_i.controller_i.instr_is_compressed_i ;
 wire \id_stage_i.controller_i.instr_valid_i ;
 wire \id_stage_i.controller_i.load_err_q ;
 wire \id_stage_i.controller_i.nmi_mode_d ;
 wire \id_stage_i.controller_i.store_err_q ;
 wire \id_stage_i.decoder_i.illegal_c_insn_i ;
 wire \id_stage_i.id_fsm_q ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_q ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net538;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire \load_store_unit_i.data_sign_ext_q ;
 wire \load_store_unit_i.data_we_q ;
 wire \load_store_unit_i.handle_misaligned_q ;
 wire \load_store_unit_i.lsu_err_q ;
 wire net437;
 wire net438;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net5782;
 wire net8153;
 wire net5781;
 wire net5780;
 wire net5832;
 wire net5779;
 wire net5778;
 wire net5783;
 wire net5802;
 wire net5809;
 wire net5827;
 wire net5788;
 wire net5787;
 wire net5789;
 wire net5786;
 wire net5785;
 wire net5796;
 wire net5795;
 wire net5794;
 wire net5793;
 wire net5792;
 wire net5797;
 wire net5803;
 wire net5801;
 wire net5800;
 wire net5799;
 wire net5798;
 wire net5807;
 wire net5806;
 wire net5805;
 wire net5804;
 wire net5808;
 wire net5815;
 wire net5814;
 wire net5813;
 wire net5812;
 wire net5811;
 wire net5810;
 wire net5822;
 wire net5831;
 wire net5823;
 wire net5821;
 wire net5820;
 wire net5834;
 wire net8151;
 wire net8150;
 wire net5833;
 wire net5837;
 wire net5836;
 wire net5835;
 wire net8149;
 wire net5858;
 wire net5842;
 wire net5863;
 wire net5841;
 wire net5840;
 wire net5839;
 wire net5838;
 wire net5857;
 wire net5843;
 wire net5856;
 wire net5855;
 wire net5849;
 wire net5851;
 wire net5848;
 wire net5850;
 wire net5844;
 wire net5846;
 wire net5845;
 wire net5854;
 wire net5847;
 wire net5852;
 wire net5862;
 wire net5861;
 wire net5853;
 wire net5860;
 wire net8135;
 wire net8134;
 wire net5880;
 wire net5867;
 wire net5878;
 wire net5877;
 wire net5876;
 wire net5875;
 wire net5872;
 wire net5873;
 wire net5868;
 wire net5871;
 wire net5870;
 wire net5885;
 wire net5883;
 wire net5881;
 wire net5882;
 wire net5911;
 wire net5890;
 wire net5889;
 wire net5899;
 wire net5888;
 wire net5887;
 wire net5891;
 wire net5898;
 wire net5897;
 wire net5896;
 wire net5895;
 wire net5904;
 wire net5903;
 wire net5902;
 wire net5901;
 wire net5900;
 wire net5953;
 wire net5910;
 wire net5909;
 wire net5952;
 wire net5908;
 wire net5905;
 wire net5916;
 wire net5906;
 wire net5915;
 wire net5914;
 wire net5913;
 wire net5907;
 wire net5912;
 wire net5920;
 wire net5919;
 wire net5921;
 wire net5918;
 wire net5917;
 wire net5950;
 wire net5949;
 wire net5948;
 wire net5947;
 wire net5946;
 wire net5945;
 wire net5942;
 wire net5944;
 wire net5943;
 wire net5941;
 wire net5926;
 wire net5927;
 wire net5961;
 wire net5933;
 wire net5930;
 wire net5931;
 wire net5979;
 wire net5957;
 wire net5954;
 wire net5966;
 wire net5990;
 wire net5965;
 wire net5964;
 wire net5963;
 wire net5962;
 wire net5980;
 wire net5971;
 wire net5972;
 wire net8103;
 wire net5989;
 wire net5988;
 wire net5983;
 wire net5987;
 wire net5986;
 wire net5985;
 wire net5991;
 wire net5981;
 wire net5977;
 wire net5978;
 wire net5976;
 wire net5975;
 wire net5968;
 wire net5970;
 wire net5967;
 wire net5973;
 wire net5969;
 wire net5974;
 wire net5984;
 wire net5982;
 wire net7919;
 wire net7918;
 wire net6042;
 wire net6007;
 wire net6006;
 wire net6005;
 wire net6004;
 wire net6003;
 wire net6002;
 wire net7915;
 wire net5992;
 wire net5993;
 wire net6040;
 wire net6011;
 wire net6050;
 wire net6010;
 wire net6039;
 wire net6009;
 wire net6041;
 wire net7917;
 wire net5994;
 wire net5995;
 wire net5996;
 wire net5997;
 wire net5998;
 wire net5999;
 wire net6000;
 wire net6001;
 wire net6008;
 wire net6015;
 wire net6033;
 wire net6014;
 wire net6013;
 wire net6012;
 wire net6027;
 wire net6022;
 wire net6021;
 wire net6020;
 wire net6018;
 wire net6016;
 wire net6028;
 wire net6019;
 wire net6017;
 wire net6026;
 wire net6025;
 wire net6024;
 wire net6023;
 wire net6038;
 wire net6032;
 wire net6031;
 wire net6030;
 wire net6029;
 wire net6037;
 wire net6036;
 wire net6035;
 wire net6034;
 wire net6046;
 wire net6045;
 wire net6044;
 wire net6043;
 wire net7912;
 wire net7911;
 wire net6067;
 wire net6055;
 wire net7914;
 wire net7913;
 wire net6054;
 wire net6053;
 wire net6052;
 wire net6051;
 wire net6079;
 wire net6065;
 wire net6064;
 wire net6063;
 wire net6077;
 wire net6062;
 wire net6056;
 wire net6078;
 wire net6066;
 wire net6075;
 wire net7910;
 wire net6076;
 wire net6059;
 wire net6057;
 wire net6061;
 wire net6058;
 wire net6060;
 wire net6068;
 wire net6069;
 wire net6091;
 wire net6074;
 wire net6090;
 wire net6089;
 wire net6084;
 wire net6088;
 wire net7909;
 wire net6085;
 wire net6087;
 wire net6070;
 wire net6071;
 wire net6072;
 wire net6073;
 wire net6083;
 wire net6166;
 wire net6108;
 wire net6107;
 wire net7906;
 wire net7905;
 wire net7908;
 wire net6094;
 wire net6093;
 wire net7904;
 wire net6095;
 wire net6106;
 wire net6105;
 wire net6104;
 wire net6165;
 wire net6113;
 wire net6112;
 wire net6111;
 wire net6110;
 wire net6114;
 wire net6096;
 wire net6097;
 wire net6098;
 wire net6099;
 wire net6100;
 wire net6101;
 wire net6102;
 wire net6103;
 wire net6120;
 wire net6119;
 wire net6118;
 wire net6109;
 wire net6115;
 wire net6163;
 wire net6117;
 wire net6116;
 wire net6162;
 wire net6161;
 wire net6153;
 wire net6155;
 wire net6130;
 wire net6132;
 wire net6171;
 wire net7900;
 wire net6176;
 wire net6175;
 wire net6136;
 wire net6169;
 wire net6133;
 wire net6135;
 wire net6174;
 wire net6137;
 wire net6138;
 wire net6139;
 wire net6141;
 wire net6142;
 wire net6143;
 wire net6144;
 wire net6145;
 wire net6147;
 wire net6149;
 wire net6150;
 wire net6152;
 wire net6154;
 wire net6156;
 wire net6158;
 wire net6159;
 wire net6160;
 wire net6173;
 wire net7899;
 wire net6182;
 wire net7898;
 wire net6181;
 wire net6180;
 wire net6185;
 wire net6179;
 wire net6178;
 wire net6177;
 wire net7897;
 wire net6186;
 wire net6192;
 wire net6188;
 wire net7896;
 wire net6191;
 wire net6187;
 wire net7895;
 wire net6190;
 wire net6198;
 wire net6197;
 wire net7894;
 wire net6199;
 wire net7804;
 wire net6196;
 wire net6200;
 wire net6195;
 wire net6194;
 wire net7803;
 wire net7802;
 wire net6203;
 wire net6208;
 wire net6202;
 wire net6207;
 wire net6206;
 wire net6205;
 wire net6201;
 wire net6213;
 wire net6212;
 wire net6215;
 wire net6211;
 wire net7801;
 wire net6210;
 wire net6209;
 wire net7800;
 wire net6214;
 wire net6220;
 wire net6219;
 wire net7799;
 wire net6218;
 wire net6224;
 wire net6223;
 wire net6222;
 wire net6221;
 wire net6217;
 wire net6227;
 wire net6226;
 wire net6267;
 wire net6229;
 wire net6228;
 wire net6225;
 wire net6232;
 wire net6231;
 wire net6230;
 wire net6238;
 wire net6237;
 wire net7798;
 wire net6234;
 wire net6240;
 wire net6236;
 wire net6235;
 wire net6239;
 wire net6233;
 wire net6247;
 wire net6246;
 wire net6249;
 wire net6245;
 wire net6244;
 wire net6248;
 wire net6243;
 wire net6242;
 wire net6241;
 wire net6251;
 wire net6258;
 wire net6250;
 wire net6257;
 wire net6256;
 wire net6254;
 wire net6255;
 wire net6253;
 wire net6252;
 wire net6263;
 wire net6262;
 wire net6261;
 wire net6266;
 wire net6265;
 wire net7797;
 wire net6259;
 wire net7796;
 wire net6264;
 wire net6260;
 wire net6270;
 wire net6269;
 wire net6273;
 wire net6294;
 wire net6268;
 wire net6276;
 wire net6275;
 wire net6272;
 wire net6278;
 wire net6277;
 wire net6282;
 wire net6285;
 wire net6281;
 wire net6279;
 wire net6284;
 wire net6280;
 wire net6290;
 wire net6293;
 wire net6287;
 wire net6292;
 wire net6288;
 wire net6289;
 wire net6291;
 wire net6286;
 wire net6355;
 wire net6303;
 wire net6300;
 wire net6299;
 wire net6298;
 wire net6302;
 wire net6296;
 wire net6295;
 wire net6297;
 wire net6301;
 wire net7794;
 wire net6308;
 wire net6307;
 wire net6306;
 wire net7793;
 wire net6305;
 wire net6304;
 wire net6310;
 wire net6309;
 wire net6314;
 wire net7792;
 wire net6318;
 wire net6317;
 wire net6313;
 wire net6312;
 wire net6311;
 wire net6316;
 wire net6315;
 wire net6322;
 wire net6321;
 wire net6320;
 wire net7791;
 wire net6319;
 wire net6326;
 wire net6325;
 wire net6324;
 wire net6323;
 wire net6345;
 wire net6333;
 wire net6332;
 wire net6329;
 wire net6331;
 wire net6328;
 wire net6330;
 wire net6334;
 wire net6327;
 wire net6335;
 wire net6343;
 wire net6342;
 wire net6341;
 wire net6340;
 wire net6339;
 wire net6338;
 wire net6336;
 wire net6344;
 wire net6337;
 wire net6348;
 wire net6347;
 wire net6352;
 wire net6346;
 wire net6351;
 wire net6354;
 wire net6350;
 wire net6349;
 wire net6358;
 wire net6357;
 wire net6356;
 wire net6362;
 wire net6361;
 wire net6360;
 wire net6393;
 wire net6359;
 wire net6363;
 wire net6392;
 wire net6365;
 wire net6376;
 wire net6368;
 wire net6367;
 wire net6366;
 wire net6364;
 wire net6375;
 wire net6374;
 wire net6369;
 wire net6372;
 wire net7783;
 wire net6370;
 wire net7782;
 wire net6371;
 wire net7790;
 wire net6394;
 wire net7789;
 wire net6380;
 wire net6379;
 wire net6390;
 wire net6378;
 wire net6377;
 wire net6382;
 wire net6381;
 wire net6391;
 wire net6384;
 wire net6383;
 wire net6389;
 wire net6388;
 wire net6387;
 wire net6386;
 wire net6385;
 wire net7787;
 wire net7786;
 wire net7785;
 wire net7784;
 wire net7788;
 wire net7781;
 wire net7779;
 wire net7780;
 wire net6395;
 wire net6413;
 wire net6414;
 wire net6429;
 wire net6430;
 wire net6428;
 wire net6397;
 wire net6418;
 wire net6447;
 wire net6421;
 wire net6419;
 wire net6440;
 wire net6420;
 wire net7778;
 wire net6432;
 wire net6431;
 wire net6439;
 wire net6453;
 wire net6438;
 wire net6434;
 wire net6433;
 wire net6437;
 wire net6435;
 wire net6436;
 wire net6446;
 wire net6474;
 wire net6462;
 wire net7777;
 wire net7776;
 wire net6472;
 wire net6473;
 wire net6443;
 wire net6442;
 wire net6444;
 wire net6445;
 wire net6441;
 wire net7775;
 wire net7747;
 wire net6461;
 wire net7745;
 wire net7746;
 wire net6457;
 wire net6454;
 wire net6455;
 wire net6478;
 wire net6465;
 wire net6511;
 wire net7585;
 wire net7744;
 wire net7743;
 wire net6501;
 wire net6500;
 wire net6479;
 wire net6456;
 wire net6458;
 wire net6464;
 wire net6459;
 wire net6460;
 wire net6463;
 wire net6468;
 wire net6471;
 wire net7742;
 wire net7741;
 wire net6467;
 wire net6466;
 wire net7740;
 wire net6469;
 wire net6470;
 wire net7739;
 wire net7738;
 wire net7717;
 wire net7716;
 wire net7715;
 wire net7712;
 wire net7714;
 wire net7713;
 wire net6494;
 wire net6496;
 wire net6510;
 wire net6503;
 wire net6504;
 wire net6502;
 wire net6509;
 wire net6512;
 wire net7584;
 wire net6531;
 wire net6530;
 wire net6529;
 wire net6516;
 wire net6515;
 wire net6517;
 wire net6514;
 wire net6513;
 wire net6521;
 wire net7583;
 wire net6536;
 wire net6528;
 wire net6520;
 wire net6519;
 wire net6522;
 wire net6535;
 wire net6518;
 wire net6524;
 wire net6523;
 wire net6527;
 wire net6532;
 wire net6526;
 wire net6525;
 wire net6541;
 wire net7582;
 wire net6540;
 wire net7581;
 wire net7580;
 wire net7579;
 wire net6537;
 wire net6533;
 wire net7578;
 wire net6539;
 wire net7549;
 wire net7280;
 wire net6557;
 wire net6568;
 wire net6534;
 wire net6538;
 wire net6546;
 wire net6552;
 wire net6542;
 wire net6545;
 wire net6543;
 wire net6550;
 wire net7290;
 wire net6551;
 wire net7324;
 wire net6544;
 wire net6547;
 wire net7376;
 wire net6549;
 wire net6548;
 wire net7375;
 wire net7374;
 wire net7373;
 wire net6553;
 wire net7360;
 wire net6554;
 wire net7372;
 wire net7371;
 wire net7362;
 wire net7361;
 wire net6590;
 wire net6571;
 wire net6573;
 wire net6575;
 wire net6583;
 wire net6578;
 wire net6582;
 wire net6589;
 wire net6585;
 wire net6588;
 wire net6592;
 wire net6600;
 wire net7238;
 wire net7239;
 wire net6604;
 wire net6605;
 wire net7095;
 wire net7089;
 wire net6669;
 wire net6610;
 wire net6667;
 wire net6617;
 wire net6625;
 wire net6666;
 wire net6665;
 wire net6632;
 wire net6631;
 wire net6629;
 wire net6635;
 wire net6636;
 wire net6637;
 wire net6644;
 wire net6638;
 wire net6639;
 wire net6643;
 wire net6642;
 wire net6657;
 wire net7038;
 wire net6652;
 wire net6650;
 wire net6651;
 wire net6649;
 wire net6656;
 wire net6725;
 wire net6662;
 wire net6655;
 wire net6654;
 wire net6724;
 wire net6653;
 wire net6658;
 wire net6661;
 wire net6659;
 wire net6660;
 wire net6677;
 wire net6727;
 wire net7058;
 wire net6672;
 wire net6671;
 wire net6670;
 wire net6723;
 wire net6821;
 wire net6793;
 wire net6676;
 wire net6673;
 wire net6675;
 wire net6722;
 wire net6721;
 wire net6681;
 wire net7037;
 wire net6720;
 wire net6731;
 wire net6730;
 wire net6792;
 wire net6791;
 wire net6823;
 wire net6680;
 wire net6674;
 wire net6678;
 wire net6679;
 wire net6694;
 wire net6685;
 wire net6684;
 wire net6683;
 wire net6682;
 wire net6686;
 wire net6689;
 wire net6688;
 wire net6687;
 wire net6693;
 wire net6692;
 wire net6691;
 wire net6690;
 wire net6719;
 wire net6698;
 wire net6697;
 wire net6696;
 wire net6695;
 wire net6702;
 wire net6701;
 wire net6700;
 wire net6699;
 wire net6718;
 wire net6711;
 wire net6704;
 wire net6703;
 wire net6706;
 wire net6705;
 wire net6768;
 wire net6767;
 wire net6728;
 wire net6710;
 wire net6707;
 wire net6717;
 wire net6708;
 wire net6709;
 wire net6713;
 wire net6712;
 wire net6747;
 wire net6714;
 wire net6716;
 wire net6822;
 wire net6715;
 wire net6735;
 wire net6729;
 wire net6733;
 wire net7460;
 wire net6734;
 wire net6748;
 wire net6752;
 wire net6766;
 wire net7382;
 wire net7370;
 wire net7357;
 wire net7363;
 wire net7369;
 wire net7384;
 wire net6732;
 wire net6739;
 wire net6738;
 wire net6737;
 wire net6736;
 wire net6744;
 wire net6743;
 wire net6750;
 wire net6746;
 wire net6745;
 wire net6751;
 wire net6764;
 wire net6741;
 wire net6742;
 wire net6740;
 wire net6765;
 wire net6749;
 wire net6753;
 wire net7353;
 wire net6763;
 wire net6869;
 wire net6755;
 wire net6820;
 wire net6870;
 wire net6754;
 wire net6756;
 wire net6758;
 wire net6757;
 wire net6776;
 wire net6761;
 wire net6759;
 wire net6762;
 wire net6775;
 wire net6769;
 wire net6760;
 wire net6773;
 wire net6771;
 wire net6774;
 wire net6770;
 wire net6772;
 wire net6797;
 wire net6780;
 wire net6779;
 wire net6789;
 wire net6778;
 wire net6788;
 wire net6781;
 wire net6777;
 wire net6790;
 wire net6803;
 wire net6784;
 wire net6786;
 wire net6794;
 wire net6819;
 wire net6785;
 wire net6787;
 wire net6802;
 wire net6796;
 wire net6783;
 wire net6812;
 wire net6782;
 wire net6818;
 wire net6811;
 wire net6795;
 wire net6857;
 wire net6826;
 wire net6800;
 wire net6801;
 wire net6846;
 wire net7036;
 wire net6851;
 wire net6842;
 wire net6843;
 wire net6798;
 wire net6799;
 wire net6810;
 wire net6805;
 wire net6804;
 wire net6806;
 wire net6809;
 wire net6807;
 wire net6808;
 wire net6824;
 wire net6813;
 wire net6969;
 wire net6817;
 wire net6816;
 wire net6814;
 wire net6815;
 wire net6871;
 wire net6841;
 wire net6840;
 wire net6839;
 wire net6838;
 wire net6837;
 wire net6827;
 wire net6825;
 wire net6829;
 wire net6835;
 wire net6868;
 wire net6834;
 wire net6867;
 wire net6831;
 wire net6833;
 wire net6830;
 wire net6832;
 wire net6847;
 wire net6836;
 wire net6828;
 wire net6968;
 wire net6844;
 wire net6845;
 wire net6877;
 wire net6850;
 wire net6874;
 wire net6872;
 wire net6873;
 wire net6876;
 wire net7350;
 wire net7352;
 wire net6849;
 wire net6848;
 wire net6854;
 wire net6856;
 wire net6852;
 wire net6855;
 wire net6853;
 wire net6859;
 wire net6858;
 wire net6866;
 wire net6875;
 wire net6865;
 wire net6864;
 wire net6863;
 wire net6907;
 wire net6861;
 wire net6860;
 wire net6862;
 wire net6912;
 wire net6878;
 wire net6879;
 wire net6906;
 wire net7351;
 wire net7354;
 wire net6886;
 wire net6880;
 wire net7349;
 wire net7347;
 wire net7348;
 wire net7344;
 wire net7044;
 wire net6885;
 wire net6881;
 wire net6882;
 wire net7345;
 wire net7346;
 wire net6899;
 wire net6884;
 wire net6883;
 wire net6905;
 wire net6891;
 wire net6889;
 wire net6887;
 wire net6896;
 wire net6888;
 wire net6897;
 wire net6898;
 wire net6901;
 wire net6890;
 wire net6893;
 wire net6892;
 wire net6894;
 wire net6895;
 wire net6900;
 wire net6902;
 wire net6911;
 wire net6903;
 wire net6904;
 wire net6908;
 wire net6909;
 wire net6910;
 wire net6913;
 wire net6915;
 wire net7039;
 wire net6916;
 wire net6914;
 wire net6919;
 wire net6939;
 wire net6918;
 wire net6917;
 wire net6929;
 wire net7032;
 wire net6928;
 wire net6922;
 wire net6921;
 wire net6920;
 wire net6945;
 wire net6967;
 wire net6925;
 wire net6923;
 wire net6924;
 wire net6941;
 wire net6927;
 wire net6938;
 wire net6926;
 wire net6940;
 wire net6932;
 wire net6931;
 wire net6930;
 wire net6942;
 wire net6937;
 wire net6933;
 wire net6936;
 wire net6944;
 wire net6935;
 wire net6943;
 wire net6934;
 wire net6947;
 wire net6946;
 wire net6960;
 wire net6958;
 wire net6957;
 wire net6959;
 wire net6956;
 wire net6951;
 wire net6948;
 wire net6966;
 wire net6949;
 wire net6953;
 wire net6965;
 wire net6950;
 wire net6952;
 wire net6954;
 wire net6955;
 wire net6964;
 wire net6963;
 wire net6961;
 wire net6962;
 wire net6976;
 wire net7030;
 wire net6970;
 wire net6977;
 wire net6971;
 wire net6972;
 wire net7027;
 wire net7031;
 wire net6973;
 wire net6974;
 wire net7043;
 wire net6975;
 wire net7023;
 wire net7035;
 wire net7024;
 wire net7029;
 wire net7028;
 wire net7033;
 wire net6980;
 wire net6979;
 wire net6978;
 wire net6981;
 wire net7025;
 wire net7022;
 wire net6982;
 wire net6988;
 wire net6983;
 wire net6984;
 wire net7026;
 wire net7016;
 wire net7004;
 wire net6985;
 wire net6987;
 wire net6986;
 wire net7021;
 wire net6996;
 wire net6989;
 wire net7020;
 wire net7019;
 wire net6995;
 wire net6992;
 wire net6990;
 wire net6991;
 wire net6999;
 wire net6994;
 wire net6993;
 wire net6997;
 wire net7003;
 wire net6998;
 wire net7018;
 wire net7001;
 wire net7000;
 wire net7002;
 wire net7015;
 wire net7013;
 wire net7010;
 wire net7005;
 wire net7012;
 wire net7006;
 wire net7011;
 wire net7008;
 wire net7009;
 wire net7014;
 wire net7007;
 wire net7017;
 wire net7034;
 wire net7041;
 wire net7042;
 wire net7049;
 wire net7048;
 wire net7057;
 wire net7040;
 wire net7046;
 wire net7056;
 wire net7055;
 wire net7060;
 wire net7047;
 wire net7054;
 wire net7059;
 wire net7289;
 wire net7088;
 wire net7342;
 wire net7050;
 wire net7051;
 wire net7063;
 wire net7087;
 wire net7053;
 wire net7064;
 wire net7052;
 wire net7077;
 wire net7086;
 wire net7062;
 wire net7061;
 wire net7078;
 wire net7079;
 wire net7085;
 wire net7094;
 wire net7065;
 wire net7070;
 wire net7067;
 wire net7073;
 wire net7068;
 wire net7069;
 wire net7066;
 wire net7071;
 wire net7072;
 wire net7082;
 wire net7074;
 wire net7075;
 wire net7076;
 wire net7080;
 wire net7081;
 wire net7083;
 wire net7090;
 wire net7084;
 wire net7091;
 wire net7093;
 wire net7092;
 wire net7101;
 wire net7171;
 wire net7097;
 wire net7165;
 wire net7166;
 wire net7096;
 wire net7099;
 wire net7098;
 wire net7287;
 wire net7100;
 wire net7281;
 wire net7276;
 wire net7285;
 wire net7288;
 wire net7117;
 wire net7108;
 wire net7102;
 wire net7129;
 wire net7103;
 wire net7275;
 wire net7116;
 wire net7107;
 wire net7274;
 wire net7105;
 wire net7104;
 wire net7106;
 wire net7115;
 wire net7109;
 wire net7110;
 wire net7124;
 wire net7123;
 wire net7119;
 wire net7111;
 wire net7112;
 wire net7113;
 wire net7114;
 wire net7118;
 wire net7122;
 wire net7267;
 wire net7128;
 wire net7120;
 wire net7197;
 wire net7269;
 wire net7127;
 wire net7121;
 wire net7126;
 wire net7125;
 wire net7154;
 wire net7132;
 wire net7131;
 wire net7130;
 wire net7155;
 wire net7233;
 wire net7135;
 wire net7133;
 wire net7139;
 wire net7175;
 wire net7174;
 wire net7138;
 wire net7134;
 wire net7151;
 wire net7143;
 wire net7137;
 wire net7136;
 wire net7142;
 wire net7140;
 wire net7141;
 wire net7145;
 wire net7144;
 wire net7147;
 wire net7146;
 wire net7150;
 wire net7149;
 wire net7148;
 wire net7153;
 wire net7152;
 wire net7161;
 wire net7156;
 wire net7158;
 wire net7157;
 wire net7160;
 wire net7159;
 wire net7170;
 wire net7173;
 wire net7164;
 wire net7162;
 wire net7163;
 wire net7169;
 wire net7168;
 wire net7167;
 wire net7208;
 wire net7180;
 wire net7176;
 wire net7228;
 wire net7178;
 wire net7187;
 wire net7177;
 wire net7179;
 wire net7186;
 wire net7181;
 wire net7183;
 wire net7182;
 wire net7194;
 wire net7185;
 wire net7184;
 wire net7265;
 wire net7188;
 wire net7190;
 wire net7189;
 wire net7193;
 wire net7192;
 wire net7191;
 wire net7264;
 wire net7195;
 wire net7254;
 wire net7196;
 wire net7200;
 wire net7198;
 wire net7199;
 wire net7207;
 wire net7203;
 wire net7202;
 wire net7201;
 wire net7216;
 wire net7206;
 wire net7205;
 wire net7204;
 wire net7215;
 wire net7210;
 wire net7209;
 wire net7212;
 wire net7278;
 wire net7224;
 wire net7211;
 wire net7279;
 wire net7214;
 wire net7213;
 wire net7220;
 wire net7219;
 wire net7217;
 wire net7218;
 wire net7222;
 wire net7221;
 wire net7223;
 wire net7227;
 wire net7226;
 wire net7225;
 wire net7246;
 wire net7231;
 wire net7229;
 wire net7230;
 wire net7232;
 wire net7237;
 wire net7236;
 wire net7234;
 wire net7235;
 wire net7245;
 wire net7244;
 wire net7241;
 wire net7243;
 wire net7249;
 wire net7247;
 wire net7242;
 wire net7248;
 wire net7250;
 wire net7258;
 wire net7251;
 wire net7252;
 wire net7253;
 wire net7263;
 wire net7256;
 wire net7257;
 wire net7255;
 wire net7271;
 wire net7268;
 wire net7277;
 wire net7259;
 wire net7273;
 wire net7260;
 wire net7261;
 wire net7266;
 wire net7262;
 wire net7272;
 wire net7270;
 wire net7282;
 wire net7283;
 wire net7294;
 wire net7286;
 wire net7284;
 wire net7296;
 wire net7295;
 wire net7291;
 wire net7292;
 wire net7341;
 wire net7298;
 wire net7300;
 wire net7340;
 wire net7293;
 wire net7297;
 wire net7299;
 wire net7301;
 wire net7312;
 wire net7305;
 wire net7304;
 wire net7339;
 wire net7311;
 wire net7310;
 wire net7302;
 wire net7358;
 wire net7337;
 wire net7359;
 wire net7303;
 wire net7306;
 wire net7316;
 wire net7307;
 wire net7317;
 wire net7308;
 wire net7309;
 wire net7315;
 wire net7313;
 wire net7323;
 wire net7314;
 wire net7322;
 wire net7321;
 wire net7318;
 wire net7320;
 wire net7319;
 wire net7327;
 wire net7325;
 wire net7343;
 wire net7334;
 wire net7326;
 wire net7338;
 wire net7332;
 wire net7335;
 wire net7331;
 wire net7333;
 wire net7336;
 wire net7328;
 wire net7329;
 wire net7330;
 wire net7356;
 wire net7355;
 wire net7365;
 wire net7367;
 wire net7366;
 wire net7368;
 wire net7510;
 wire net7377;
 wire net7364;
 wire net7429;
 wire net7383;
 wire net7379;
 wire net7380;
 wire net7381;
 wire net7509;
 wire net7378;
 wire clknet_1_1_0__06563_;
 wire net7385;
 wire clknet_3_6_0__06563_;
 wire net7428;
 wire net7398;
 wire net7387;
 wire clknet_leaf_49__06563_;
 wire net7427;
 wire net7413;
 wire net7408;
 wire delaynet_2_core_clock;
 wire clknet_1_0_0__06563_;
 wire clknet_0__06563_;
 wire clknet_leaf_51__06563_;
 wire clknet_leaf_50__06563_;
 wire net7386;
 wire net7389;
 wire delaynet_1_core_clock;
 wire clknet_leaf_44__06563_;
 wire clknet_leaf_48__06563_;
 wire clknet_leaf_47__06563_;
 wire clknet_leaf_46__06563_;
 wire delaynet_0_core_clock;
 wire net7388;
 wire net7391;
 wire net7390;
 wire net7394;
 wire net7393;
 wire net7392;
 wire clknet_leaf_28__06563_;
 wire net7395;
 wire net7396;
 wire net7397;
 wire clknet_leaf_43__06563_;
 wire net7399;
 wire net7403;
 wire net7402;
 wire net7400;
 wire net7401;
 wire clknet_leaf_32__06563_;
 wire clknet_leaf_36__06563_;
 wire clknet_leaf_35__06563_;
 wire clknet_leaf_34__06563_;
 wire net7405;
 wire net7404;
 wire net8102;
 wire net7407;
 wire net7406;
 wire net8030;
 wire net7412;
 wire net7409;
 wire net7417;
 wire net7411;
 wire net7410;
 wire net7416;
 wire net7415;
 wire net7414;
 wire net7418;
 wire net7419;
 wire net7423;
 wire net7420;
 wire net7923;
 wire net7455;
 wire net7434;
 wire net7422;
 wire net7421;
 wire net7454;
 wire net7922;
 wire net7426;
 wire net7424;
 wire net7425;
 wire net7430;
 wire net7453;
 wire net7445;
 wire net7947;
 wire net7945;
 wire net7925;
 wire net7431;
 wire net8002;
 wire net7921;
 wire net7920;
 wire net7432;
 wire net7433;
 wire net7436;
 wire net7435;
 wire net7437;
 wire net7441;
 wire net7444;
 wire net7438;
 wire net7439;
 wire net7440;
 wire net7442;
 wire net7449;
 wire net7443;
 wire net7446;
 wire net7452;
 wire net7447;
 wire net7459;
 wire net7448;
 wire net7450;
 wire net7458;
 wire net7451;
 wire net7457;
 wire net7456;
 wire net7470;
 wire net7469;
 wire net7462;
 wire net7464;
 wire net7463;
 wire net7924;
 wire net7465;
 wire net7468;
 wire net7467;
 wire net7946;
 wire net7508;
 wire net7466;
 wire net7472;
 wire net7492;
 wire net7473;
 wire net7471;
 wire net7480;
 wire net7474;
 wire net8101;
 wire net7491;
 wire net7481;
 wire net8001;
 wire net8073;
 wire net7475;
 wire net7476;
 wire net8052;
 wire net7479;
 wire net7477;
 wire net7490;
 wire net7478;
 wire net7482;
 wire net7486;
 wire net7484;
 wire net7485;
 wire net7483;
 wire net8051;
 wire net7489;
 wire net7496;
 wire net7498;
 wire net7488;
 wire net7487;
 wire net7495;
 wire net7497;
 wire net7494;
 wire net7493;
 wire net7503;
 wire net7507;
 wire net7499;
 wire net7506;
 wire net7505;
 wire net7500;
 wire net7502;
 wire net7501;
 wire net8031;
 wire net7512;
 wire net7711;
 wire net7511;
 wire net7524;
 wire net7710;
 wire net7515;
 wire net7504;
 wire net7514;
 wire net7513;
 wire net7518;
 wire net7517;
 wire net7523;
 wire net7519;
 wire net7516;
 wire net7591;
 wire net7547;
 wire net7522;
 wire net7521;
 wire net7520;
 wire net7540;
 wire net7566;
 wire net7526;
 wire net7534;
 wire net7539;
 wire net7525;
 wire net7527;
 wire net7533;
 wire net7541;
 wire net7538;
 wire net7546;
 wire net7529;
 wire net7528;
 wire net7532;
 wire net7530;
 wire net7531;
 wire net7536;
 wire net7537;
 wire net7535;
 wire net7542;
 wire net7545;
 wire net7544;
 wire net7543;
 wire net7565;
 wire net7553;
 wire net7556;
 wire net7555;
 wire net7554;
 wire net7552;
 wire net7551;
 wire net7550;
 wire net7560;
 wire net7559;
 wire net7557;
 wire net7588;
 wire net7592;
 wire net7558;
 wire net7587;
 wire net7708;
 wire net7705;
 wire net7709;
 wire net7707;
 wire net7586;
 wire net7561;
 wire net7564;
 wire net7577;
 wire net7563;
 wire net7562;
 wire net7569;
 wire net7571;
 wire net7568;
 wire net7567;
 wire net7570;
 wire net7576;
 wire net7575;
 wire net7574;
 wire net7572;
 wire net7573;
 wire net7648;
 wire net7706;
 wire net7647;
 wire net7625;
 wire net7646;
 wire net7645;
 wire net7590;
 wire net7589;
 wire net7596;
 wire net7606;
 wire net7805;
 wire net7893;
 wire net7829;
 wire net7891;
 wire net7828;
 wire net7812;
 wire net7811;
 wire net7827;
 wire net7813;
 wire net7826;
 wire net7806;
 wire net7816;
 wire net7892;
 wire net7595;
 wire net7594;
 wire net7593;
 wire net7604;
 wire net7601;
 wire net7605;
 wire net7597;
 wire net7624;
 wire net7598;
 wire net7815;
 wire net7890;
 wire net7814;
 wire net7599;
 wire net7607;
 wire net7600;
 wire net7603;
 wire net7602;
 wire net7623;
 wire net7615;
 wire net7608;
 wire net7609;
 wire net7834;
 wire net7832;
 wire net7831;
 wire net7610;
 wire net7611;
 wire net7612;
 wire net7830;
 wire net7613;
 wire net7833;
 wire net7614;
 wire net7889;
 wire net7616;
 wire net7617;
 wire net7858;
 wire net7618;
 wire net7619;
 wire net7620;
 wire net7857;
 wire net7621;
 wire net7704;
 wire net7622;
 wire net7644;
 wire net7639;
 wire net7626;
 wire net7634;
 wire net7627;
 wire net7652;
 wire net7654;
 wire net7653;
 wire net7628;
 wire net7631;
 wire net7629;
 wire net7633;
 wire net7630;
 wire net7632;
 wire net7635;
 wire net7636;
 wire net7650;
 wire net7637;
 wire net7638;
 wire net7643;
 wire net7642;
 wire net7640;
 wire net7651;
 wire net7641;
 wire net7656;
 wire net7649;
 wire net7655;
 wire net7690;
 wire net7671;
 wire net7659;
 wire net7670;
 wire net7703;
 wire net7657;
 wire net7663;
 wire net7664;
 wire net7835;
 wire net7691;
 wire net7856;
 wire net7718;
 wire net7658;
 wire net7737;
 wire net7720;
 wire net7719;
 wire net7722;
 wire net7750;
 wire net7749;
 wire net7748;
 wire net7774;
 wire net7660;
 wire net7661;
 wire net7669;
 wire net7665;
 wire net7662;
 wire net7668;
 wire net7689;
 wire net7666;
 wire net7672;
 wire net7688;
 wire net7667;
 wire net7687;
 wire net7674;
 wire net7673;
 wire net7726;
 wire net7724;
 wire net7725;
 wire net7736;
 wire net7721;
 wire net7675;
 wire net7686;
 wire net7676;
 wire net7735;
 wire net7723;
 wire net7677;
 wire net7697;
 wire net7696;
 wire net7678;
 wire net7679;
 wire net7680;
 wire net7694;
 wire net7681;
 wire net7695;
 wire net7682;
 wire net7683;
 wire net7684;
 wire net7685;
 wire net7693;
 wire net7692;
 wire net7734;
 wire net7730;
 wire net7700;
 wire net7702;
 wire net7699;
 wire net7698;
 wire net7701;
 wire net7731;
 wire net7729;
 wire net7733;
 wire net7732;
 wire net7728;
 wire net7727;
 wire net7760;
 wire net7762;
 wire net7759;
 wire net7758;
 wire net7757;
 wire net7772;
 wire net7756;
 wire net7753;
 wire net7761;
 wire net7771;
 wire net7751;
 wire net7768;
 wire net7764;
 wire net7763;
 wire net7767;
 wire net7752;
 wire net7765;
 wire net7770;
 wire net7766;
 wire net7769;
 wire net7755;
 wire net7754;
 wire net7773;
 wire net7861;
 wire net7868;
 wire net7873;
 wire net7872;
 wire net7867;
 wire net7863;
 wire net7866;
 wire net7855;
 wire net7865;
 wire net7864;
 wire net7869;
 wire net7888;
 wire net7887;
 wire net7871;
 wire net7862;
 wire net7870;
 wire net7859;
 wire net7874;
 wire net7885;
 wire net7875;
 wire net7886;
 wire net7884;
 wire net7883;
 wire net7876;
 wire net7882;
 wire net7881;
 wire net7877;
 wire net7878;
 wire net7879;
 wire net7880;
 wire net7860;
 wire net7854;
 wire net7808;
 wire net7849;
 wire net7853;
 wire net7848;
 wire net7807;
 wire net7836;
 wire net7823;
 wire net7825;
 wire net7822;
 wire net7837;
 wire net8075;
 wire net7850;
 wire net7852;
 wire net7851;
 wire net8080;
 wire net8050;
 wire net8079;
 wire net8078;
 wire net8077;
 wire net8033;
 wire net8083;
 wire net8064;
 wire net8072;
 wire net8100;
 wire net8053;
 wire net8071;
 wire net8067;
 wire net8066;
 wire net8065;
 wire net8063;
 wire net8062;
 wire net8070;
 wire net8069;
 wire net8068;
 wire net8061;
 wire net8060;
 wire net8057;
 wire net8059;
 wire net8056;
 wire net8055;
 wire net8054;
 wire net8058;
 wire net8049;
 wire net8048;
 wire net8047;
 wire net8039;
 wire net8038;
 wire net8043;
 wire net8045;
 wire net8040;
 wire net8034;
 wire net8037;
 wire net8044;
 wire net8042;
 wire net8041;
 wire net8046;
 wire net8036;
 wire net8035;
 wire net8032;
 wire net7810;
 wire net7809;
 wire net7818;
 wire net7819;
 wire net7824;
 wire net7820;
 wire net7821;
 wire net7817;
 wire net7845;
 wire net7841;
 wire net7847;
 wire net7844;
 wire net7839;
 wire net7843;
 wire net7838;
 wire net7846;
 wire net7842;
 wire net7840;
 wire net8088;
 wire net8084;
 wire net8087;
 wire net8076;
 wire net8086;
 wire net8082;
 wire net8098;
 wire net8097;
 wire net8096;
 wire net8095;
 wire net8085;
 wire net8094;
 wire net8081;
 wire net8093;
 wire net8090;
 wire net8089;
 wire net8092;
 wire net8091;
 wire net8099;
 wire net8074;
 wire net7944;
 wire clknet_2_3_0_clk_i_regs;
 wire clknet_leaf_1_clk_i_regs;
 wire net7926;
 wire net7942;
 wire clknet_1_0__leaf_clk_i;
 wire net7928;
 wire net7927;
 wire net7943;
 wire clknet_0_clk_i;
 wire clknet_leaf_22_clk_i_regs;
 wire clknet_leaf_11_clk_i_regs;
 wire clknet_leaf_8_clk_i_regs;
 wire clknet_leaf_5_clk_i_regs;
 wire clknet_leaf_2_clk_i_regs;
 wire clknet_leaf_10_clk_i_regs;
 wire clknet_leaf_4_clk_i_regs;
 wire clknet_leaf_3_clk_i_regs;
 wire clknet_leaf_6_clk_i_regs;
 wire clknet_leaf_26_clk_i_regs;
 wire clknet_leaf_7_clk_i_regs;
 wire clknet_leaf_9_clk_i_regs;
 wire clknet_leaf_16_clk_i_regs;
 wire clknet_leaf_24_clk_i_regs;
 wire clknet_leaf_15_clk_i_regs;
 wire clknet_leaf_14_clk_i_regs;
 wire clknet_leaf_12_clk_i_regs;
 wire clknet_leaf_13_clk_i_regs;
 wire clknet_leaf_31__06563_;
 wire clknet_leaf_20_clk_i_regs;
 wire clknet_leaf_19_clk_i_regs;
 wire clknet_leaf_17_clk_i_regs;
 wire clknet_leaf_21__06563_;
 wire clknet_leaf_18_clk_i_regs;
 wire clknet_leaf_20__06563_;
 wire clknet_2_2_0_clk_i_regs;
 wire clknet_leaf_25_clk_i_regs;
 wire clknet_leaf_23_clk_i_regs;
 wire clknet_leaf_21_clk_i_regs;
 wire clknet_leaf_19__06563_;
 wire clknet_3_3_0_clk_i_regs;
 wire clknet_3_2_0_clk_i_regs;
 wire clknet_leaf_1__06563_;
 wire clknet_3_1_0_clk_i_regs;
 wire clknet_leaf_27__06563_;
 wire clknet_3_0_0_clk_i_regs;
 wire clknet_leaf_0__06563_;
 wire clknet_3_7_0_clk_i_regs;
 wire clknet_3_6_0_clk_i_regs;
 wire clknet_3_5_0_clk_i_regs;
 wire clknet_leaf_24__06563_;
 wire clknet_leaf_23__06563_;
 wire clknet_leaf_30__06563_;
 wire clknet_leaf_18__06563_;
 wire clknet_leaf_2__06563_;
 wire clknet_leaf_6__06563_;
 wire clknet_leaf_17__06563_;
 wire clknet_leaf_4__06563_;
 wire clknet_leaf_5__06563_;
 wire clknet_leaf_3__06563_;
 wire clknet_leaf_15__06563_;
 wire clknet_leaf_33__06563_;
 wire clknet_leaf_14__06563_;
 wire clknet_leaf_7__06563_;
 wire clknet_leaf_22__06563_;
 wire clknet_leaf_12__06563_;
 wire clknet_leaf_9__06563_;
 wire clknet_leaf_16__06563_;
 wire clknet_leaf_8__06563_;
 wire clknet_leaf_13__06563_;
 wire clknet_leaf_10__06563_;
 wire clknet_leaf_11__06563_;
 wire clknet_leaf_42__06563_;
 wire clknet_leaf_26__06563_;
 wire clknet_3_4_0_clk_i_regs;
 wire clknet_leaf_25__06563_;
 wire clknet_leaf_41__06563_;
 wire clknet_leaf_45__06563_;
 wire clknet_leaf_38__06563_;
 wire clknet_leaf_37__06563_;
 wire clknet_leaf_40__06563_;
 wire clknet_leaf_39__06563_;
 wire clknet_leaf_29__06563_;
 wire net7930;
 wire net7929;
 wire net7976;
 wire net7951;
 wire net7931;
 wire net7950;
 wire net7955;
 wire clk_i_regs;
 wire net7935;
 wire net7934;
 wire net7932;
 wire net7936;
 wire net7933;
 wire net7940;
 wire net7941;
 wire net7949;
 wire net7948;
 wire net7937;
 wire net7939;
 wire net7953;
 wire net7966;
 wire net7938;
 wire net7952;
 wire net7954;
 wire net7956;
 wire net7965;
 wire net7959;
 wire net7964;
 wire net7957;
 wire net7958;
 wire net8286;
 wire net7960;
 wire net7961;
 wire clknet_leaf_0_clk_i_regs;
 wire net7962;
 wire net7963;
 wire net8287;
 wire net7975;
 wire net7968;
 wire net7967;
 wire net7974;
 wire net7971;
 wire net7969;
 wire net7973;
 wire clknet_2_1_0_clk_i_regs;
 wire net7970;
 wire net7972;
 wire clknet_leaf_27_clk_i_regs;
 wire net7999;
 wire net7998;
 wire net7990;
 wire net7989;
 wire net7983;
 wire net7977;
 wire clknet_2_0_0_clk_i_regs;
 wire net7997;
 wire net7991;
 wire net8000;
 wire net8029;
 wire net7978;
 wire net8003;
 wire net7986;
 wire net8028;
 wire net7996;
 wire clknet_1_0_0_clk_i_regs;
 wire clknet_leaf_34_clk_i_regs;
 wire clknet_leaf_44_clk_i_regs;
 wire clknet_1_1_0_clk_i_regs;
 wire clknet_leaf_28_clk_i_regs;
 wire net7979;
 wire net7980;
 wire net7981;
 wire net7982;
 wire net7984;
 wire net7985;
 wire net7992;
 wire net7995;
 wire net7988;
 wire net7987;
 wire net7994;
 wire net7993;
 wire net8005;
 wire net8008;
 wire net8004;
 wire net8007;
 wire net8027;
 wire net8006;
 wire net8026;
 wire net8015;
 wire clknet_leaf_33_clk_i_regs;
 wire net8013;
 wire net8010;
 wire net8009;
 wire clknet_leaf_31_clk_i_regs;
 wire clknet_leaf_40_clk_i_regs;
 wire net8014;
 wire clknet_leaf_43_clk_i_regs;
 wire clknet_leaf_30_clk_i_regs;
 wire clknet_leaf_32_clk_i_regs;
 wire clknet_leaf_29_clk_i_regs;
 wire net8011;
 wire net8025;
 wire net8012;
 wire net8022;
 wire clknet_leaf_39_clk_i_regs;
 wire clknet_leaf_35_clk_i_regs;
 wire net8016;
 wire net8020;
 wire net8017;
 wire clknet_leaf_42_clk_i_regs;
 wire clknet_leaf_36_clk_i_regs;
 wire clknet_leaf_38_clk_i_regs;
 wire clknet_leaf_37_clk_i_regs;
 wire net8018;
 wire clknet_leaf_41_clk_i_regs;
 wire net8019;
 wire clknet_0_clk_i_regs;
 wire net8021;
 wire clknet_leaf_45_clk_i_regs;
 wire net8024;
 wire net8023;
 wire clknet_leaf_47_clk_i_regs;
 wire clknet_leaf_46_clk_i_regs;
 wire clknet_leaf_48_clk_i_regs;
 wire net5761;
 wire net8142;
 wire net8162;
 wire net5765;
 wire net5762;
 wire net5764;
 wire net5763;
 wire net5766;
 wire net8155;
 wire net5767;
 wire net5768;
 wire net5819;
 wire net5769;
 wire net5771;
 wire net5770;
 wire net5818;
 wire net8161;
 wire net8160;
 wire net8157;
 wire net8156;
 wire net8158;
 wire net8159;
 wire net8163;
 wire net8171;
 wire net8164;
 wire net8165;
 wire net8170;
 wire net8166;
 wire net8168;
 wire net8167;
 wire net8169;
 wire net8187;
 wire net8186;
 wire net8185;
 wire net8183;
 wire net8175;
 wire net8173;
 wire net8172;
 wire net8174;
 wire net8182;
 wire net8180;
 wire net8176;
 wire net8178;
 wire net8177;
 wire net8179;
 wire net8181;
 wire net8184;
 wire net8248;
 wire net8189;
 wire net8188;
 wire net8200;
 wire net8190;
 wire net8199;
 wire net8192;
 wire net8191;
 wire net8193;
 wire net8198;
 wire net8195;
 wire net8194;
 wire net8196;
 wire net8197;
 wire net8247;
 wire net8203;
 wire net8202;
 wire net8201;
 wire net8220;
 wire net8204;
 wire net8205;
 wire net8219;
 wire net8206;
 wire net8210;
 wire net8209;
 wire net8208;
 wire net8207;
 wire net8218;
 wire net8211;
 wire net8212;
 wire net8217;
 wire net8215;
 wire net8214;
 wire net8213;
 wire net8216;
 wire net8246;
 wire net8224;
 wire net8222;
 wire net8221;
 wire net8223;
 wire net8225;
 wire net8245;
 wire net8226;
 wire net8228;
 wire net8227;
 wire net8243;
 wire net8242;
 wire net8234;
 wire net8229;
 wire net8233;
 wire net8231;
 wire net8230;
 wire net8232;
 wire net8241;
 wire net8235;
 wire net8239;
 wire net8236;
 wire net8238;
 wire net8237;
 wire net8240;
 wire net8244;
 wire net8249;
 wire net8255;
 wire net8250;
 wire net8251;
 wire net8254;
 wire net8252;
 wire net8253;
 wire net8279;
 wire net8259;
 wire net8257;
 wire net8256;
 wire net8258;
 wire net8260;
 wire net8278;
 wire net8262;
 wire net8261;
 wire net8264;
 wire net8263;
 wire net8277;
 wire net8266;
 wire net8265;
 wire net8276;
 wire net8274;
 wire net8273;
 wire net8268;
 wire net8267;
 wire net8272;
 wire net8269;
 wire net8270;
 wire net8271;
 wire net8275;
 wire net8280;
 wire net8283;
 wire net8281;
 wire net8282;
 wire net8284;
 wire net8285;
 wire net5773;
 wire net5772;
 wire net5817;
 wire net5816;
 wire net5774;
 wire net5791;
 wire net5784;
 wire net5777;
 wire net5776;
 wire net5775;
 wire net5790;
 wire net5826;
 wire net5825;
 wire net5824;
 wire net5830;
 wire net5829;
 wire net5828;
 wire net8154;
 wire net8140;
 wire net8139;
 wire net8141;
 wire net8138;
 wire net8148;
 wire net8147;
 wire net8143;
 wire net8146;
 wire net8144;
 wire net8145;
 wire net8152;
 wire net5859;
 wire net8137;
 wire net5866;
 wire net5865;
 wire net5864;
 wire net8136;
 wire net5874;
 wire net5879;
 wire net5869;
 wire net5884;
 wire net8133;
 wire net5893;
 wire net5892;
 wire net5886;
 wire net8132;
 wire net8124;
 wire net8123;
 wire net5894;
 wire net8131;
 wire net8126;
 wire net8125;
 wire net8130;
 wire net8128;
 wire net8127;
 wire net8129;
 wire net8122;
 wire net5951;
 wire net5940;
 wire net5922;
 wire net5939;
 wire net5923;
 wire net5929;
 wire net5928;
 wire net5938;
 wire net5924;
 wire net5925;
 wire net5934;
 wire net5932;
 wire net5936;
 wire net5935;
 wire net5937;
 wire net5960;
 wire net5955;
 wire net5959;
 wire net5958;
 wire net8119;
 wire net8117;
 wire net8116;
 wire net8115;
 wire net8105;
 wire net8104;
 wire net8114;
 wire net8107;
 wire net8106;
 wire net8113;
 wire net8110;
 wire net8109;
 wire net8108;
 wire net8112;
 wire net8111;
 wire net8118;
 wire net8120;
 wire net8121;
 wire net6049;
 wire net6048;
 wire net6047;
 wire net7916;
 wire net6082;
 wire net6080;
 wire net6081;
 wire net6086;
 wire net6092;
 wire net7901;
 wire net6168;
 wire net6167;
 wire net7903;
 wire net7902;
 wire net7907;
 wire net6157;
 wire net6121;
 wire net6164;
 wire net6128;
 wire net6129;
 wire net6127;
 wire net6125;
 wire net6126;
 wire net6131;
 wire net6134;
 wire net6151;
 wire net6140;
 wire net6146;
 wire net6148;
 wire net6170;
 wire net6172;
 wire net6183;
 wire net6184;
 wire net6189;
 wire net6193;
 wire net6204;
 wire net6216;
 wire net7795;
 wire net6271;
 wire net6274;
 wire net6283;
 wire net6353;
 wire net6373;
 wire net6399;
 wire net6398;
 wire net6400;
 wire net6412;
 wire net6411;
 wire net6410;
 wire net6409;
 wire net6408;
 wire net6407;
 wire net6406;
 wire net6405;
 wire net6422;
 wire net6417;
 wire net6416;
 wire net6415;
 wire net6427;
 wire net6426;
 wire net6423;
 wire net6424;
 wire net6425;
 wire net6452;
 wire net6450;
 wire net6449;
 wire net6448;
 wire net6451;
 wire net6499;
 wire net6498;
 wire net6497;
 wire net6492;
 wire net6491;
 wire net6490;
 wire net6489;
 wire net6487;
 wire net6488;
 wire net6493;
 wire net6495;
 wire net6507;
 wire net6506;
 wire net6505;
 wire net6508;
 wire net6567;
 wire net6569;
 wire net6591;
 wire net6570;
 wire net6572;
 wire net6574;
 wire net6576;
 wire net6577;
 wire net6580;
 wire net6579;
 wire net6581;
 wire net6584;
 wire net6586;
 wire net6587;
 wire net7240;
 wire net6599;
 wire net7172;
 wire net6602;
 wire net6601;
 wire net6603;
 wire net6606;
 wire net6607;
 wire net6608;
 wire net6609;
 wire net6668;
 wire net6611;
 wire net6613;
 wire net6612;
 wire net6615;
 wire net6614;
 wire net6621;
 wire net6620;
 wire net6623;
 wire net6622;
 wire net6624;
 wire net6626;
 wire net6627;
 wire net6628;
 wire net6630;
 wire net6663;
 wire net6664;
 wire net6640;
 wire net6641;
 wire net6645;
 wire net6646;
 wire net6648;
 wire net6647;
 wire net6726;
 wire net7045;
 wire net7461;
 wire net7548;
 wire clknet_3_4_0__06563_;
 wire clknet_3_3_0__06563_;
 wire clknet_2_1_0__06563_;
 wire clknet_2_0_0__06563_;
 wire clknet_3_2_0__06563_;
 wire clknet_3_0_0__06563_;
 wire clknet_2_2_0__06563_;
 wire clknet_2_3_0__06563_;
 wire clknet_3_1_0__06563_;
 wire clknet_3_5_0__06563_;
 wire clknet_3_7_0__06563_;

 sg13g2_tielo _15585__1 (.L_LO(alert_major_o));
 sg13g2_tielo _15586__2 (.L_LO(alert_minor_o));
 sg13g2_tielo _15587__3 (.L_LO(data_addr_o[0]));
 sg13g2_tielo _15588__4 (.L_LO(data_addr_o[1]));
 sg13g2_tielo _15589__5 (.L_LO(instr_addr_o[0]));
 sg13g2_tielo _15590__6 (.L_LO(instr_addr_o[1]));
 ALU_34_0_34_0_34_KOGGE_STONE _15591_ (.A({_06506_,
    _06463_,
    _06407_,
    _06322_,
    _06234_,
    _06141_,
    _06064_,
    _05955_,
    _05861_,
    _05741_,
    _05631_,
    _05527_,
    _05417_,
    _05275_,
    _05172_,
    _05051_,
    _04949_,
    _04831_,
    _04705_,
    _04604_,
    _04524_,
    _04443_,
    _04364_,
    _04288_,
    _04211_,
    _04141_,
    _04077_,
    _04003_,
    _03961_,
    _03930_,
    _03896_,
    _03865_,
    _03844_,
    _03832_}),
    .B({_06562_,
    _06559_,
    _06551_,
    _06549_,
    _06545_,
    _06541_,
    _06540_,
    _06539_,
    _06537_,
    _06534_,
    _06530_,
    _06528_,
    _06526_,
    _06525_,
    _06524_,
    _06523_,
    _06520_,
    _06519_,
    _06516_,
    _06515_,
    _06514_,
    _06513_,
    _06511_,
    _06510_,
    _06509_,
    _04076_,
    _04001_,
    _03960_,
    _06507_,
    _03895_,
    net_4,
    net_3,
    net_2,
    net_1}),
    .BI(net),
    .CI(net_5),
    .CO({_00070_,
    _00069_,
    _00068_,
    _00067_,
    _00065_,
    _00064_,
    _00063_,
    _00062_,
    _00061_,
    _00060_,
    _00059_,
    _00058_,
    _00057_,
    _00056_,
    _00054_,
    _00053_,
    _00052_,
    _00051_,
    _00050_,
    _00049_,
    _00048_,
    _00047_,
    _00046_,
    _00045_,
    _00077_,
    _00076_,
    _00075_,
    _00074_,
    _00073_,
    _00072_,
    _00071_,
    _00066_,
    _00055_,
    _00044_}),
    .X({_00036_,
    _00035_,
    _00034_,
    _00033_,
    _00031_,
    _00030_,
    _00029_,
    _00028_,
    _00027_,
    _00026_,
    _00025_,
    _00024_,
    _00023_,
    _00022_,
    _00020_,
    _00019_,
    _00018_,
    _00017_,
    _00016_,
    _00015_,
    _00014_,
    _00013_,
    _00012_,
    _00011_,
    _00043_,
    _00042_,
    _00041_,
    _00040_,
    _00039_,
    _00038_,
    _00037_,
    _00032_,
    _00021_,
    _00010_}),
    .Y({_00104_,
    _00103_,
    _00102_,
    _00101_,
    _00099_,
    _00098_,
    _00097_,
    _00096_,
    _00095_,
    _00094_,
    _00093_,
    _00092_,
    _00091_,
    _00090_,
    _00088_,
    _00087_,
    _00086_,
    _00085_,
    _00084_,
    _00083_,
    _00082_,
    _00081_,
    _00080_,
    _00079_,
    _00111_,
    _00110_,
    _00109_,
    _00108_,
    _00107_,
    _00106_,
    _00105_,
    _00100_,
    _00089_,
    _00078_}));
 sg13g2_tielo _15591__10 (.L_LO(net_3));
 sg13g2_tielo _15591__11 (.L_LO(net_4));
 sg13g2_tielo _15591__12 (.L_LO(net_5));
 sg13g2_tielo _15591__7 (.L_LO(net));
 sg13g2_tielo _15591__8 (.L_LO(net_1));
 sg13g2_tielo _15591__9 (.L_LO(net_2));
 sg13g2_o21ai_1 _15592_ (.B1(_15578_),
    .Y(_02012_),
    .A1(_15581_),
    .A2(_15582_));
 sg13g2_inv_1 _15593_ (.Y(_02013_),
    .A(_01680_));
 sg13g2_mux4_1 _15594_ (.S0(net7772),
    .A0(_01072_),
    .A1(_01107_),
    .A2(_01142_),
    .A3(_01177_),
    .S1(net7723),
    .X(_02014_));
 sg13g2_nand2b_1 _15595_ (.Y(_02015_),
    .B(net7433),
    .A_N(_02014_));
 sg13g2_inv_1 _15596_ (.Y(_02016_),
    .A(_01679_));
 sg13g2_mux4_1 _15597_ (.S0(net7772),
    .A0(_01212_),
    .A1(_01248_),
    .A2(_01283_),
    .A3(_01318_),
    .S1(net7723),
    .X(_02017_));
 sg13g2_or2_1 _15598_ (.X(_02018_),
    .B(_02017_),
    .A(net7587));
 sg13g2_mux2_1 _15599_ (.A0(_01494_),
    .A1(_01529_),
    .S(net7767),
    .X(_02019_));
 sg13g2_nor3_1 _15600_ (.A(net7579),
    .B(net7563),
    .C(_02019_),
    .Y(_02020_));
 sg13g2_mux2_1 _15601_ (.A0(_01424_),
    .A1(_01459_),
    .S(net7767),
    .X(_02021_));
 sg13g2_nor3_1 _15602_ (.A(net7582),
    .B(net7569),
    .C(_02021_),
    .Y(_02022_));
 sg13g2_mux2_1 _15603_ (.A0(_01353_),
    .A1(_01388_),
    .S(net7767),
    .X(_02023_));
 sg13g2_nor3_1 _15604_ (.A(net7579),
    .B(net7559),
    .C(_02023_),
    .Y(_02024_));
 sg13g2_inv_1 _15605_ (.Y(_02025_),
    .A(_01676_));
 sg13g2_mux2_1 _15606_ (.A0(_01564_),
    .A1(_00608_),
    .S(net7767),
    .X(_02026_));
 sg13g2_nor2_1 _15607_ (.A(net7553),
    .B(_02026_),
    .Y(_02027_));
 sg13g2_nor4_1 _15608_ (.A(_02020_),
    .B(_02022_),
    .C(_02024_),
    .D(_02027_),
    .Y(_02028_));
 sg13g2_inv_1 _15609_ (.Y(_02029_),
    .A(_01675_));
 sg13g2_nand4_1 _15610_ (.B(_02015_),
    .C(_02018_),
    .A(_02012_),
    .Y(_02030_),
    .D(_02028_));
 sg13g2_nor2_1 _15611_ (.A(net7291),
    .B(net7271),
    .Y(_02031_));
 sg13g2_a21oi_1 _15612_ (.A1(net7681),
    .A2(net7039),
    .Y(_02032_),
    .B1(_02031_));
 sg13g2_inv_1 _15613_ (.Y(_02033_),
    .A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_q ));
 sg13g2_nand2b_1 _15614_ (.Y(_02034_),
    .B(net8000),
    .A_N(_01641_));
 sg13g2_o21ai_1 _15615_ (.B1(_02034_),
    .Y(_02035_),
    .A1(_01671_),
    .A2(net7479));
 sg13g2_mux2_1 _15616_ (.A0(_01564_),
    .A1(_00608_),
    .S(net7865),
    .X(_02036_));
 sg13g2_nor2_1 _15617_ (.A(_10982_),
    .B(_02036_),
    .Y(_02037_));
 sg13g2_mux2_1 _15618_ (.A0(_01494_),
    .A1(_01529_),
    .S(net7865),
    .X(_02038_));
 sg13g2_nor3_1 _15619_ (.A(net7504),
    .B(net7490),
    .C(_02038_),
    .Y(_02039_));
 sg13g2_mux2_1 _15620_ (.A0(_00796_),
    .A1(_00828_),
    .S(_01892_),
    .X(_02040_));
 sg13g2_nor3_1 _15621_ (.A(_08892_),
    .B(_10182_),
    .C(_02040_),
    .Y(_02041_));
 sg13g2_mux2_1 _15622_ (.A0(_00860_),
    .A1(_00896_),
    .S(_01892_),
    .X(_02042_));
 sg13g2_nor3_1 _15623_ (.A(_08892_),
    .B(net7456),
    .C(_02042_),
    .Y(_02043_));
 sg13g2_nor4_1 _15624_ (.A(_02037_),
    .B(_02039_),
    .C(_02041_),
    .D(_02043_),
    .Y(_02044_));
 sg13g2_mux2_1 _15625_ (.A0(_01001_),
    .A1(_01036_),
    .S(net7865),
    .X(_02045_));
 sg13g2_nor3_1 _15626_ (.A(_08892_),
    .B(net7524),
    .C(_02045_),
    .Y(_02046_));
 sg13g2_mux2_1 _15627_ (.A0(_00931_),
    .A1(_00966_),
    .S(net7865),
    .X(_02047_));
 sg13g2_nor3_1 _15628_ (.A(_08892_),
    .B(net7504),
    .C(_02047_),
    .Y(_02048_));
 sg13g2_mux2_1 _15629_ (.A0(_01353_),
    .A1(_01388_),
    .S(net7865),
    .X(_02049_));
 sg13g2_nor3_1 _15630_ (.A(net7490),
    .B(_10182_),
    .C(_02049_),
    .Y(_02050_));
 sg13g2_mux2_1 _15631_ (.A0(_01424_),
    .A1(_01459_),
    .S(net7865),
    .X(_02051_));
 sg13g2_nor3_1 _15632_ (.A(net7490),
    .B(_10191_),
    .C(_02051_),
    .Y(_02052_));
 sg13g2_nor4_1 _15633_ (.A(_02046_),
    .B(_02048_),
    .C(_02050_),
    .D(_02052_),
    .Y(_02053_));
 sg13g2_mux2_1 _15634_ (.A0(_01302_),
    .A1(_00636_),
    .S(net7880),
    .X(_02054_));
 sg13g2_inv_1 _15635_ (.Y(_02055_),
    .A(_01667_));
 sg13g2_and2_1 _15636_ (.A(net7880),
    .B(_00950_),
    .X(_02056_));
 sg13g2_mux2_1 _15637_ (.A0(_00668_),
    .A1(_00700_),
    .S(net7880),
    .X(_02057_));
 sg13g2_mux2_1 _15638_ (.A0(_00732_),
    .A1(_00764_),
    .S(net7880),
    .X(_02058_));
 sg13g2_mux4_1 _15639_ (.S0(net7815),
    .A0(_02056_),
    .A1(_02057_),
    .A2(_02054_),
    .A3(_02058_),
    .S1(net7834),
    .X(_02059_));
 sg13g2_or2_1 _15640_ (.X(_02060_),
    .B(_02059_),
    .A(_08974_));
 sg13g2_mux4_1 _15641_ (.S0(net7918),
    .A0(_01072_),
    .A1(_01107_),
    .A2(_01142_),
    .A3(_01177_),
    .S1(net7831),
    .X(_02061_));
 sg13g2_nor3_1 _15642_ (.A(net7816),
    .B(_09073_),
    .C(_02061_),
    .Y(_02062_));
 sg13g2_mux4_1 _15643_ (.S0(net7918),
    .A0(_01212_),
    .A1(_01248_),
    .A2(_01283_),
    .A3(_01318_),
    .S1(net7831),
    .X(_02063_));
 sg13g2_nor2_1 _15644_ (.A(net7445),
    .B(_02063_),
    .Y(_02064_));
 sg13g2_nor2_1 _15645_ (.A(_02062_),
    .B(_02064_),
    .Y(_02065_));
 sg13g2_and4_1 _15646_ (.A(_02044_),
    .B(_02053_),
    .C(_02060_),
    .D(_02065_),
    .X(_02066_));
 sg13g2_nand4_1 _15647_ (.B(_02053_),
    .C(_02060_),
    .A(_02044_),
    .Y(_02067_),
    .D(_02065_));
 sg13g2_a221oi_1 _15648_ (.B2(net8006),
    .C1(_02035_),
    .B1(_02067_),
    .A1(net7354),
    .Y(_02068_),
    .A2(net7271));
 sg13g2_nand2_1 _15649_ (.Y(_02069_),
    .A(net6981),
    .B(_02032_));
 sg13g2_o21ai_1 _15650_ (.B1(_02069_),
    .Y(_02070_),
    .A1(_08251_),
    .A2(_02032_));
 sg13g2_o21ai_1 _15651_ (.B1(_02070_),
    .Y(_02071_),
    .A1(net7364),
    .A2(_02068_));
 sg13g2_mux4_1 _15652_ (.S0(net7776),
    .A0(_00797_),
    .A1(_00829_),
    .A2(_00861_),
    .A3(_00897_),
    .S1(net7728),
    .X(_02072_));
 sg13g2_and2_1 _15653_ (.A(_08255_),
    .B(_02072_),
    .X(_02073_));
 sg13g2_nand2_1 _15654_ (.Y(_02074_),
    .A(net7714),
    .B(_00765_));
 sg13g2_nand2b_1 _15655_ (.Y(_02075_),
    .B(_00637_),
    .A_N(net7714));
 sg13g2_a21oi_1 _15656_ (.A1(_02074_),
    .A2(_02075_),
    .Y(_02076_),
    .B1(net7600));
 sg13g2_nand3b_1 _15657_ (.B(net7775),
    .C(_00961_),
    .Y(_02077_),
    .A_N(net7726));
 sg13g2_nand3b_1 _15658_ (.B(_01313_),
    .C(net7726),
    .Y(_02078_),
    .A_N(net7775));
 sg13g2_a21oi_1 _15659_ (.A1(_02077_),
    .A2(_02078_),
    .Y(_02079_),
    .B1(net7598));
 sg13g2_nor4_1 _15660_ (.A(net7686),
    .B(_02073_),
    .C(_02076_),
    .D(_02079_),
    .Y(_02080_));
 sg13g2_inv_1 _15661_ (.Y(_02081_),
    .A(_01656_));
 sg13g2_mux4_1 _15662_ (.S0(net7776),
    .A0(_00932_),
    .A1(_00967_),
    .A2(_01002_),
    .A3(_01037_),
    .S1(net7727),
    .X(_02082_));
 sg13g2_mux2_1 _15663_ (.A0(_00669_),
    .A1(_00701_),
    .S(net7775),
    .X(_02083_));
 sg13g2_a221oi_1 _15664_ (.B2(net7518),
    .C1(net7695),
    .B1(_02083_),
    .A1(_00733_),
    .Y(_02084_),
    .A2(net7595));
 sg13g2_o21ai_1 _15665_ (.B1(net7713),
    .Y(_02085_),
    .A1(net7533),
    .A2(_02082_));
 sg13g2_o21ai_1 _15666_ (.B1(_02080_),
    .Y(_02086_),
    .A1(_02084_),
    .A2(_02085_));
 sg13g2_mux4_1 _15667_ (.S0(net7771),
    .A0(_01073_),
    .A1(_01108_),
    .A2(_01143_),
    .A3(_01178_),
    .S1(net7724),
    .X(_02087_));
 sg13g2_nor3_1 _15668_ (.A(net7712),
    .B(_08385_),
    .C(_02087_),
    .Y(_02088_));
 sg13g2_inv_1 _15669_ (.Y(_02089_),
    .A(_01651_));
 sg13g2_mux4_1 _15670_ (.S0(net7769),
    .A0(_01213_),
    .A1(_01249_),
    .A2(_01284_),
    .A3(_01319_),
    .S1(net7724),
    .X(_02090_));
 sg13g2_nor2_1 _15671_ (.A(net7588),
    .B(_02090_),
    .Y(_02091_));
 sg13g2_mux2_1 _15672_ (.A0(_01354_),
    .A1(_01389_),
    .S(net7768),
    .X(_02092_));
 sg13g2_nor3_1 _15673_ (.A(net7577),
    .B(_08503_),
    .C(_02092_),
    .Y(_02093_));
 sg13g2_mux2_1 _15674_ (.A0(_01425_),
    .A1(_01460_),
    .S(net7768),
    .X(_02094_));
 sg13g2_nor3_1 _15675_ (.A(net7577),
    .B(net7569),
    .C(_02094_),
    .Y(_02095_));
 sg13g2_mux2_1 _15676_ (.A0(_01495_),
    .A1(_01530_),
    .S(net7768),
    .X(_02096_));
 sg13g2_nor3_1 _15677_ (.A(net7577),
    .B(net7561),
    .C(_02096_),
    .Y(_02097_));
 sg13g2_inv_1 _15678_ (.Y(_02098_),
    .A(_01648_));
 sg13g2_mux2_1 _15679_ (.A0(_01565_),
    .A1(_00609_),
    .S(net7768),
    .X(_02099_));
 sg13g2_nor2_1 _15680_ (.A(net7556),
    .B(_02099_),
    .Y(_02100_));
 sg13g2_or4_1 _15681_ (.A(_02093_),
    .B(_02095_),
    .C(_02097_),
    .D(_02100_),
    .X(_02101_));
 sg13g2_nor3_1 _15682_ (.A(_02088_),
    .B(_02091_),
    .C(_02101_),
    .Y(_02102_));
 sg13g2_and2_1 _15683_ (.A(_02086_),
    .B(_02102_),
    .X(_02103_));
 sg13g2_inv_1 _15684_ (.Y(_02104_),
    .A(_02103_));
 sg13g2_a22oi_1 _15685_ (.Y(_02105_),
    .B1(_02103_),
    .B2(_08639_),
    .A2(_13410_),
    .A1(_01907_));
 sg13g2_mux2_1 _15686_ (.A0(_01313_),
    .A1(_00637_),
    .S(net7879),
    .X(_02106_));
 sg13g2_a22oi_1 _15687_ (.Y(_02107_),
    .B1(_02106_),
    .B2(net7833),
    .A2(net7527),
    .A1(_00961_));
 sg13g2_nand2b_1 _15688_ (.Y(_02108_),
    .B(net7879),
    .A_N(_00701_));
 sg13g2_o21ai_1 _15689_ (.B1(_02108_),
    .Y(_02109_),
    .A1(net7879),
    .A2(_00669_));
 sg13g2_mux2_1 _15690_ (.A0(_00733_),
    .A1(_00765_),
    .S(net7878),
    .X(_02110_));
 sg13g2_o21ai_1 _15691_ (.B1(net7530),
    .Y(_02111_),
    .A1(net7520),
    .A2(_02110_));
 sg13g2_a221oi_1 _15692_ (.B2(net7515),
    .C1(_02111_),
    .B1(_02109_),
    .A1(net7484),
    .Y(_02112_),
    .A2(_02107_));
 sg13g2_mux2_1 _15693_ (.A0(_01284_),
    .A1(_01319_),
    .S(net7864),
    .X(_02113_));
 sg13g2_nor2_1 _15694_ (.A(net7520),
    .B(_02113_),
    .Y(_02114_));
 sg13g2_mux2_1 _15695_ (.A0(_01073_),
    .A1(_01108_),
    .S(net7917),
    .X(_02115_));
 sg13g2_nor2_1 _15696_ (.A(_10182_),
    .B(_02115_),
    .Y(_02116_));
 sg13g2_mux2_1 _15697_ (.A0(_01143_),
    .A1(_01178_),
    .S(net7917),
    .X(_02117_));
 sg13g2_nor2_1 _15698_ (.A(net7460),
    .B(_02117_),
    .Y(_02118_));
 sg13g2_mux2_1 _15699_ (.A0(_01213_),
    .A1(_01249_),
    .S(net7864),
    .X(_02119_));
 sg13g2_o21ai_1 _15700_ (.B1(net7502),
    .Y(_02120_),
    .A1(net7504),
    .A2(_02119_));
 sg13g2_nor4_1 _15701_ (.A(_02114_),
    .B(_02116_),
    .C(_02118_),
    .D(_02120_),
    .Y(_02121_));
 sg13g2_mux2_1 _15702_ (.A0(_01354_),
    .A1(_01389_),
    .S(net7876),
    .X(_02122_));
 sg13g2_nand3_1 _15703_ (.B(_10179_),
    .C(_02122_),
    .A(net7497),
    .Y(_02123_));
 sg13g2_mux2_1 _15704_ (.A0(_01425_),
    .A1(_01460_),
    .S(net7876),
    .X(_02124_));
 sg13g2_nand3_1 _15705_ (.B(_10189_),
    .C(_02124_),
    .A(net7497),
    .Y(_02125_));
 sg13g2_mux2_1 _15706_ (.A0(_01495_),
    .A1(_01530_),
    .S(net7876),
    .X(_02126_));
 sg13g2_nand3_1 _15707_ (.B(net7497),
    .C(_02126_),
    .A(net7513),
    .Y(_02127_));
 sg13g2_mux2_1 _15708_ (.A0(_01565_),
    .A1(_00609_),
    .S(net7876),
    .X(_02128_));
 sg13g2_nand2_1 _15709_ (.Y(_02129_),
    .A(_10980_),
    .B(_02128_));
 sg13g2_mux2_1 _15710_ (.A0(_00861_),
    .A1(_00897_),
    .S(net7877),
    .X(_02130_));
 sg13g2_nand3_1 _15711_ (.B(_10189_),
    .C(_02130_),
    .A(net7545),
    .Y(_02131_));
 sg13g2_mux2_1 _15712_ (.A0(_00797_),
    .A1(_00829_),
    .S(net7877),
    .X(_02132_));
 sg13g2_nand3_1 _15713_ (.B(_10179_),
    .C(_02132_),
    .A(net7545),
    .Y(_02133_));
 sg13g2_mux2_1 _15714_ (.A0(_00932_),
    .A1(_00967_),
    .S(net7876),
    .X(_02134_));
 sg13g2_nand3_1 _15715_ (.B(net7513),
    .C(_02134_),
    .A(net7545),
    .Y(_02135_));
 sg13g2_mux2_1 _15716_ (.A0(_01002_),
    .A1(_01037_),
    .S(net7877),
    .X(_02136_));
 sg13g2_nand3_1 _15717_ (.B(net7526),
    .C(_02136_),
    .A(net7545),
    .Y(_02137_));
 sg13g2_nand4_1 _15718_ (.B(_02125_),
    .C(_02131_),
    .A(_02123_),
    .Y(_02138_),
    .D(_02133_));
 sg13g2_nand4_1 _15719_ (.B(_02129_),
    .C(_02135_),
    .A(_02127_),
    .Y(_02139_),
    .D(_02137_));
 sg13g2_nor4_1 _15720_ (.A(_02112_),
    .B(_02121_),
    .C(_02138_),
    .D(_02139_),
    .Y(_02140_));
 sg13g2_or4_1 _15721_ (.A(_02112_),
    .B(_02121_),
    .C(_02138_),
    .D(_02139_),
    .X(_02141_));
 sg13g2_nand2b_1 _15722_ (.Y(_02142_),
    .B(net8000),
    .A_N(_01642_));
 sg13g2_o21ai_1 _15723_ (.B1(_02142_),
    .Y(_02143_),
    .A1(_01672_),
    .A2(net7479));
 sg13g2_a221oi_1 _15724_ (.B2(net8006),
    .C1(_02143_),
    .B1(net7349),
    .A1(net7354),
    .Y(_02144_),
    .A2(_02104_));
 sg13g2_mux2_1 _15725_ (.A0(_08254_),
    .A1(net6981),
    .S(_02105_),
    .X(_02145_));
 sg13g2_o21ai_1 _15726_ (.B1(_02145_),
    .Y(_02146_),
    .A1(net7364),
    .A2(_02144_));
 sg13g2_mux4_1 _15727_ (.S0(net7753),
    .A0(_00798_),
    .A1(_00830_),
    .A2(_00863_),
    .A3(_00898_),
    .S1(net7735),
    .X(_02147_));
 sg13g2_nand2_1 _15728_ (.Y(_02148_),
    .A(net7606),
    .B(_02147_));
 sg13g2_mux2_1 _15729_ (.A0(_00638_),
    .A1(_00766_),
    .S(net7701),
    .X(_02149_));
 sg13g2_a21oi_1 _15730_ (.A1(_00972_),
    .A2(net7422),
    .Y(_02150_),
    .B1(net7685));
 sg13g2_a22oi_1 _15731_ (.Y(_02151_),
    .B1(_02149_),
    .B2(net7436),
    .A2(net7424),
    .A1(_01324_));
 sg13g2_mux4_1 _15732_ (.S0(net7753),
    .A0(_00933_),
    .A1(_00968_),
    .A2(_01003_),
    .A3(_01039_),
    .S1(net7735),
    .X(_02152_));
 sg13g2_mux2_1 _15733_ (.A0(_00670_),
    .A1(_00702_),
    .S(net7762),
    .X(_02153_));
 sg13g2_a22oi_1 _15734_ (.Y(_02154_),
    .B1(_02153_),
    .B2(_09011_),
    .A2(_08313_),
    .A1(_00734_));
 sg13g2_o21ai_1 _15735_ (.B1(net7701),
    .Y(_02155_),
    .A1(_08946_),
    .A2(_02152_));
 sg13g2_a21o_1 _15736_ (.A2(_02154_),
    .A1(_08946_),
    .B1(_02155_),
    .X(_02156_));
 sg13g2_nand4_1 _15737_ (.B(_02150_),
    .C(_02151_),
    .A(_02148_),
    .Y(_02157_),
    .D(_02156_));
 sg13g2_mux4_1 _15738_ (.S0(net7749),
    .A0(_01074_),
    .A1(_01109_),
    .A2(_01144_),
    .A3(_01179_),
    .S1(net7721),
    .X(_02158_));
 sg13g2_nand2b_1 _15739_ (.Y(_02159_),
    .B(net7433),
    .A_N(_02158_));
 sg13g2_mux4_1 _15740_ (.S0(net7752),
    .A0(_01215_),
    .A1(_01250_),
    .A2(_01285_),
    .A3(_01320_),
    .S1(net7718),
    .X(_02160_));
 sg13g2_or2_1 _15741_ (.X(_02161_),
    .B(_02160_),
    .A(net7586));
 sg13g2_mux2_1 _15742_ (.A0(_01567_),
    .A1(_00610_),
    .S(net7759),
    .X(_02162_));
 sg13g2_nor2_1 _15743_ (.A(net7553),
    .B(_02162_),
    .Y(_02163_));
 sg13g2_mux2_1 _15744_ (.A0(_01426_),
    .A1(_01461_),
    .S(net7754),
    .X(_02164_));
 sg13g2_nor3_1 _15745_ (.A(net7584),
    .B(net7568),
    .C(_02164_),
    .Y(_02165_));
 sg13g2_mux2_1 _15746_ (.A0(_01496_),
    .A1(_01531_),
    .S(net7754),
    .X(_02166_));
 sg13g2_nor3_1 _15747_ (.A(net7583),
    .B(net7565),
    .C(_02166_),
    .Y(_02167_));
 sg13g2_mux2_1 _15748_ (.A0(_01355_),
    .A1(_01391_),
    .S(net7754),
    .X(_02168_));
 sg13g2_nor3_1 _15749_ (.A(net7584),
    .B(net7560),
    .C(_02168_),
    .Y(_02169_));
 sg13g2_nor4_1 _15750_ (.A(_02163_),
    .B(_02165_),
    .C(_02167_),
    .D(_02169_),
    .Y(_02170_));
 sg13g2_and4_1 _15751_ (.A(_02157_),
    .B(_02159_),
    .C(_02161_),
    .D(_02170_),
    .X(_02171_));
 sg13g2_inv_1 _15752_ (.Y(_02172_),
    .A(net7033));
 sg13g2_a22oi_1 _15753_ (.Y(_02173_),
    .B1(_02171_),
    .B2(_08639_),
    .A2(net7039),
    .A1(_01909_));
 sg13g2_nor2b_1 _15754_ (.A(net6980),
    .B_N(_02173_),
    .Y(_02174_));
 sg13g2_mux2_1 _15755_ (.A0(_01567_),
    .A1(_00610_),
    .S(net7912),
    .X(_02175_));
 sg13g2_nor2_1 _15756_ (.A(net7448),
    .B(_02175_),
    .Y(_02176_));
 sg13g2_mux2_1 _15757_ (.A0(_01496_),
    .A1(_01531_),
    .S(net7903),
    .X(_02177_));
 sg13g2_nor3_1 _15758_ (.A(net7508),
    .B(net7489),
    .C(_02177_),
    .Y(_02178_));
 sg13g2_mux2_1 _15759_ (.A0(_00798_),
    .A1(_00830_),
    .S(net7856),
    .X(_02179_));
 sg13g2_nor3_1 _15760_ (.A(net7538),
    .B(net7467),
    .C(_02179_),
    .Y(_02180_));
 sg13g2_mux2_1 _15761_ (.A0(_00863_),
    .A1(_00898_),
    .S(net7856),
    .X(_02181_));
 sg13g2_nor3_1 _15762_ (.A(net7538),
    .B(net7458),
    .C(_02181_),
    .Y(_02182_));
 sg13g2_nor4_1 _15763_ (.A(_02176_),
    .B(_02178_),
    .C(_02180_),
    .D(_02182_),
    .Y(_02183_));
 sg13g2_mux2_1 _15764_ (.A0(_01003_),
    .A1(_01039_),
    .S(net7862),
    .X(_02184_));
 sg13g2_nor3_1 _15765_ (.A(net7538),
    .B(net7522),
    .C(_02184_),
    .Y(_02185_));
 sg13g2_mux2_1 _15766_ (.A0(_00933_),
    .A1(_00968_),
    .S(net7856),
    .X(_02186_));
 sg13g2_nor3_1 _15767_ (.A(net7538),
    .B(net7506),
    .C(_02186_),
    .Y(_02187_));
 sg13g2_mux2_1 _15768_ (.A0(_01355_),
    .A1(_01391_),
    .S(net7906),
    .X(_02188_));
 sg13g2_nor3_1 _15769_ (.A(net7488),
    .B(net7469),
    .C(_02188_),
    .Y(_02189_));
 sg13g2_mux2_1 _15770_ (.A0(_01426_),
    .A1(_01461_),
    .S(net7902),
    .X(_02190_));
 sg13g2_nor3_1 _15771_ (.A(net7488),
    .B(net7459),
    .C(_02190_),
    .Y(_02191_));
 sg13g2_nor4_1 _15772_ (.A(_02185_),
    .B(_02187_),
    .C(_02189_),
    .D(_02191_),
    .Y(_02192_));
 sg13g2_mux2_1 _15773_ (.A0(_01324_),
    .A1(_00638_),
    .S(net7842),
    .X(_02193_));
 sg13g2_and2_1 _15774_ (.A(net7842),
    .B(_00972_),
    .X(_02194_));
 sg13g2_mux2_1 _15775_ (.A0(_00670_),
    .A1(_00702_),
    .S(net7842),
    .X(_02195_));
 sg13g2_mux2_1 _15776_ (.A0(_00734_),
    .A1(_00766_),
    .S(net7842),
    .X(_02196_));
 sg13g2_mux4_1 _15777_ (.S0(net7813),
    .A0(_02194_),
    .A1(_02195_),
    .A2(_02193_),
    .A3(_02196_),
    .S1(net7821),
    .X(_02197_));
 sg13g2_or2_1 _15778_ (.X(_02198_),
    .B(_02197_),
    .A(net7528));
 sg13g2_mux4_1 _15779_ (.S0(net7900),
    .A0(_01074_),
    .A1(_01109_),
    .A2(_01144_),
    .A3(_01179_),
    .S1(net7818),
    .X(_02199_));
 sg13g2_nor3_1 _15780_ (.A(net7809),
    .B(net7499),
    .C(_02199_),
    .Y(_02200_));
 sg13g2_inv_1 _15781_ (.Y(_02201_),
    .A(net7981));
 sg13g2_mux4_1 _15782_ (.S0(net7897),
    .A0(_01215_),
    .A1(_01250_),
    .A2(_01285_),
    .A3(_01320_),
    .S1(net7818),
    .X(_02202_));
 sg13g2_nor2_1 _15783_ (.A(net7444),
    .B(_02202_),
    .Y(_02203_));
 sg13g2_nor2_1 _15784_ (.A(_02200_),
    .B(_02203_),
    .Y(_02204_));
 sg13g2_and4_1 _15785_ (.A(_02183_),
    .B(_02192_),
    .C(_02198_),
    .D(_02204_),
    .X(_02205_));
 sg13g2_nand4_1 _15786_ (.B(_02192_),
    .C(_02198_),
    .A(_02183_),
    .Y(_02206_),
    .D(_02204_));
 sg13g2_nand2b_1 _15787_ (.Y(_02207_),
    .B(net8000),
    .A_N(_01643_));
 sg13g2_o21ai_1 _15788_ (.B1(_02207_),
    .Y(_02208_),
    .A1(_01608_),
    .A2(net7479));
 sg13g2_a21oi_1 _15789_ (.A1(net8006),
    .A2(net7348),
    .Y(_02209_),
    .B1(_02208_));
 sg13g2_o21ai_1 _15790_ (.B1(_02209_),
    .Y(_02210_),
    .A1(_09277_),
    .A2(_02171_));
 sg13g2_inv_1 _15791_ (.Y(_02211_),
    .A(\cs_registers_i.nmi_mode_i ));
 sg13g2_a21oi_1 _15792_ (.A1(net7385),
    .A2(_02210_),
    .Y(_02212_),
    .B1(_02174_));
 sg13g2_o21ai_1 _15793_ (.B1(_02212_),
    .Y(_02213_),
    .A1(_08254_),
    .A2(_02173_));
 sg13g2_nand3_1 _15794_ (.B(_08800_),
    .C(_08808_),
    .A(net7748),
    .Y(_02214_));
 sg13g2_nand2b_1 _15795_ (.Y(_02215_),
    .B(_01915_),
    .A_N(_08785_));
 sg13g2_nand3_1 _15796_ (.B(_08665_),
    .C(_08784_),
    .A(net7677),
    .Y(_02216_));
 sg13g2_a21oi_1 _15797_ (.A1(_02215_),
    .A2(_02216_),
    .Y(_02217_),
    .B1(_08819_));
 sg13g2_nor2_1 _15798_ (.A(_08614_),
    .B(_02217_),
    .Y(_02218_));
 sg13g2_mux4_1 _15799_ (.S0(net7776),
    .A0(_00799_),
    .A1(_00831_),
    .A2(_00864_),
    .A3(_00899_),
    .S1(net7727),
    .X(_02219_));
 sg13g2_and2_1 _15800_ (.A(_08255_),
    .B(_02219_),
    .X(_02220_));
 sg13g2_nand2_1 _15801_ (.Y(_02221_),
    .A(net7713),
    .B(_00767_));
 sg13g2_nand2b_1 _15802_ (.Y(_02222_),
    .B(_00639_),
    .A_N(net7713));
 sg13g2_a21oi_1 _15803_ (.A1(_02221_),
    .A2(_02222_),
    .Y(_02223_),
    .B1(net7600));
 sg13g2_nand3b_1 _15804_ (.B(net7775),
    .C(_00983_),
    .Y(_02224_),
    .A_N(net7726));
 sg13g2_nand3b_1 _15805_ (.B(_01335_),
    .C(net7726),
    .Y(_02225_),
    .A_N(net7775));
 sg13g2_inv_1 _15806_ (.Y(_02226_),
    .A(net7984));
 sg13g2_a21oi_1 _15807_ (.A1(_02224_),
    .A2(_02225_),
    .Y(_02227_),
    .B1(net7598));
 sg13g2_nor4_1 _15808_ (.A(net7686),
    .B(_02220_),
    .C(_02223_),
    .D(_02227_),
    .Y(_02228_));
 sg13g2_mux4_1 _15809_ (.S0(net7776),
    .A0(_00934_),
    .A1(_00969_),
    .A2(_01004_),
    .A3(_01040_),
    .S1(net7727),
    .X(_02229_));
 sg13g2_mux2_1 _15810_ (.A0(_00671_),
    .A1(_00703_),
    .S(net7776),
    .X(_02230_));
 sg13g2_a221oi_1 _15811_ (.B2(net7518),
    .C1(net7695),
    .B1(_02230_),
    .A1(_00735_),
    .Y(_02231_),
    .A2(net7595));
 sg13g2_inv_1 _15812_ (.Y(_02232_),
    .A(\id_stage_i.controller_i.controller_run_o ));
 sg13g2_o21ai_1 _15813_ (.B1(net7713),
    .Y(_02233_),
    .A1(net7533),
    .A2(_02229_));
 sg13g2_o21ai_1 _15814_ (.B1(_02228_),
    .Y(_02234_),
    .A1(_02231_),
    .A2(_02233_));
 sg13g2_inv_1 _15815_ (.Y(_02235_),
    .A(_01605_));
 sg13g2_mux4_1 _15816_ (.S0(net7771),
    .A0(_01075_),
    .A1(_01110_),
    .A2(_01145_),
    .A3(_01180_),
    .S1(net7724),
    .X(_02236_));
 sg13g2_nand2b_1 _15817_ (.Y(_02237_),
    .B(_08387_),
    .A_N(_02236_));
 sg13g2_inv_1 _15818_ (.Y(_02238_),
    .A(net7986));
 sg13g2_mux4_1 _15819_ (.S0(net7769),
    .A0(_01216_),
    .A1(_01251_),
    .A2(_01286_),
    .A3(_01321_),
    .S1(net7728),
    .X(_02239_));
 sg13g2_or2_1 _15820_ (.X(_02240_),
    .B(_02239_),
    .A(net7588));
 sg13g2_mux2_1 _15821_ (.A0(_01356_),
    .A1(_01392_),
    .S(net7769),
    .X(_02241_));
 sg13g2_nor3_1 _15822_ (.A(net7578),
    .B(_08503_),
    .C(_02241_),
    .Y(_02242_));
 sg13g2_mux2_1 _15823_ (.A0(_01568_),
    .A1(_00611_),
    .S(net7771),
    .X(_02243_));
 sg13g2_nor2_1 _15824_ (.A(net7556),
    .B(_02243_),
    .Y(_02244_));
 sg13g2_inv_1 _15825_ (.Y(_02245_),
    .A(_01601_));
 sg13g2_mux2_1 _15826_ (.A0(_01427_),
    .A1(_01462_),
    .S(net7769),
    .X(_02246_));
 sg13g2_nor3_1 _15827_ (.A(net7578),
    .B(net7569),
    .C(_02246_),
    .Y(_02247_));
 sg13g2_mux2_1 _15828_ (.A0(_01497_),
    .A1(_01532_),
    .S(net7771),
    .X(_02248_));
 sg13g2_nor3_1 _15829_ (.A(net7578),
    .B(net7561),
    .C(_02248_),
    .Y(_02249_));
 sg13g2_nor4_1 _15830_ (.A(_02242_),
    .B(_02244_),
    .C(_02247_),
    .D(_02249_),
    .Y(_02250_));
 sg13g2_inv_1 _15831_ (.Y(_02251_),
    .A(_00006_));
 sg13g2_inv_1 _15832_ (.Y(_02252_),
    .A(net7269));
 sg13g2_nand4_1 _15833_ (.B(_02237_),
    .C(_02240_),
    .A(_02234_),
    .Y(_02253_),
    .D(_02250_));
 sg13g2_a221oi_1 _15834_ (.B2(_08614_),
    .C1(net7360),
    .B1(net7269),
    .A1(_02214_),
    .Y(_02254_),
    .A2(_02218_));
 sg13g2_mux4_1 _15835_ (.S0(net7864),
    .A0(_01356_),
    .A1(_01392_),
    .A2(_01427_),
    .A3(_01462_),
    .S1(net7830),
    .X(_02255_));
 sg13g2_or3_1 _15836_ (.A(net7814),
    .B(net7490),
    .C(_02255_),
    .X(_02256_));
 sg13g2_mux4_1 _15837_ (.S0(net7917),
    .A0(_01497_),
    .A1(_01532_),
    .A2(_01568_),
    .A3(_00611_),
    .S1(net7830),
    .X(_02257_));
 sg13g2_o21ai_1 _15838_ (.B1(_02256_),
    .Y(_02258_),
    .A1(_10018_),
    .A2(_02257_));
 sg13g2_mux2_1 _15839_ (.A0(_00671_),
    .A1(_00703_),
    .S(net7878),
    .X(_02259_));
 sg13g2_mux2_1 _15840_ (.A0(_00735_),
    .A1(_00767_),
    .S(net7878),
    .X(_02260_));
 sg13g2_mux2_1 _15841_ (.A0(_01335_),
    .A1(_00639_),
    .S(net7878),
    .X(_02261_));
 sg13g2_and2_1 _15842_ (.A(net7878),
    .B(_00983_),
    .X(_02262_));
 sg13g2_mux4_1 _15843_ (.S0(net7833),
    .A0(_02259_),
    .A1(_02260_),
    .A2(_02262_),
    .A3(_02261_),
    .S1(net7484),
    .X(_02263_));
 sg13g2_nor2_1 _15844_ (.A(net7529),
    .B(_02263_),
    .Y(_02264_));
 sg13g2_mux4_1 _15845_ (.S0(net7917),
    .A0(_01075_),
    .A1(_01110_),
    .A2(_01145_),
    .A3(_01180_),
    .S1(net7830),
    .X(_02265_));
 sg13g2_mux4_1 _15846_ (.S0(net7864),
    .A0(_01216_),
    .A1(_01251_),
    .A2(_01286_),
    .A3(_01321_),
    .S1(net7830),
    .X(_02266_));
 sg13g2_or2_1 _15847_ (.X(_02267_),
    .B(_02266_),
    .A(net7445));
 sg13g2_o21ai_1 _15848_ (.B1(_02267_),
    .Y(_02268_),
    .A1(net7421),
    .A2(_02265_));
 sg13g2_nand2_1 _15849_ (.Y(_02269_),
    .A(net7869),
    .B(_01040_));
 sg13g2_nand2b_1 _15850_ (.Y(_02270_),
    .B(_01004_),
    .A_N(net7869));
 sg13g2_nand4_1 _15851_ (.B(net7526),
    .C(_02269_),
    .A(net7545),
    .Y(_02271_),
    .D(_02270_));
 sg13g2_nand2_1 _15852_ (.Y(_02272_),
    .A(net7869),
    .B(_00899_));
 sg13g2_nand2b_1 _15853_ (.Y(_02273_),
    .B(_00864_),
    .A_N(net7869));
 sg13g2_nand4_1 _15854_ (.B(_10189_),
    .C(_02272_),
    .A(net7544),
    .Y(_02274_),
    .D(_02273_));
 sg13g2_nand2_1 _15855_ (.Y(_02275_),
    .A(net7869),
    .B(_00831_));
 sg13g2_nand2b_1 _15856_ (.Y(_02276_),
    .B(_00799_),
    .A_N(net7869));
 sg13g2_nand4_1 _15857_ (.B(_10179_),
    .C(_02275_),
    .A(net7545),
    .Y(_02277_),
    .D(_02276_));
 sg13g2_nand2_1 _15858_ (.Y(_02278_),
    .A(net7869),
    .B(_00969_));
 sg13g2_nand2b_1 _15859_ (.Y(_02279_),
    .B(_00934_),
    .A_N(net7869));
 sg13g2_nand4_1 _15860_ (.B(net7513),
    .C(_02278_),
    .A(net7545),
    .Y(_02280_),
    .D(_02279_));
 sg13g2_nand4_1 _15861_ (.B(_02274_),
    .C(_02277_),
    .A(_02271_),
    .Y(_02281_),
    .D(_02280_));
 sg13g2_nor4_1 _15862_ (.A(_02258_),
    .B(_02264_),
    .C(_02268_),
    .D(_02281_),
    .Y(_02282_));
 sg13g2_or4_1 _15863_ (.A(_02258_),
    .B(_02264_),
    .C(_02268_),
    .D(_02281_),
    .X(_02283_));
 sg13g2_nand2b_1 _15864_ (.Y(_02284_),
    .B(net8000),
    .A_N(_01644_));
 sg13g2_o21ai_1 _15865_ (.B1(_02284_),
    .Y(_02285_),
    .A1(_01609_),
    .A2(net7479));
 sg13g2_a221oi_1 _15866_ (.B2(net8006),
    .C1(_02285_),
    .B1(_02283_),
    .A1(net7354),
    .Y(_02286_),
    .A2(net7269));
 sg13g2_nor2_1 _15867_ (.A(net7364),
    .B(_02286_),
    .Y(_02287_));
 sg13g2_a21oi_1 _15868_ (.A1(_08251_),
    .A2(_02254_),
    .Y(_02288_),
    .B1(_02287_));
 sg13g2_o21ai_1 _15869_ (.B1(_02288_),
    .Y(_02289_),
    .A1(net6980),
    .A2(_02254_));
 sg13g2_and2_1 _15870_ (.A(_08777_),
    .B(_08797_),
    .X(_02290_));
 sg13g2_nor2_1 _15871_ (.A(_08819_),
    .B(net7268),
    .Y(_02291_));
 sg13g2_a21oi_1 _15872_ (.A1(net7677),
    .A2(_02291_),
    .Y(_02292_),
    .B1(_08614_));
 sg13g2_a21o_1 _15873_ (.A2(_08808_),
    .A1(_08800_),
    .B1(_02290_),
    .X(_02293_));
 sg13g2_nand2_1 _15874_ (.Y(_02294_),
    .A(net7930),
    .B(_02293_));
 sg13g2_mux2_1 _15875_ (.A0(_01498_),
    .A1(_01534_),
    .S(net7786),
    .X(_02295_));
 sg13g2_nor3_1 _15876_ (.A(net7574),
    .B(net7562),
    .C(_02295_),
    .Y(_02296_));
 sg13g2_mux2_1 _15877_ (.A0(_01428_),
    .A1(_01463_),
    .S(net7786),
    .X(_02297_));
 sg13g2_nor3_1 _15878_ (.A(net7574),
    .B(net7571),
    .C(_02297_),
    .Y(_02298_));
 sg13g2_mux2_1 _15879_ (.A0(_01569_),
    .A1(_00612_),
    .S(net7786),
    .X(_02299_));
 sg13g2_nor2_1 _15880_ (.A(net7556),
    .B(_02299_),
    .Y(_02300_));
 sg13g2_mux2_1 _15881_ (.A0(_01358_),
    .A1(_01393_),
    .S(net7786),
    .X(_02301_));
 sg13g2_nor3_1 _15882_ (.A(net7574),
    .B(net7558),
    .C(_02301_),
    .Y(_02302_));
 sg13g2_or4_1 _15883_ (.A(_02296_),
    .B(_02298_),
    .C(_02300_),
    .D(_02302_),
    .X(_02303_));
 sg13g2_mux4_1 _15884_ (.S0(net7787),
    .A0(_01217_),
    .A1(_01252_),
    .A2(_01287_),
    .A3(_01322_),
    .S1(net7727),
    .X(_02304_));
 sg13g2_mux4_1 _15885_ (.S0(net7786),
    .A0(_01076_),
    .A1(_01111_),
    .A2(_01146_),
    .A3(_01182_),
    .S1(net7727),
    .X(_02305_));
 sg13g2_nand2b_1 _15886_ (.Y(_02306_),
    .B(net7713),
    .A_N(_02304_));
 sg13g2_o21ai_1 _15887_ (.B1(_02306_),
    .Y(_02307_),
    .A1(net7713),
    .A2(_02305_));
 sg13g2_a21oi_1 _15888_ (.A1(net7591),
    .A2(_02307_),
    .Y(_02308_),
    .B1(_02303_));
 sg13g2_mux4_1 _15889_ (.S0(net7787),
    .A0(_00800_),
    .A1(_00832_),
    .A2(_00865_),
    .A3(_00900_),
    .S1(net7745),
    .X(_02309_));
 sg13g2_and2_1 _15890_ (.A(net7602),
    .B(_02309_),
    .X(_02310_));
 sg13g2_nand2_1 _15891_ (.Y(_02311_),
    .A(net7711),
    .B(_00768_));
 sg13g2_nand2b_1 _15892_ (.Y(_02312_),
    .B(_00640_),
    .A_N(net7711));
 sg13g2_a21oi_1 _15893_ (.A1(_02311_),
    .A2(_02312_),
    .Y(_02313_),
    .B1(net7600));
 sg13g2_nand3b_1 _15894_ (.B(net7783),
    .C(_00994_),
    .Y(_02314_),
    .A_N(net7747));
 sg13g2_nand3b_1 _15895_ (.B(_01346_),
    .C(net7747),
    .Y(_02315_),
    .A_N(net7783));
 sg13g2_a21oi_1 _15896_ (.A1(_02314_),
    .A2(_02315_),
    .Y(_02316_),
    .B1(net7598));
 sg13g2_nor4_1 _15897_ (.A(net7690),
    .B(_02310_),
    .C(_02313_),
    .D(_02316_),
    .Y(_02317_));
 sg13g2_mux4_1 _15898_ (.S0(net7784),
    .A0(_00935_),
    .A1(_00970_),
    .A2(_01006_),
    .A3(_01041_),
    .S1(net7745),
    .X(_02318_));
 sg13g2_nand2b_1 _15899_ (.Y(_02319_),
    .B(net7695),
    .A_N(_02318_));
 sg13g2_mux2_1 _15900_ (.A0(_00672_),
    .A1(_00704_),
    .S(net7774),
    .X(_02320_));
 sg13g2_a221oi_1 _15901_ (.B2(net7518),
    .C1(net7695),
    .B1(_02320_),
    .A1(_00736_),
    .Y(_02321_),
    .A2(net7595));
 sg13g2_nand3b_1 _15902_ (.B(net7711),
    .C(_02319_),
    .Y(_02322_),
    .A_N(_02321_));
 sg13g2_nand2_1 _15903_ (.Y(_02323_),
    .A(_02317_),
    .B(_02322_));
 sg13g2_a221oi_1 _15904_ (.B2(_02322_),
    .C1(_02303_),
    .B1(_02317_),
    .A1(net7591),
    .Y(_02324_),
    .A2(_02307_));
 sg13g2_nand2_1 _15905_ (.Y(_02325_),
    .A(_02308_),
    .B(_02323_));
 sg13g2_a221oi_1 _15906_ (.B2(net7363),
    .C1(net7361),
    .B1(_02325_),
    .A1(_02292_),
    .Y(_02326_),
    .A2(_02294_));
 sg13g2_mux2_1 _15907_ (.A0(_01346_),
    .A1(_00640_),
    .S(net7868),
    .X(_02327_));
 sg13g2_a221oi_1 _15908_ (.B2(net7833),
    .C1(net7815),
    .B1(_02327_),
    .A1(_00994_),
    .Y(_02328_),
    .A2(net7527));
 sg13g2_mux2_1 _15909_ (.A0(_00736_),
    .A1(_00768_),
    .S(net7868),
    .X(_02329_));
 sg13g2_nor2_1 _15910_ (.A(net7520),
    .B(_02329_),
    .Y(_02330_));
 sg13g2_mux2_1 _15911_ (.A0(_00672_),
    .A1(_00704_),
    .S(net7871),
    .X(_02331_));
 sg13g2_o21ai_1 _15912_ (.B1(net7530),
    .Y(_02332_),
    .A1(net7509),
    .A2(_02331_));
 sg13g2_or3_1 _15913_ (.A(_02328_),
    .B(_02330_),
    .C(_02332_),
    .X(_02333_));
 sg13g2_mux2_1 _15914_ (.A0(_01287_),
    .A1(_01322_),
    .S(net7870),
    .X(_02334_));
 sg13g2_nor2_1 _15915_ (.A(net7520),
    .B(_02334_),
    .Y(_02335_));
 sg13g2_mux2_1 _15916_ (.A0(_01076_),
    .A1(_01111_),
    .S(net7870),
    .X(_02336_));
 sg13g2_nor2_1 _15917_ (.A(net7465),
    .B(_02336_),
    .Y(_02337_));
 sg13g2_mux2_1 _15918_ (.A0(_01146_),
    .A1(_01182_),
    .S(net7870),
    .X(_02338_));
 sg13g2_nor2_1 _15919_ (.A(net7456),
    .B(_02338_),
    .Y(_02339_));
 sg13g2_mux2_1 _15920_ (.A0(_01217_),
    .A1(_01252_),
    .S(net7870),
    .X(_02340_));
 sg13g2_o21ai_1 _15921_ (.B1(net7501),
    .Y(_02341_),
    .A1(net7509),
    .A2(_02340_));
 sg13g2_or4_1 _15922_ (.A(_02335_),
    .B(_02337_),
    .C(_02339_),
    .D(_02341_),
    .X(_02342_));
 sg13g2_mux2_1 _15923_ (.A0(_01569_),
    .A1(_00612_),
    .S(net7872),
    .X(_02343_));
 sg13g2_nand2_1 _15924_ (.Y(_02344_),
    .A(net7450),
    .B(_02343_));
 sg13g2_mux2_1 _15925_ (.A0(_01498_),
    .A1(_01534_),
    .S(net7872),
    .X(_02345_));
 sg13g2_nand3_1 _15926_ (.B(net7493),
    .C(_02345_),
    .A(net7514),
    .Y(_02346_));
 sg13g2_mux2_1 _15927_ (.A0(_01428_),
    .A1(_01463_),
    .S(net7872),
    .X(_02347_));
 sg13g2_nand3_1 _15928_ (.B(net7463),
    .C(_02347_),
    .A(net7493),
    .Y(_02348_));
 sg13g2_mux2_1 _15929_ (.A0(_01358_),
    .A1(_01393_),
    .S(net7872),
    .X(_02349_));
 sg13g2_nand3_1 _15930_ (.B(net7472),
    .C(_02349_),
    .A(net7493),
    .Y(_02350_));
 sg13g2_mux2_1 _15931_ (.A0(_00865_),
    .A1(_00900_),
    .S(net7872),
    .X(_02351_));
 sg13g2_nand3_1 _15932_ (.B(net7463),
    .C(_02351_),
    .A(net7543),
    .Y(_02352_));
 sg13g2_mux2_1 _15933_ (.A0(_00800_),
    .A1(_00832_),
    .S(net7872),
    .X(_02353_));
 sg13g2_nand3_1 _15934_ (.B(net7472),
    .C(_02353_),
    .A(net7543),
    .Y(_02354_));
 sg13g2_mux2_1 _15935_ (.A0(_00935_),
    .A1(_00970_),
    .S(net7875),
    .X(_02355_));
 sg13g2_nand3_1 _15936_ (.B(net7514),
    .C(_02355_),
    .A(net7543),
    .Y(_02356_));
 sg13g2_mux2_1 _15937_ (.A0(_01006_),
    .A1(_01041_),
    .S(net7875),
    .X(_02357_));
 sg13g2_nand3_1 _15938_ (.B(net7526),
    .C(_02357_),
    .A(net7543),
    .Y(_02358_));
 sg13g2_and4_1 _15939_ (.A(_02344_),
    .B(_02348_),
    .C(_02350_),
    .D(_02356_),
    .X(_02359_));
 sg13g2_and4_1 _15940_ (.A(_02346_),
    .B(_02352_),
    .C(_02354_),
    .D(_02358_),
    .X(_02360_));
 sg13g2_and4_1 _15941_ (.A(_02333_),
    .B(_02342_),
    .C(_02359_),
    .D(_02360_),
    .X(_02361_));
 sg13g2_nand4_1 _15942_ (.B(_02342_),
    .C(_02359_),
    .A(_02333_),
    .Y(_02362_),
    .D(_02360_));
 sg13g2_nand2b_1 _15943_ (.Y(_02363_),
    .B(net8000),
    .A_N(_01645_));
 sg13g2_o21ai_1 _15944_ (.B1(_02363_),
    .Y(_02364_),
    .A1(_01610_),
    .A2(net7480));
 sg13g2_a221oi_1 _15945_ (.B2(net8007),
    .C1(_02364_),
    .B1(_02361_),
    .A1(net7354),
    .Y(_02365_),
    .A2(net7266));
 sg13g2_nor2_1 _15946_ (.A(net7375),
    .B(_02365_),
    .Y(_02366_));
 sg13g2_a21oi_1 _15947_ (.A1(net6919),
    .A2(_02326_),
    .Y(_02367_),
    .B1(_02366_));
 sg13g2_o21ai_1 _15948_ (.B1(_02367_),
    .Y(_02368_),
    .A1(net6980),
    .A2(_02326_));
 sg13g2_nand2_1 _15949_ (.Y(_02369_),
    .A(net7926),
    .B(_02293_));
 sg13g2_mux2_1 _15950_ (.A0(_01359_),
    .A1(_01394_),
    .S(net7801),
    .X(_02370_));
 sg13g2_nor3_1 _15951_ (.A(net7572),
    .B(net7558),
    .C(_02370_),
    .Y(_02371_));
 sg13g2_mux2_1 _15952_ (.A0(_01499_),
    .A1(_01535_),
    .S(net7801),
    .X(_02372_));
 sg13g2_nor3_1 _15953_ (.A(net7572),
    .B(net7562),
    .C(_02372_),
    .Y(_02373_));
 sg13g2_mux2_1 _15954_ (.A0(_01429_),
    .A1(_01464_),
    .S(net7801),
    .X(_02374_));
 sg13g2_nor3_1 _15955_ (.A(net7572),
    .B(net7571),
    .C(_02374_),
    .Y(_02375_));
 sg13g2_mux2_1 _15956_ (.A0(_01570_),
    .A1(_00613_),
    .S(net7801),
    .X(_02376_));
 sg13g2_nor2_1 _15957_ (.A(net7555),
    .B(_02376_),
    .Y(_02377_));
 sg13g2_or4_1 _15958_ (.A(_02371_),
    .B(_02373_),
    .C(_02375_),
    .D(_02377_),
    .X(_02378_));
 sg13g2_mux4_1 _15959_ (.S0(net7801),
    .A0(_01218_),
    .A1(_01253_),
    .A2(_01288_),
    .A3(_01323_),
    .S1(net7746),
    .X(_02379_));
 sg13g2_mux4_1 _15960_ (.S0(net7801),
    .A0(_01077_),
    .A1(_01112_),
    .A2(_01147_),
    .A3(_01183_),
    .S1(net7746),
    .X(_02380_));
 sg13g2_nand2b_1 _15961_ (.Y(_02381_),
    .B(net7709),
    .A_N(_02379_));
 sg13g2_o21ai_1 _15962_ (.B1(_02381_),
    .Y(_02382_),
    .A1(net7709),
    .A2(_02380_));
 sg13g2_a21oi_1 _15963_ (.A1(net7591),
    .A2(_02382_),
    .Y(_02383_),
    .B1(_02378_));
 sg13g2_mux4_1 _15964_ (.S0(net7799),
    .A0(_00801_),
    .A1(_00833_),
    .A2(_00866_),
    .A3(_00901_),
    .S1(net7746),
    .X(_02384_));
 sg13g2_and2_1 _15965_ (.A(net7602),
    .B(_02384_),
    .X(_02385_));
 sg13g2_nand2_1 _15966_ (.Y(_02386_),
    .A(net7710),
    .B(_00769_));
 sg13g2_nand2b_1 _15967_ (.Y(_02387_),
    .B(_00641_),
    .A_N(net7710));
 sg13g2_a21oi_1 _15968_ (.A1(_02386_),
    .A2(_02387_),
    .Y(_02388_),
    .B1(net7600));
 sg13g2_nand3b_1 _15969_ (.B(net7799),
    .C(_01005_),
    .Y(_02389_),
    .A_N(net7747));
 sg13g2_nand3b_1 _15970_ (.B(_01357_),
    .C(net7747),
    .Y(_02390_),
    .A_N(net7799));
 sg13g2_a21oi_1 _15971_ (.A1(_02389_),
    .A2(_02390_),
    .Y(_02391_),
    .B1(net7598));
 sg13g2_nor4_1 _15972_ (.A(net7690),
    .B(_02385_),
    .C(_02388_),
    .D(_02391_),
    .Y(_02392_));
 sg13g2_mux4_1 _15973_ (.S0(net7799),
    .A0(_00936_),
    .A1(_00971_),
    .A2(_01007_),
    .A3(_01042_),
    .S1(net7746),
    .X(_02393_));
 sg13g2_nand2b_1 _15974_ (.Y(_02394_),
    .B(net7694),
    .A_N(_02393_));
 sg13g2_mux2_1 _15975_ (.A0(_00673_),
    .A1(_00705_),
    .S(net7800),
    .X(_02395_));
 sg13g2_a221oi_1 _15976_ (.B2(net7516),
    .C1(net7694),
    .B1(_02395_),
    .A1(_00737_),
    .Y(_02396_),
    .A2(net7595));
 sg13g2_nand3b_1 _15977_ (.B(net7710),
    .C(_02394_),
    .Y(_02397_),
    .A_N(_02396_));
 sg13g2_nand2_1 _15978_ (.Y(_02398_),
    .A(_02392_),
    .B(_02397_));
 sg13g2_a221oi_1 _15979_ (.B2(_02397_),
    .C1(_02378_),
    .B1(_02392_),
    .A1(net7591),
    .Y(_02399_),
    .A2(_02382_));
 sg13g2_nand2_1 _15980_ (.Y(_02400_),
    .A(_02383_),
    .B(_02398_));
 sg13g2_a221oi_1 _15981_ (.B2(net7363),
    .C1(net7361),
    .B1(_02400_),
    .A1(_02292_),
    .Y(_02401_),
    .A2(_02369_));
 sg13g2_nand2b_1 _15982_ (.Y(_02402_),
    .B(_01570_),
    .A_N(net7889));
 sg13g2_nand2_1 _15983_ (.Y(_02403_),
    .A(net7889),
    .B(_00613_));
 sg13g2_nand3_1 _15984_ (.B(_02402_),
    .C(_02403_),
    .A(net7450),
    .Y(_02404_));
 sg13g2_nand2_1 _15985_ (.Y(_02405_),
    .A(net7891),
    .B(_01535_));
 sg13g2_nand2b_1 _15986_ (.Y(_02406_),
    .B(_01499_),
    .A_N(net7891));
 sg13g2_nand4_1 _15987_ (.B(net7495),
    .C(_02405_),
    .A(net7514),
    .Y(_02407_),
    .D(_02406_));
 sg13g2_nand2_1 _15988_ (.Y(_02408_),
    .A(net7886),
    .B(_01042_));
 sg13g2_nand2b_1 _15989_ (.Y(_02409_),
    .B(_01007_),
    .A_N(net7886));
 sg13g2_nand4_1 _15990_ (.B(net7525),
    .C(_02408_),
    .A(net7549),
    .Y(_02410_),
    .D(_02409_));
 sg13g2_nand2_1 _15991_ (.Y(_02411_),
    .A(net7886),
    .B(_00971_));
 sg13g2_nand2b_1 _15992_ (.Y(_02412_),
    .B(_00936_),
    .A_N(net7886));
 sg13g2_nand4_1 _15993_ (.B(net7514),
    .C(_02411_),
    .A(net7549),
    .Y(_02413_),
    .D(_02412_));
 sg13g2_nand2_1 _15994_ (.Y(_02414_),
    .A(net7886),
    .B(_00833_));
 sg13g2_nand2b_1 _15995_ (.Y(_02415_),
    .B(_00801_),
    .A_N(net7886));
 sg13g2_nand4_1 _15996_ (.B(net7472),
    .C(_02414_),
    .A(net7549),
    .Y(_02416_),
    .D(_02415_));
 sg13g2_nand2_1 _15997_ (.Y(_02417_),
    .A(net7890),
    .B(_00901_));
 sg13g2_nand2b_1 _15998_ (.Y(_02418_),
    .B(_00866_),
    .A_N(net7891));
 sg13g2_nand4_1 _15999_ (.B(net7463),
    .C(_02417_),
    .A(net7549),
    .Y(_02419_),
    .D(_02418_));
 sg13g2_nand2_1 _16000_ (.Y(_02420_),
    .A(net7889),
    .B(_01394_));
 sg13g2_nand2b_1 _16001_ (.Y(_02421_),
    .B(_01359_),
    .A_N(net7889));
 sg13g2_nand4_1 _16002_ (.B(net7472),
    .C(_02420_),
    .A(net7493),
    .Y(_02422_),
    .D(_02421_));
 sg13g2_nand2_1 _16003_ (.Y(_02423_),
    .A(net7889),
    .B(_01464_));
 sg13g2_nand2b_1 _16004_ (.Y(_02424_),
    .B(_01429_),
    .A_N(net7888));
 sg13g2_nand4_1 _16005_ (.B(net7463),
    .C(_02423_),
    .A(net7493),
    .Y(_02425_),
    .D(_02424_));
 sg13g2_nand4_1 _16006_ (.B(_02416_),
    .C(_02422_),
    .A(_02410_),
    .Y(_02426_),
    .D(_02425_));
 sg13g2_nand4_1 _16007_ (.B(_02407_),
    .C(_02413_),
    .A(_02404_),
    .Y(_02427_),
    .D(_02419_));
 sg13g2_mux2_1 _16008_ (.A0(_01357_),
    .A1(_00641_),
    .S(net7885),
    .X(_02428_));
 sg13g2_and2_1 _16009_ (.A(net7885),
    .B(_01005_),
    .X(_02429_));
 sg13g2_mux2_1 _16010_ (.A0(_00673_),
    .A1(_00705_),
    .S(net7884),
    .X(_02430_));
 sg13g2_mux2_1 _16011_ (.A0(_00737_),
    .A1(_00769_),
    .S(net7885),
    .X(_02431_));
 sg13g2_mux4_1 _16012_ (.S0(net7815),
    .A0(_02429_),
    .A1(_02430_),
    .A2(_02428_),
    .A3(_02431_),
    .S1(net7824),
    .X(_02432_));
 sg13g2_nor2_1 _16013_ (.A(net7529),
    .B(_02432_),
    .Y(_02433_));
 sg13g2_mux4_1 _16014_ (.S0(net7888),
    .A0(_01077_),
    .A1(_01112_),
    .A2(_01147_),
    .A3(_01183_),
    .S1(net7824),
    .X(_02434_));
 sg13g2_mux4_1 _16015_ (.S0(net7888),
    .A0(_01218_),
    .A1(_01253_),
    .A2(_01288_),
    .A3(_01323_),
    .S1(net7824),
    .X(_02435_));
 sg13g2_or2_1 _16016_ (.X(_02436_),
    .B(_02435_),
    .A(net7443));
 sg13g2_o21ai_1 _16017_ (.B1(_02436_),
    .Y(_02437_),
    .A1(net7421),
    .A2(_02434_));
 sg13g2_nor4_1 _16018_ (.A(_02426_),
    .B(_02427_),
    .C(_02433_),
    .D(_02437_),
    .Y(_02438_));
 sg13g2_or4_1 _16019_ (.A(_02426_),
    .B(_02427_),
    .C(_02433_),
    .D(_02437_),
    .X(_02439_));
 sg13g2_nand2b_1 _16020_ (.Y(_02440_),
    .B(net8001),
    .A_N(_01646_));
 sg13g2_o21ai_1 _16021_ (.B1(_02440_),
    .Y(_02441_),
    .A1(_01611_),
    .A2(net7478));
 sg13g2_a221oi_1 _16022_ (.B2(net8007),
    .C1(_02441_),
    .B1(_02439_),
    .A1(_09275_),
    .Y(_02442_),
    .A2(net7265));
 sg13g2_nor2_1 _16023_ (.A(net7375),
    .B(_02442_),
    .Y(_02443_));
 sg13g2_a21oi_1 _16024_ (.A1(net6918),
    .A2(_02401_),
    .Y(_02444_),
    .B1(_02443_));
 sg13g2_o21ai_1 _16025_ (.B1(_02444_),
    .Y(_02445_),
    .A1(net6978),
    .A2(_02401_));
 sg13g2_nand2_1 _16026_ (.Y(_02446_),
    .A(net7924),
    .B(_02293_));
 sg13g2_mux2_1 _16027_ (.A0(_01571_),
    .A1(_00614_),
    .S(net7770),
    .X(_02447_));
 sg13g2_nor2_1 _16028_ (.A(net7551),
    .B(_02447_),
    .Y(_02448_));
 sg13g2_mux2_1 _16029_ (.A0(_01430_),
    .A1(_01465_),
    .S(net7767),
    .X(_02449_));
 sg13g2_nor3_1 _16030_ (.A(net7579),
    .B(net7567),
    .C(_02449_),
    .Y(_02450_));
 sg13g2_mux2_1 _16031_ (.A0(_01360_),
    .A1(_01395_),
    .S(net7767),
    .X(_02451_));
 sg13g2_nor3_1 _16032_ (.A(net7579),
    .B(net7559),
    .C(_02451_),
    .Y(_02452_));
 sg13g2_mux2_1 _16033_ (.A0(_01501_),
    .A1(_01536_),
    .S(net7767),
    .X(_02453_));
 sg13g2_nor3_1 _16034_ (.A(net7579),
    .B(net7563),
    .C(_02453_),
    .Y(_02454_));
 sg13g2_or4_1 _16035_ (.A(_02448_),
    .B(_02450_),
    .C(_02452_),
    .D(_02454_),
    .X(_02455_));
 sg13g2_mux4_1 _16036_ (.S0(net7766),
    .A0(_01219_),
    .A1(_01254_),
    .A2(_01289_),
    .A3(_01325_),
    .S1(net7723),
    .X(_02456_));
 sg13g2_mux4_1 _16037_ (.S0(net7766),
    .A0(_01078_),
    .A1(_01113_),
    .A2(_01149_),
    .A3(_01184_),
    .S1(net7723),
    .X(_02457_));
 sg13g2_nand2b_1 _16038_ (.Y(_02458_),
    .B(net7703),
    .A_N(_02456_));
 sg13g2_o21ai_1 _16039_ (.B1(_02458_),
    .Y(_02459_),
    .A1(net7703),
    .A2(_02457_));
 sg13g2_a21o_1 _16040_ (.A2(_02459_),
    .A1(net7590),
    .B1(_02455_),
    .X(_02460_));
 sg13g2_mux4_1 _16041_ (.S0(net7770),
    .A0(_00937_),
    .A1(_00973_),
    .A2(_01008_),
    .A3(_01043_),
    .S1(net7723),
    .X(_02461_));
 sg13g2_and2_1 _16042_ (.A(_01901_),
    .B(net7706),
    .X(_02462_));
 sg13g2_and2_1 _16043_ (.A(_02461_),
    .B(net7640),
    .X(_02463_));
 sg13g2_mux4_1 _16044_ (.S0(net7765),
    .A0(_00802_),
    .A1(_00834_),
    .A2(_00867_),
    .A3(_00902_),
    .S1(net7725),
    .X(_02464_));
 sg13g2_and3_1 _16045_ (.X(_02465_),
    .A(_01016_),
    .B(net7599),
    .C(net7597));
 sg13g2_nand2_1 _16046_ (.Y(_02466_),
    .A(net7703),
    .B(_00770_));
 sg13g2_nand2b_1 _16047_ (.Y(_02467_),
    .B(_00642_),
    .A_N(net7703));
 sg13g2_a21oi_1 _16048_ (.A1(_02466_),
    .A2(_02467_),
    .Y(_02468_),
    .B1(net7601));
 sg13g2_and3_1 _16049_ (.X(_02469_),
    .A(_01368_),
    .B(net7599),
    .C(net7594));
 sg13g2_nor4_1 _16050_ (.A(net7687),
    .B(_02465_),
    .C(_02468_),
    .D(_02469_),
    .Y(_02470_));
 sg13g2_mux2_1 _16051_ (.A0(_00674_),
    .A1(_00706_),
    .S(net7765),
    .X(_02471_));
 sg13g2_nor2b_1 _16052_ (.A(net7765),
    .B_N(_00738_),
    .Y(_02472_));
 sg13g2_mux2_1 _16053_ (.A0(_02471_),
    .A1(_02472_),
    .S(net7725),
    .X(_02473_));
 sg13g2_a221oi_1 _16054_ (.B2(net7442),
    .C1(_02463_),
    .B1(_02473_),
    .A1(net7605),
    .Y(_02474_),
    .A2(_02464_));
 sg13g2_a221oi_1 _16055_ (.B2(_02474_),
    .C1(_02455_),
    .B1(_02470_),
    .A1(net7590),
    .Y(_02475_),
    .A2(_02459_));
 sg13g2_a21o_1 _16056_ (.A2(_02474_),
    .A1(_02470_),
    .B1(_02460_),
    .X(_02476_));
 sg13g2_a221oi_1 _16057_ (.B2(net7363),
    .C1(net7361),
    .B1(_02476_),
    .A1(_02292_),
    .Y(_02477_),
    .A2(_02446_));
 sg13g2_mux4_1 _16058_ (.S0(net7915),
    .A0(_01078_),
    .A1(_01113_),
    .A2(_01149_),
    .A3(_01184_),
    .S1(net7828),
    .X(_02478_));
 sg13g2_inv_1 _16059_ (.Y(_02479_),
    .A(_02478_));
 sg13g2_mux4_1 _16060_ (.S0(net7915),
    .A0(_01219_),
    .A1(_01254_),
    .A2(_01289_),
    .A3(_01325_),
    .S1(net7828),
    .X(_02480_));
 sg13g2_nor2_1 _16061_ (.A(net7445),
    .B(_02480_),
    .Y(_02481_));
 sg13g2_mux2_1 _16062_ (.A0(_00674_),
    .A1(_00706_),
    .S(net7858),
    .X(_02482_));
 sg13g2_mux2_1 _16063_ (.A0(_00738_),
    .A1(_00770_),
    .S(net7858),
    .X(_02483_));
 sg13g2_mux2_1 _16064_ (.A0(_01368_),
    .A1(_00642_),
    .S(net7858),
    .X(_02484_));
 sg13g2_and2_1 _16065_ (.A(net7858),
    .B(_01016_),
    .X(_02485_));
 sg13g2_mux4_1 _16066_ (.S0(net7829),
    .A0(_02482_),
    .A1(_02483_),
    .A2(_02485_),
    .A3(_02484_),
    .S1(net7484),
    .X(_02486_));
 sg13g2_nand2b_1 _16067_ (.Y(_02487_),
    .B(_08973_),
    .A_N(_02486_));
 sg13g2_mux4_1 _16068_ (.S0(net7916),
    .A0(_00937_),
    .A1(_00973_),
    .A2(_01008_),
    .A3(_01043_),
    .S1(net7828),
    .X(_02488_));
 sg13g2_nand2_1 _16069_ (.Y(_02489_),
    .A(net7814),
    .B(_02488_));
 sg13g2_mux4_1 _16070_ (.S0(net7913),
    .A0(_00802_),
    .A1(_00834_),
    .A2(_00867_),
    .A3(_00902_),
    .S1(net7828),
    .X(_02490_));
 sg13g2_a21oi_1 _16071_ (.A1(net7484),
    .A2(_02490_),
    .Y(_02491_),
    .B1(net7540));
 sg13g2_mux2_1 _16072_ (.A0(_01430_),
    .A1(_01465_),
    .S(net7916),
    .X(_02492_));
 sg13g2_nor3_1 _16073_ (.A(_09152_),
    .B(net7460),
    .C(_02492_),
    .Y(_02493_));
 sg13g2_mux2_1 _16074_ (.A0(_01360_),
    .A1(_01395_),
    .S(net7916),
    .X(_02494_));
 sg13g2_nor3_1 _16075_ (.A(_09152_),
    .B(net7470),
    .C(_02494_),
    .Y(_02495_));
 sg13g2_mux2_1 _16076_ (.A0(_01501_),
    .A1(_01536_),
    .S(net7916),
    .X(_02496_));
 sg13g2_nor3_1 _16077_ (.A(_09028_),
    .B(_09152_),
    .C(_02496_),
    .Y(_02497_));
 sg13g2_mux2_1 _16078_ (.A0(_01571_),
    .A1(_00614_),
    .S(net7916),
    .X(_02498_));
 sg13g2_nor2_1 _16079_ (.A(net7449),
    .B(_02498_),
    .Y(_02499_));
 sg13g2_nor4_1 _16080_ (.A(_02493_),
    .B(_02495_),
    .C(_02497_),
    .D(_02499_),
    .Y(_02500_));
 sg13g2_a221oi_1 _16081_ (.B2(_02491_),
    .C1(_02481_),
    .B1(_02489_),
    .A1(_12135_),
    .Y(_02501_),
    .A2(_02479_));
 sg13g2_and3_1 _16082_ (.X(_02502_),
    .A(_02487_),
    .B(_02500_),
    .C(_02501_));
 sg13g2_nand3_1 _16083_ (.B(_02500_),
    .C(_02501_),
    .A(_02487_),
    .Y(_02503_));
 sg13g2_nand2b_1 _16084_ (.Y(_02504_),
    .B(net8001),
    .A_N(_01647_));
 sg13g2_o21ai_1 _16085_ (.B1(_02504_),
    .Y(_02505_),
    .A1(_01612_),
    .A2(net7480));
 sg13g2_a221oi_1 _16086_ (.B2(net8005),
    .C1(_02505_),
    .B1(net7347),
    .A1(net7352),
    .Y(_02506_),
    .A2(_02476_));
 sg13g2_nor2_1 _16087_ (.A(net7375),
    .B(_02506_),
    .Y(_02507_));
 sg13g2_a21oi_1 _16088_ (.A1(net6919),
    .A2(_02477_),
    .Y(_02508_),
    .B1(_02507_));
 sg13g2_o21ai_1 _16089_ (.B1(_02508_),
    .Y(_02509_),
    .A1(net6980),
    .A2(_02477_));
 sg13g2_nand2_1 _16090_ (.Y(_02510_),
    .A(net7843),
    .B(_02293_));
 sg13g2_mux2_1 _16091_ (.A0(_01431_),
    .A1(_01466_),
    .S(net7789),
    .X(_02511_));
 sg13g2_nor3_1 _16092_ (.A(net7576),
    .B(net7570),
    .C(_02511_),
    .Y(_02512_));
 sg13g2_mux2_1 _16093_ (.A0(_01361_),
    .A1(_01396_),
    .S(net7789),
    .X(_02513_));
 sg13g2_nor3_1 _16094_ (.A(net7576),
    .B(net7557),
    .C(_02513_),
    .Y(_02514_));
 sg13g2_mux2_1 _16095_ (.A0(_01502_),
    .A1(_01537_),
    .S(net7789),
    .X(_02515_));
 sg13g2_nor3_1 _16096_ (.A(net7576),
    .B(net7566),
    .C(_02515_),
    .Y(_02516_));
 sg13g2_mux2_1 _16097_ (.A0(_01572_),
    .A1(_00615_),
    .S(net7789),
    .X(_02517_));
 sg13g2_nor2_1 _16098_ (.A(net7554),
    .B(_02517_),
    .Y(_02518_));
 sg13g2_nor4_1 _16099_ (.A(_02512_),
    .B(_02514_),
    .C(_02516_),
    .D(_02518_),
    .Y(_02519_));
 sg13g2_mux4_1 _16100_ (.S0(net7789),
    .A0(_01220_),
    .A1(_01255_),
    .A2(_01290_),
    .A3(_01326_),
    .S1(net7737),
    .X(_02520_));
 sg13g2_or2_1 _16101_ (.X(_02521_),
    .B(_02520_),
    .A(net7587));
 sg13g2_mux4_1 _16102_ (.S0(net7789),
    .A0(_01079_),
    .A1(_01114_),
    .A2(_01150_),
    .A3(_01185_),
    .S1(net7737),
    .X(_02522_));
 sg13g2_nand2b_1 _16103_ (.Y(_02523_),
    .B(net7434),
    .A_N(_02522_));
 sg13g2_mux4_1 _16104_ (.S0(net7788),
    .A0(_00803_),
    .A1(_00835_),
    .A2(_00868_),
    .A3(_00903_),
    .S1(net7743),
    .X(_02524_));
 sg13g2_mux4_1 _16105_ (.S0(net7788),
    .A0(_00938_),
    .A1(_00974_),
    .A2(_01009_),
    .A3(_01044_),
    .S1(net7743),
    .X(_02525_));
 sg13g2_a22oi_1 _16106_ (.Y(_02526_),
    .B1(_02525_),
    .B2(_02462_),
    .A2(_02524_),
    .A1(net7604));
 sg13g2_mux2_1 _16107_ (.A0(_00643_),
    .A1(_00771_),
    .S(net7717),
    .X(_02527_));
 sg13g2_a22oi_1 _16108_ (.Y(_02528_),
    .B1(_02527_),
    .B2(_08288_),
    .A2(_10463_),
    .A1(_01027_));
 sg13g2_a21oi_1 _16109_ (.A1(_01379_),
    .A2(_10449_),
    .Y(_02529_),
    .B1(net7688));
 sg13g2_mux2_1 _16110_ (.A0(_00675_),
    .A1(_00707_),
    .S(net7781),
    .X(_02530_));
 sg13g2_a22oi_1 _16111_ (.Y(_02531_),
    .B1(_02530_),
    .B2(net7517),
    .A2(net7596),
    .A1(_00739_));
 sg13g2_nand2b_1 _16112_ (.Y(_02532_),
    .B(_14476_),
    .A_N(_02531_));
 sg13g2_nand4_1 _16113_ (.B(_02528_),
    .C(_02529_),
    .A(_02526_),
    .Y(_02533_),
    .D(_02532_));
 sg13g2_nand4_1 _16114_ (.B(_02521_),
    .C(_02523_),
    .A(_02519_),
    .Y(_02534_),
    .D(_02533_));
 sg13g2_a221oi_1 _16115_ (.B2(net7363),
    .C1(net7361),
    .B1(_02534_),
    .A1(_02292_),
    .Y(_02535_),
    .A2(_02510_));
 sg13g2_mux4_1 _16116_ (.S0(net7845),
    .A0(_01220_),
    .A1(_01255_),
    .A2(_01290_),
    .A3(_01326_),
    .S1(net7822),
    .X(_02536_));
 sg13g2_mux4_1 _16117_ (.S0(net7845),
    .A0(_01079_),
    .A1(_01114_),
    .A2(_01150_),
    .A3(_01185_),
    .S1(net7822),
    .X(_02537_));
 sg13g2_mux4_1 _16118_ (.S0(net7845),
    .A0(_01361_),
    .A1(_01396_),
    .A2(_01431_),
    .A3(_01466_),
    .S1(net7822),
    .X(_02538_));
 sg13g2_mux4_1 _16119_ (.S0(net7845),
    .A0(_01502_),
    .A1(_01537_),
    .A2(_01572_),
    .A3(_00615_),
    .S1(net7822),
    .X(_02539_));
 sg13g2_mux4_1 _16120_ (.S0(net7483),
    .A0(_02536_),
    .A1(_02537_),
    .A2(_02539_),
    .A3(_02538_),
    .S1(net7807),
    .X(_02540_));
 sg13g2_nand2b_1 _16121_ (.Y(_02541_),
    .B(net7805),
    .A_N(_02540_));
 sg13g2_mux4_1 _16122_ (.S0(net7843),
    .A0(_00675_),
    .A1(_00707_),
    .A2(_00739_),
    .A3(_00771_),
    .S1(net7823),
    .X(_02542_));
 sg13g2_mux2_1 _16123_ (.A0(_01379_),
    .A1(_00643_),
    .S(net7843),
    .X(_02543_));
 sg13g2_and2_1 _16124_ (.A(net7843),
    .B(_01027_),
    .X(_02544_));
 sg13g2_mux2_1 _16125_ (.A0(_02544_),
    .A1(_02543_),
    .S(net7823),
    .X(_02545_));
 sg13g2_mux4_1 _16126_ (.S0(net7855),
    .A0(_00938_),
    .A1(_00974_),
    .A2(_01009_),
    .A3(_01044_),
    .S1(net7822),
    .X(_02546_));
 sg13g2_mux4_1 _16127_ (.S0(net7844),
    .A0(_00803_),
    .A1(_00835_),
    .A2(_00868_),
    .A3(_00903_),
    .S1(net7822),
    .X(_02547_));
 sg13g2_mux4_1 _16128_ (.S0(net7483),
    .A0(_02542_),
    .A1(_02545_),
    .A2(_02546_),
    .A3(_02547_),
    .S1(net7807),
    .X(_02548_));
 sg13g2_o21ai_1 _16129_ (.B1(_02541_),
    .Y(_02549_),
    .A1(net7805),
    .A2(_02548_));
 sg13g2_nand2_1 _16130_ (.Y(_02550_),
    .A(_02098_),
    .B(net7999));
 sg13g2_o21ai_1 _16131_ (.B1(_02550_),
    .Y(_02551_),
    .A1(_01613_),
    .A2(net7478));
 sg13g2_a221oi_1 _16132_ (.B2(net8004),
    .C1(_02551_),
    .B1(_02549_),
    .A1(net7352),
    .Y(_02552_),
    .A2(_02534_));
 sg13g2_nor2_1 _16133_ (.A(net7375),
    .B(_02552_),
    .Y(_02553_));
 sg13g2_a21oi_1 _16134_ (.A1(net6918),
    .A2(_02535_),
    .Y(_02554_),
    .B1(_02553_));
 sg13g2_o21ai_1 _16135_ (.B1(_02554_),
    .Y(_02555_),
    .A1(net6978),
    .A2(_02535_));
 sg13g2_nand2_1 _16136_ (.Y(_02556_),
    .A(net7823),
    .B(_02293_));
 sg13g2_mux2_1 _16137_ (.A0(_01432_),
    .A1(_01468_),
    .S(net7763),
    .X(_02557_));
 sg13g2_nor3_1 _16138_ (.A(net7582),
    .B(net7567),
    .C(_02557_),
    .Y(_02558_));
 sg13g2_mux2_1 _16139_ (.A0(_01362_),
    .A1(_01397_),
    .S(net7763),
    .X(_02559_));
 sg13g2_nor3_1 _16140_ (.A(net7582),
    .B(net7559),
    .C(_02559_),
    .Y(_02560_));
 sg13g2_mux2_1 _16141_ (.A0(_01503_),
    .A1(_01538_),
    .S(net7763),
    .X(_02561_));
 sg13g2_nor3_1 _16142_ (.A(net7582),
    .B(net7564),
    .C(_02561_),
    .Y(_02562_));
 sg13g2_mux2_1 _16143_ (.A0(_01573_),
    .A1(_00616_),
    .S(net7763),
    .X(_02563_));
 sg13g2_nor2_1 _16144_ (.A(net7551),
    .B(_02563_),
    .Y(_02564_));
 sg13g2_or4_1 _16145_ (.A(_02558_),
    .B(_02560_),
    .C(_02562_),
    .D(_02564_),
    .X(_02565_));
 sg13g2_mux4_1 _16146_ (.S0(net7751),
    .A0(_01221_),
    .A1(_01256_),
    .A2(_01292_),
    .A3(_01327_),
    .S1(net7720),
    .X(_02566_));
 sg13g2_mux4_1 _16147_ (.S0(net7751),
    .A0(_01080_),
    .A1(_01116_),
    .A2(_01151_),
    .A3(_01186_),
    .S1(net7720),
    .X(_02567_));
 sg13g2_nand2b_1 _16148_ (.Y(_02568_),
    .B(net7698),
    .A_N(_02566_));
 sg13g2_o21ai_1 _16149_ (.B1(_02568_),
    .Y(_02569_),
    .A1(net7698),
    .A2(_02567_));
 sg13g2_a21o_1 _16150_ (.A2(_02569_),
    .A1(net7590),
    .B1(_02565_),
    .X(_02570_));
 sg13g2_mux4_1 _16151_ (.S0(net7763),
    .A0(_00804_),
    .A1(_00836_),
    .A2(_00869_),
    .A3(_00904_),
    .S1(net7725),
    .X(_02571_));
 sg13g2_mux4_1 _16152_ (.S0(net7763),
    .A0(_00940_),
    .A1(_00975_),
    .A2(_01010_),
    .A3(_01045_),
    .S1(net7725),
    .X(_02572_));
 sg13g2_and2_1 _16153_ (.A(net7640),
    .B(_02572_),
    .X(_02573_));
 sg13g2_and3_1 _16154_ (.X(_02574_),
    .A(_01038_),
    .B(net7599),
    .C(net7597));
 sg13g2_nand2_1 _16155_ (.Y(_02575_),
    .A(net7705),
    .B(_00772_));
 sg13g2_nand2b_1 _16156_ (.Y(_02576_),
    .B(_00644_),
    .A_N(net7705));
 sg13g2_a21oi_1 _16157_ (.A1(_02575_),
    .A2(_02576_),
    .Y(_02577_),
    .B1(net7601));
 sg13g2_and3_1 _16158_ (.X(_02578_),
    .A(_01390_),
    .B(net7599),
    .C(net7594));
 sg13g2_nor4_1 _16159_ (.A(net7687),
    .B(_02574_),
    .C(_02577_),
    .D(_02578_),
    .Y(_02579_));
 sg13g2_mux2_1 _16160_ (.A0(_00676_),
    .A1(_00708_),
    .S(net7765),
    .X(_02580_));
 sg13g2_nor2b_1 _16161_ (.A(net7773),
    .B_N(_00740_),
    .Y(_02581_));
 sg13g2_mux2_1 _16162_ (.A0(_02580_),
    .A1(_02581_),
    .S(net7722),
    .X(_02582_));
 sg13g2_a221oi_1 _16163_ (.B2(net7442),
    .C1(_02573_),
    .B1(_02582_),
    .A1(net7605),
    .Y(_02583_),
    .A2(_02571_));
 sg13g2_a221oi_1 _16164_ (.B2(_02583_),
    .C1(_02565_),
    .B1(_02579_),
    .A1(net7590),
    .Y(_02584_),
    .A2(_02569_));
 sg13g2_a21o_1 _16165_ (.A2(_02583_),
    .A1(_02579_),
    .B1(_02570_),
    .X(_02585_));
 sg13g2_a221oi_1 _16166_ (.B2(net7363),
    .C1(net7361),
    .B1(_02585_),
    .A1(_02292_),
    .Y(_02586_),
    .A2(_02556_));
 sg13g2_mux2_1 _16167_ (.A0(_00804_),
    .A1(_00836_),
    .S(net7914),
    .X(_02587_));
 sg13g2_nor2_1 _16168_ (.A(net7467),
    .B(_02587_),
    .Y(_02588_));
 sg13g2_mux2_1 _16169_ (.A0(_00869_),
    .A1(_00904_),
    .S(net7914),
    .X(_02589_));
 sg13g2_nor2_1 _16170_ (.A(net7457),
    .B(_02589_),
    .Y(_02590_));
 sg13g2_mux2_1 _16171_ (.A0(_01010_),
    .A1(_01045_),
    .S(net7913),
    .X(_02591_));
 sg13g2_nor2_1 _16172_ (.A(net7524),
    .B(_02591_),
    .Y(_02592_));
 sg13g2_mux2_1 _16173_ (.A0(_00940_),
    .A1(_00975_),
    .S(net7913),
    .X(_02593_));
 sg13g2_o21ai_1 _16174_ (.B1(net7542),
    .Y(_02594_),
    .A1(_09028_),
    .A2(_02593_));
 sg13g2_nor4_1 _16175_ (.A(_02588_),
    .B(_02590_),
    .C(_02592_),
    .D(_02594_),
    .Y(_02595_));
 sg13g2_mux2_1 _16176_ (.A0(_01080_),
    .A1(_01116_),
    .S(net7898),
    .X(_02596_));
 sg13g2_nor2_1 _16177_ (.A(net7468),
    .B(_02596_),
    .Y(_02597_));
 sg13g2_mux2_1 _16178_ (.A0(_01151_),
    .A1(_01186_),
    .S(net7898),
    .X(_02598_));
 sg13g2_nor2_1 _16179_ (.A(net7459),
    .B(_02598_),
    .Y(_02599_));
 sg13g2_mux2_1 _16180_ (.A0(_01292_),
    .A1(_01327_),
    .S(net7898),
    .X(_02600_));
 sg13g2_nor2_1 _16181_ (.A(net7523),
    .B(_02600_),
    .Y(_02601_));
 sg13g2_mux2_1 _16182_ (.A0(_01221_),
    .A1(_01256_),
    .S(net7898),
    .X(_02602_));
 sg13g2_o21ai_1 _16183_ (.B1(net7503),
    .Y(_02603_),
    .A1(net7508),
    .A2(_02602_));
 sg13g2_nor4_1 _16184_ (.A(_02597_),
    .B(_02599_),
    .C(_02601_),
    .D(_02603_),
    .Y(_02604_));
 sg13g2_mux4_1 _16185_ (.S0(net7913),
    .A0(_01503_),
    .A1(_01538_),
    .A2(_01573_),
    .A3(_00616_),
    .S1(net7828),
    .X(_02605_));
 sg13g2_nand2_1 _16186_ (.Y(_02606_),
    .A(net7810),
    .B(_02605_));
 sg13g2_mux4_1 _16187_ (.S0(net7913),
    .A0(_01362_),
    .A1(_01397_),
    .A2(_01432_),
    .A3(_01468_),
    .S1(net7828),
    .X(_02607_));
 sg13g2_nand2_1 _16188_ (.Y(_02608_),
    .A(net7485),
    .B(_02607_));
 sg13g2_a21oi_1 _16189_ (.A1(_02606_),
    .A2(_02608_),
    .Y(_02609_),
    .B1(net7487));
 sg13g2_mux4_1 _16190_ (.S0(net7860),
    .A0(_00676_),
    .A1(_00708_),
    .A2(_00740_),
    .A3(_00772_),
    .S1(net7829),
    .X(_02610_));
 sg13g2_mux2_1 _16191_ (.A0(_01390_),
    .A1(_00644_),
    .S(net7860),
    .X(_02611_));
 sg13g2_a22oi_1 _16192_ (.Y(_02612_),
    .B1(_02611_),
    .B2(net7829),
    .A2(_08988_),
    .A1(_01038_));
 sg13g2_o21ai_1 _16193_ (.B1(_08973_),
    .Y(_02613_),
    .A1(net7485),
    .A2(_02610_));
 sg13g2_a21oi_1 _16194_ (.A1(net7485),
    .A2(_02612_),
    .Y(_02614_),
    .B1(_02613_));
 sg13g2_nor4_1 _16195_ (.A(_02595_),
    .B(net7418),
    .C(_02609_),
    .D(_02614_),
    .Y(_02615_));
 sg13g2_or4_1 _16196_ (.A(_02595_),
    .B(net7418),
    .C(_02609_),
    .D(_02614_),
    .X(_02616_));
 sg13g2_nand2b_1 _16197_ (.Y(_02617_),
    .B(net7999),
    .A_N(_01650_));
 sg13g2_o21ai_1 _16198_ (.B1(_02617_),
    .Y(_02618_),
    .A1(_01614_),
    .A2(net7480));
 sg13g2_a21oi_1 _16199_ (.A1(net8007),
    .A2(_02615_),
    .Y(_02619_),
    .B1(_02618_));
 sg13g2_o21ai_1 _16200_ (.B1(_02619_),
    .Y(_02620_),
    .A1(_09277_),
    .A2(_02584_));
 sg13g2_a22oi_1 _16201_ (.Y(_02621_),
    .B1(_02620_),
    .B2(net7377),
    .A2(_02586_),
    .A1(net6919));
 sg13g2_o21ai_1 _16202_ (.B1(_02621_),
    .Y(_02622_),
    .A1(net6980),
    .A2(_02586_));
 sg13g2_nand2_1 _16203_ (.Y(_02623_),
    .A(net7812),
    .B(_02293_));
 sg13g2_mux2_1 _16204_ (.A0(_01504_),
    .A1(_01539_),
    .S(net7756),
    .X(_02624_));
 sg13g2_nor3_1 _16205_ (.A(net7583),
    .B(net7565),
    .C(_02624_),
    .Y(_02625_));
 sg13g2_mux2_1 _16206_ (.A0(_01574_),
    .A1(_00617_),
    .S(net7756),
    .X(_02626_));
 sg13g2_nor2_1 _16207_ (.A(net7552),
    .B(_02626_),
    .Y(_02627_));
 sg13g2_mux2_1 _16208_ (.A0(_01363_),
    .A1(_01398_),
    .S(net7757),
    .X(_02628_));
 sg13g2_nor3_1 _16209_ (.A(net7583),
    .B(net7560),
    .C(_02628_),
    .Y(_02629_));
 sg13g2_mux2_1 _16210_ (.A0(_01433_),
    .A1(_01469_),
    .S(net7757),
    .X(_02630_));
 sg13g2_nor3_1 _16211_ (.A(net7583),
    .B(net7568),
    .C(_02630_),
    .Y(_02631_));
 sg13g2_or4_1 _16212_ (.A(_02625_),
    .B(_02627_),
    .C(_02629_),
    .D(_02631_),
    .X(_02632_));
 sg13g2_mux4_1 _16213_ (.S0(net7750),
    .A0(_01081_),
    .A1(_01117_),
    .A2(_01152_),
    .A3(_01187_),
    .S1(net7718),
    .X(_02633_));
 sg13g2_mux4_1 _16214_ (.S0(net7750),
    .A0(_01222_),
    .A1(_01257_),
    .A2(_01293_),
    .A3(_01328_),
    .S1(net7718),
    .X(_02634_));
 sg13g2_nand2b_1 _16215_ (.Y(_02635_),
    .B(net7698),
    .A_N(_02634_));
 sg13g2_o21ai_1 _16216_ (.B1(_02635_),
    .Y(_02636_),
    .A1(net7698),
    .A2(_02633_));
 sg13g2_a21o_1 _16217_ (.A2(_02636_),
    .A1(net7589),
    .B1(_02632_),
    .X(_02637_));
 sg13g2_mux4_1 _16218_ (.S0(net7749),
    .A0(_00805_),
    .A1(_00837_),
    .A2(_00870_),
    .A3(_00905_),
    .S1(net7719),
    .X(_02638_));
 sg13g2_mux4_1 _16219_ (.S0(net7749),
    .A0(_00941_),
    .A1(_00976_),
    .A2(_01011_),
    .A3(_01046_),
    .S1(net7719),
    .X(_02639_));
 sg13g2_and2_1 _16220_ (.A(net7640),
    .B(_02639_),
    .X(_02640_));
 sg13g2_and3_1 _16221_ (.X(_02641_),
    .A(_01049_),
    .B(net7599),
    .C(net7597));
 sg13g2_nand2_1 _16222_ (.Y(_02642_),
    .A(net7700),
    .B(_00773_));
 sg13g2_nand2b_1 _16223_ (.Y(_02643_),
    .B(_00645_),
    .A_N(net7701));
 sg13g2_a21oi_1 _16224_ (.A1(_02642_),
    .A2(_02643_),
    .Y(_02644_),
    .B1(net7601));
 sg13g2_and3_1 _16225_ (.X(_02645_),
    .A(_01401_),
    .B(net7599),
    .C(net7593));
 sg13g2_nor4_1 _16226_ (.A(net7689),
    .B(_02641_),
    .C(_02644_),
    .D(_02645_),
    .Y(_02646_));
 sg13g2_mux2_1 _16227_ (.A0(_00677_),
    .A1(_00709_),
    .S(net7760),
    .X(_02647_));
 sg13g2_nor2b_1 _16228_ (.A(net7760),
    .B_N(_00741_),
    .Y(_02648_));
 sg13g2_mux2_1 _16229_ (.A0(_02647_),
    .A1(_02648_),
    .S(net7735),
    .X(_02649_));
 sg13g2_a221oi_1 _16230_ (.B2(net7442),
    .C1(_02640_),
    .B1(_02649_),
    .A1(net7606),
    .Y(_02650_),
    .A2(_02638_));
 sg13g2_a221oi_1 _16231_ (.B2(_02650_),
    .C1(_02632_),
    .B1(_02646_),
    .A1(net7589),
    .Y(_02651_),
    .A2(_02636_));
 sg13g2_a21o_1 _16232_ (.A2(_02650_),
    .A1(_02646_),
    .B1(_02637_),
    .X(_02652_));
 sg13g2_a221oi_1 _16233_ (.B2(net7363),
    .C1(net7361),
    .B1(_02652_),
    .A1(_02292_),
    .Y(_02653_),
    .A2(_02623_));
 sg13g2_mux2_1 _16234_ (.A0(_00870_),
    .A1(_00905_),
    .S(net7907),
    .X(_02654_));
 sg13g2_nor2_1 _16235_ (.A(net7458),
    .B(_02654_),
    .Y(_02655_));
 sg13g2_mux2_1 _16236_ (.A0(_00805_),
    .A1(_00837_),
    .S(net7907),
    .X(_02656_));
 sg13g2_nor2_1 _16237_ (.A(net7469),
    .B(_02656_),
    .Y(_02657_));
 sg13g2_mux2_1 _16238_ (.A0(_01011_),
    .A1(_01046_),
    .S(net7906),
    .X(_02658_));
 sg13g2_nor2_1 _16239_ (.A(net7522),
    .B(_02658_),
    .Y(_02659_));
 sg13g2_mux2_1 _16240_ (.A0(_00941_),
    .A1(_00976_),
    .S(net7901),
    .X(_02660_));
 sg13g2_o21ai_1 _16241_ (.B1(net7541),
    .Y(_02661_),
    .A1(net7507),
    .A2(_02660_));
 sg13g2_nor4_1 _16242_ (.A(_02655_),
    .B(_02657_),
    .C(_02659_),
    .D(_02661_),
    .Y(_02662_));
 sg13g2_mux2_1 _16243_ (.A0(_01081_),
    .A1(_01117_),
    .S(net7897),
    .X(_02663_));
 sg13g2_nor2_1 _16244_ (.A(net7468),
    .B(_02663_),
    .Y(_02664_));
 sg13g2_mux2_1 _16245_ (.A0(_01152_),
    .A1(_01187_),
    .S(net7897),
    .X(_02665_));
 sg13g2_nor2_1 _16246_ (.A(net7459),
    .B(_02665_),
    .Y(_02666_));
 sg13g2_mux2_1 _16247_ (.A0(_01293_),
    .A1(_01328_),
    .S(net7896),
    .X(_02667_));
 sg13g2_nor2_1 _16248_ (.A(net7523),
    .B(_02667_),
    .Y(_02668_));
 sg13g2_mux2_1 _16249_ (.A0(_01222_),
    .A1(_01257_),
    .S(net7896),
    .X(_02669_));
 sg13g2_o21ai_1 _16250_ (.B1(net7503),
    .Y(_02670_),
    .A1(net7507),
    .A2(_02669_));
 sg13g2_nor4_1 _16251_ (.A(_02664_),
    .B(_02666_),
    .C(_02668_),
    .D(_02670_),
    .Y(_02671_));
 sg13g2_mux4_1 _16252_ (.S0(net7838),
    .A0(_00677_),
    .A1(_00709_),
    .A2(_00741_),
    .A3(_00773_),
    .S1(net7823),
    .X(_02672_));
 sg13g2_mux2_1 _16253_ (.A0(_01401_),
    .A1(_00645_),
    .S(net7836),
    .X(_02673_));
 sg13g2_a22oi_1 _16254_ (.Y(_02674_),
    .B1(_02673_),
    .B2(net7829),
    .A2(_08988_),
    .A1(_01049_));
 sg13g2_o21ai_1 _16255_ (.B1(_08973_),
    .Y(_02675_),
    .A1(net7486),
    .A2(_02672_));
 sg13g2_a21oi_1 _16256_ (.A1(net7486),
    .A2(_02674_),
    .Y(_02676_),
    .B1(_02675_));
 sg13g2_mux4_1 _16257_ (.S0(net7905),
    .A0(_01504_),
    .A1(_01539_),
    .A2(_01574_),
    .A3(_00617_),
    .S1(net7817),
    .X(_02677_));
 sg13g2_mux4_1 _16258_ (.S0(net7905),
    .A0(_01363_),
    .A1(_01398_),
    .A2(_01433_),
    .A3(_01469_),
    .S1(net7817),
    .X(_02678_));
 sg13g2_nand2_1 _16259_ (.Y(_02679_),
    .A(net7809),
    .B(_02677_));
 sg13g2_nand2_1 _16260_ (.Y(_02680_),
    .A(net7486),
    .B(_02678_));
 sg13g2_a21oi_1 _16261_ (.A1(_02679_),
    .A2(_02680_),
    .Y(_02681_),
    .B1(net7488));
 sg13g2_nor4_1 _16262_ (.A(_02662_),
    .B(_02671_),
    .C(_02676_),
    .D(_02681_),
    .Y(_02682_));
 sg13g2_nor2_1 _16263_ (.A(_01615_),
    .B(net7480),
    .Y(_02683_));
 sg13g2_a221oi_1 _16264_ (.B2(net7344),
    .C1(_02683_),
    .B1(net8005),
    .A1(_02089_),
    .Y(_02684_),
    .A2(net8001));
 sg13g2_o21ai_1 _16265_ (.B1(_02684_),
    .Y(_02685_),
    .A1(_09277_),
    .A2(net7345));
 sg13g2_a22oi_1 _16266_ (.Y(_02686_),
    .B1(_02685_),
    .B2(net7377),
    .A2(_02653_),
    .A1(net6919));
 sg13g2_o21ai_1 _16267_ (.B1(_02686_),
    .Y(_02687_),
    .A1(net6979),
    .A2(_02653_));
 sg13g2_nand2_1 _16268_ (.Y(_02688_),
    .A(net7807),
    .B(_02293_));
 sg13g2_mux2_1 _16269_ (.A0(_01575_),
    .A1(_00619_),
    .S(net7755),
    .X(_02689_));
 sg13g2_nor2_1 _16270_ (.A(net7553),
    .B(_02689_),
    .Y(_02690_));
 sg13g2_mux2_1 _16271_ (.A0(_01505_),
    .A1(_01540_),
    .S(net7756),
    .X(_02691_));
 sg13g2_nor3_1 _16272_ (.A(net7581),
    .B(net7564),
    .C(_02691_),
    .Y(_02692_));
 sg13g2_mux2_1 _16273_ (.A0(_01435_),
    .A1(_01470_),
    .S(net7755),
    .X(_02693_));
 sg13g2_nor3_1 _16274_ (.A(net7581),
    .B(net7568),
    .C(_02693_),
    .Y(_02694_));
 sg13g2_mux2_1 _16275_ (.A0(_01364_),
    .A1(_01399_),
    .S(net7756),
    .X(_02695_));
 sg13g2_nor3_1 _16276_ (.A(net7581),
    .B(net7560),
    .C(_02695_),
    .Y(_02696_));
 sg13g2_nor4_1 _16277_ (.A(_02690_),
    .B(_02692_),
    .C(_02694_),
    .D(_02696_),
    .Y(_02697_));
 sg13g2_mux4_1 _16278_ (.S0(net7750),
    .A0(_01083_),
    .A1(_01118_),
    .A2(_01153_),
    .A3(_01188_),
    .S1(net7718),
    .X(_02698_));
 sg13g2_inv_1 _16279_ (.Y(_02699_),
    .A(_02698_));
 sg13g2_mux4_1 _16280_ (.S0(net7751),
    .A0(_01223_),
    .A1(_01259_),
    .A2(_01294_),
    .A3(_01329_),
    .S1(net7720),
    .X(_02700_));
 sg13g2_nor2_1 _16281_ (.A(net7586),
    .B(_02700_),
    .Y(_02701_));
 sg13g2_a21oi_1 _16282_ (.A1(net7433),
    .A2(_02699_),
    .Y(_02702_),
    .B1(_02701_));
 sg13g2_a21oi_1 _16283_ (.A1(_01412_),
    .A2(net7424),
    .Y(_02703_),
    .B1(net7688));
 sg13g2_mux2_1 _16284_ (.A0(_00646_),
    .A1(_00774_),
    .S(net7701),
    .X(_02704_));
 sg13g2_a22oi_1 _16285_ (.Y(_02705_),
    .B1(_02704_),
    .B2(_08288_),
    .A2(net7422),
    .A1(_01060_));
 sg13g2_mux2_1 _16286_ (.A0(_00678_),
    .A1(_00710_),
    .S(net7753),
    .X(_02706_));
 sg13g2_a22oi_1 _16287_ (.Y(_02707_),
    .B1(_02706_),
    .B2(net7519),
    .A2(net7593),
    .A1(_00742_));
 sg13g2_nand2b_1 _16288_ (.Y(_02708_),
    .B(net7442),
    .A_N(_02707_));
 sg13g2_mux4_1 _16289_ (.S0(net7762),
    .A0(_00806_),
    .A1(_00838_),
    .A2(_00871_),
    .A3(_00907_),
    .S1(net7730),
    .X(_02709_));
 sg13g2_mux4_1 _16290_ (.S0(net7762),
    .A0(_00942_),
    .A1(_00977_),
    .A2(_01012_),
    .A3(_01047_),
    .S1(net7730),
    .X(_02710_));
 sg13g2_a22oi_1 _16291_ (.Y(_02711_),
    .B1(_02710_),
    .B2(net7640),
    .A2(_02709_),
    .A1(net7606));
 sg13g2_nand4_1 _16292_ (.B(_02705_),
    .C(_02708_),
    .A(_02703_),
    .Y(_02712_),
    .D(_02711_));
 sg13g2_inv_1 _16293_ (.Y(_02713_),
    .A(net7263));
 sg13g2_nand3_1 _16294_ (.B(_02702_),
    .C(_02712_),
    .A(_02697_),
    .Y(_02714_));
 sg13g2_a221oi_1 _16295_ (.B2(net7363),
    .C1(net7361),
    .B1(_02714_),
    .A1(_02292_),
    .Y(_02715_),
    .A2(_02688_));
 sg13g2_mux2_1 _16296_ (.A0(_01575_),
    .A1(_00619_),
    .S(net7903),
    .X(_02716_));
 sg13g2_nor2_1 _16297_ (.A(net7448),
    .B(_02716_),
    .Y(_02717_));
 sg13g2_mux2_1 _16298_ (.A0(_01505_),
    .A1(_01540_),
    .S(net7904),
    .X(_02718_));
 sg13g2_nor3_1 _16299_ (.A(net7508),
    .B(net7487),
    .C(_02718_),
    .Y(_02719_));
 sg13g2_mux2_1 _16300_ (.A0(_01012_),
    .A1(_01047_),
    .S(net7911),
    .X(_02720_));
 sg13g2_nor3_1 _16301_ (.A(net7539),
    .B(net7522),
    .C(_02720_),
    .Y(_02721_));
 sg13g2_mux2_1 _16302_ (.A0(_00942_),
    .A1(_00977_),
    .S(net7907),
    .X(_02722_));
 sg13g2_nor3_1 _16303_ (.A(net7537),
    .B(net7505),
    .C(_02722_),
    .Y(_02723_));
 sg13g2_nor4_1 _16304_ (.A(_02717_),
    .B(_02719_),
    .C(_02721_),
    .D(_02723_),
    .Y(_02724_));
 sg13g2_mux2_1 _16305_ (.A0(_00806_),
    .A1(_00838_),
    .S(net7911),
    .X(_02725_));
 sg13g2_nor3_1 _16306_ (.A(net7539),
    .B(net7467),
    .C(_02725_),
    .Y(_02726_));
 sg13g2_mux2_1 _16307_ (.A0(_00871_),
    .A1(_00907_),
    .S(net7911),
    .X(_02727_));
 sg13g2_nor3_1 _16308_ (.A(net7539),
    .B(net7458),
    .C(_02727_),
    .Y(_02728_));
 sg13g2_mux2_1 _16309_ (.A0(_01364_),
    .A1(_01399_),
    .S(net7904),
    .X(_02729_));
 sg13g2_nor3_1 _16310_ (.A(net7487),
    .B(net7467),
    .C(_02729_),
    .Y(_02730_));
 sg13g2_mux2_1 _16311_ (.A0(_01435_),
    .A1(_01470_),
    .S(net7903),
    .X(_02731_));
 sg13g2_nor3_1 _16312_ (.A(net7487),
    .B(net7457),
    .C(_02731_),
    .Y(_02732_));
 sg13g2_nor4_1 _16313_ (.A(_02726_),
    .B(_02728_),
    .C(_02730_),
    .D(_02732_),
    .Y(_02733_));
 sg13g2_mux2_1 _16314_ (.A0(_01412_),
    .A1(_00646_),
    .S(net7836),
    .X(_02734_));
 sg13g2_and2_1 _16315_ (.A(net7836),
    .B(_01060_),
    .X(_02735_));
 sg13g2_mux2_1 _16316_ (.A0(_00678_),
    .A1(_00710_),
    .S(net7836),
    .X(_02736_));
 sg13g2_mux2_1 _16317_ (.A0(_00742_),
    .A1(_00774_),
    .S(net7836),
    .X(_02737_));
 sg13g2_mux4_1 _16318_ (.S0(net7810),
    .A0(_02735_),
    .A1(_02736_),
    .A2(_02734_),
    .A3(_02737_),
    .S1(net7820),
    .X(_02738_));
 sg13g2_or2_1 _16319_ (.X(_02739_),
    .B(_02738_),
    .A(net7528));
 sg13g2_mux4_1 _16320_ (.S0(net7896),
    .A0(_01223_),
    .A1(_01259_),
    .A2(_01294_),
    .A3(_01329_),
    .S1(net7818),
    .X(_02740_));
 sg13g2_nor2_1 _16321_ (.A(net7444),
    .B(_02740_),
    .Y(_02741_));
 sg13g2_mux4_1 _16322_ (.S0(net7897),
    .A0(_01083_),
    .A1(_01118_),
    .A2(_01153_),
    .A3(_01188_),
    .S1(net7818),
    .X(_02742_));
 sg13g2_nor3_1 _16323_ (.A(net7809),
    .B(net7499),
    .C(_02742_),
    .Y(_02743_));
 sg13g2_nor2_1 _16324_ (.A(_02741_),
    .B(_02743_),
    .Y(_02744_));
 sg13g2_and4_1 _16325_ (.A(_02724_),
    .B(_02733_),
    .C(_02739_),
    .D(_02744_),
    .X(_02745_));
 sg13g2_nand4_1 _16326_ (.B(_02733_),
    .C(_02739_),
    .A(_02724_),
    .Y(_02746_),
    .D(_02744_));
 sg13g2_nand2b_1 _16327_ (.Y(_02747_),
    .B(net7998),
    .A_N(_01652_));
 sg13g2_o21ai_1 _16328_ (.B1(_02747_),
    .Y(_02748_),
    .A1(_01616_),
    .A2(net7479));
 sg13g2_a221oi_1 _16329_ (.B2(net8006),
    .C1(_02748_),
    .B1(net7343),
    .A1(net7354),
    .Y(_02749_),
    .A2(net7263));
 sg13g2_nor2_1 _16330_ (.A(net7376),
    .B(_02749_),
    .Y(_02750_));
 sg13g2_a21oi_1 _16331_ (.A1(_08251_),
    .A2(_02715_),
    .Y(_02751_),
    .B1(_02750_));
 sg13g2_o21ai_1 _16332_ (.B1(_02751_),
    .Y(_02752_),
    .A1(net6980),
    .A2(_02715_));
 sg13g2_nand2_1 _16333_ (.Y(_02753_),
    .A(net7805),
    .B(_02293_));
 sg13g2_mux2_1 _16334_ (.A0(_01576_),
    .A1(_00620_),
    .S(net7758),
    .X(_02754_));
 sg13g2_nor2_1 _16335_ (.A(net7551),
    .B(_02754_),
    .Y(_02755_));
 sg13g2_mux2_1 _16336_ (.A0(_01506_),
    .A1(_01541_),
    .S(net7758),
    .X(_02756_));
 sg13g2_nor3_1 _16337_ (.A(net7582),
    .B(net7564),
    .C(_02756_),
    .Y(_02757_));
 sg13g2_mux2_1 _16338_ (.A0(_01436_),
    .A1(_01471_),
    .S(net7758),
    .X(_02758_));
 sg13g2_nor3_1 _16339_ (.A(net7580),
    .B(net7567),
    .C(_02758_),
    .Y(_02759_));
 sg13g2_mux2_1 _16340_ (.A0(_01365_),
    .A1(_01400_),
    .S(net7758),
    .X(_02760_));
 sg13g2_nor3_1 _16341_ (.A(net7580),
    .B(net7559),
    .C(_02760_),
    .Y(_02761_));
 sg13g2_nor4_1 _16342_ (.A(_02755_),
    .B(_02757_),
    .C(_02759_),
    .D(_02761_),
    .Y(_02762_));
 sg13g2_mux4_1 _16343_ (.S0(net7751),
    .A0(_01084_),
    .A1(_01119_),
    .A2(_01154_),
    .A3(_01189_),
    .S1(net7720),
    .X(_02763_));
 sg13g2_inv_1 _16344_ (.Y(_02764_),
    .A(_02763_));
 sg13g2_mux4_1 _16345_ (.S0(net7751),
    .A0(_01224_),
    .A1(_01260_),
    .A2(_01295_),
    .A3(_01330_),
    .S1(net7720),
    .X(_02765_));
 sg13g2_nor2_1 _16346_ (.A(net7586),
    .B(_02765_),
    .Y(_02766_));
 sg13g2_a21oi_1 _16347_ (.A1(net7434),
    .A2(_02764_),
    .Y(_02767_),
    .B1(_02766_));
 sg13g2_a21oi_1 _16348_ (.A1(_01423_),
    .A2(net7424),
    .Y(_02768_),
    .B1(net7687));
 sg13g2_mux2_1 _16349_ (.A0(_00647_),
    .A1(_00775_),
    .S(net7705),
    .X(_02769_));
 sg13g2_a22oi_1 _16350_ (.Y(_02770_),
    .B1(_02769_),
    .B2(_08288_),
    .A2(_10463_),
    .A1(_01071_));
 sg13g2_mux2_1 _16351_ (.A0(_00679_),
    .A1(_00711_),
    .S(net7764),
    .X(_02771_));
 sg13g2_a22oi_1 _16352_ (.Y(_02772_),
    .B1(_02771_),
    .B2(net7519),
    .A2(net7593),
    .A1(_00743_));
 sg13g2_nand2b_1 _16353_ (.Y(_02773_),
    .B(net7442),
    .A_N(_02772_));
 sg13g2_mux4_1 _16354_ (.S0(net7763),
    .A0(_00807_),
    .A1(_00839_),
    .A2(_00872_),
    .A3(_00908_),
    .S1(net7722),
    .X(_02774_));
 sg13g2_mux4_1 _16355_ (.S0(net7763),
    .A0(_00943_),
    .A1(_00978_),
    .A2(_01013_),
    .A3(_01048_),
    .S1(net7725),
    .X(_02775_));
 sg13g2_a22oi_1 _16356_ (.Y(_02776_),
    .B1(_02775_),
    .B2(net7640),
    .A2(_02774_),
    .A1(net7605));
 sg13g2_nand4_1 _16357_ (.B(_02770_),
    .C(_02773_),
    .A(_02768_),
    .Y(_02777_),
    .D(_02776_));
 sg13g2_inv_1 _16358_ (.Y(_02778_),
    .A(_02779_));
 sg13g2_nand3_1 _16359_ (.B(_02767_),
    .C(_02777_),
    .A(_02762_),
    .Y(_02779_));
 sg13g2_a221oi_1 _16360_ (.B2(net7363),
    .C1(net7361),
    .B1(_02779_),
    .A1(_02292_),
    .Y(_02780_),
    .A2(_02753_));
 sg13g2_nand2b_1 _16361_ (.Y(_02781_),
    .B(_01576_),
    .A_N(net7908));
 sg13g2_nand2_1 _16362_ (.Y(_02782_),
    .A(net7908),
    .B(_00620_));
 sg13g2_nand3_1 _16363_ (.B(_02781_),
    .C(_02782_),
    .A(_10980_),
    .Y(_02783_));
 sg13g2_nand2_1 _16364_ (.Y(_02784_),
    .A(net7908),
    .B(_01541_));
 sg13g2_nand2b_1 _16365_ (.Y(_02785_),
    .B(_01506_),
    .A_N(net7908));
 sg13g2_nand4_1 _16366_ (.B(_09150_),
    .C(_02784_),
    .A(net7511),
    .Y(_02786_),
    .D(_02785_));
 sg13g2_nand2_1 _16367_ (.Y(_02787_),
    .A(net7910),
    .B(_01048_));
 sg13g2_nand2b_1 _16368_ (.Y(_02788_),
    .B(_01013_),
    .A_N(net7910));
 sg13g2_nand4_1 _16369_ (.B(_09001_),
    .C(_02787_),
    .A(net7542),
    .Y(_02789_),
    .D(_02788_));
 sg13g2_nand2_1 _16370_ (.Y(_02790_),
    .A(net7914),
    .B(_00978_));
 sg13g2_nand2b_1 _16371_ (.Y(_02791_),
    .B(_00943_),
    .A_N(net7910));
 sg13g2_nand4_1 _16372_ (.B(net7511),
    .C(_02790_),
    .A(net7542),
    .Y(_02792_),
    .D(_02791_));
 sg13g2_nand2_1 _16373_ (.Y(_02793_),
    .A(net7910),
    .B(_00839_));
 sg13g2_nand2b_1 _16374_ (.Y(_02794_),
    .B(_00807_),
    .A_N(net7910));
 sg13g2_nand4_1 _16375_ (.B(net7473),
    .C(_02793_),
    .A(net7542),
    .Y(_02795_),
    .D(_02794_));
 sg13g2_nand2_1 _16376_ (.Y(_02796_),
    .A(net7914),
    .B(_00908_));
 sg13g2_nand2b_1 _16377_ (.Y(_02797_),
    .B(_00872_),
    .A_N(net7914));
 sg13g2_nand4_1 _16378_ (.B(net7464),
    .C(_02796_),
    .A(net7542),
    .Y(_02798_),
    .D(_02797_));
 sg13g2_nand2_1 _16379_ (.Y(_02799_),
    .A(net7908),
    .B(_01400_));
 sg13g2_nand2b_1 _16380_ (.Y(_02800_),
    .B(_01365_),
    .A_N(net7908));
 sg13g2_nand4_1 _16381_ (.B(net7473),
    .C(_02799_),
    .A(net7498),
    .Y(_02801_),
    .D(_02800_));
 sg13g2_nand2_1 _16382_ (.Y(_02802_),
    .A(net7908),
    .B(_01471_));
 sg13g2_nand2b_1 _16383_ (.Y(_02803_),
    .B(_01436_),
    .A_N(net7908));
 sg13g2_nand4_1 _16384_ (.B(net7464),
    .C(_02802_),
    .A(_09150_),
    .Y(_02804_),
    .D(_02803_));
 sg13g2_nand4_1 _16385_ (.B(_02795_),
    .C(_02801_),
    .A(_02789_),
    .Y(_02805_),
    .D(_02804_));
 sg13g2_nand4_1 _16386_ (.B(_02786_),
    .C(_02792_),
    .A(_02783_),
    .Y(_02806_),
    .D(_02798_));
 sg13g2_mux2_1 _16387_ (.A0(_01423_),
    .A1(_00647_),
    .S(net7857),
    .X(_02807_));
 sg13g2_and2_1 _16388_ (.A(net7857),
    .B(_01071_),
    .X(_02808_));
 sg13g2_mux2_1 _16389_ (.A0(_00679_),
    .A1(_00711_),
    .S(net7861),
    .X(_02809_));
 sg13g2_mux2_1 _16390_ (.A0(_00743_),
    .A1(_00775_),
    .S(net7857),
    .X(_02810_));
 sg13g2_mux4_1 _16391_ (.S0(net7810),
    .A0(_02808_),
    .A1(_02809_),
    .A2(_02807_),
    .A3(_02810_),
    .S1(net7829),
    .X(_02811_));
 sg13g2_nor2_1 _16392_ (.A(net7528),
    .B(_02811_),
    .Y(_02812_));
 sg13g2_mux4_1 _16393_ (.S0(net7898),
    .A0(_01084_),
    .A1(_01119_),
    .A2(_01154_),
    .A3(_01189_),
    .S1(net7817),
    .X(_02813_));
 sg13g2_mux4_1 _16394_ (.S0(net7896),
    .A0(_01224_),
    .A1(_01260_),
    .A2(_01295_),
    .A3(_01330_),
    .S1(net7817),
    .X(_02814_));
 sg13g2_or2_1 _16395_ (.X(_02815_),
    .B(_02814_),
    .A(net7445));
 sg13g2_o21ai_1 _16396_ (.B1(_02815_),
    .Y(_02816_),
    .A1(_12139_),
    .A2(_02813_));
 sg13g2_nor4_1 _16397_ (.A(_02805_),
    .B(_02806_),
    .C(_02812_),
    .D(_02816_),
    .Y(_02817_));
 sg13g2_or4_1 _16398_ (.A(_02805_),
    .B(_02806_),
    .C(_02812_),
    .D(_02816_),
    .X(_02818_));
 sg13g2_nand2b_1 _16399_ (.Y(_02819_),
    .B(net7999),
    .A_N(_01653_));
 sg13g2_o21ai_1 _16400_ (.B1(_02819_),
    .Y(_02820_),
    .A1(_01617_),
    .A2(_09260_));
 sg13g2_a221oi_1 _16401_ (.B2(net8005),
    .C1(_02820_),
    .B1(_02818_),
    .A1(net7352),
    .Y(_02821_),
    .A2(net7262));
 sg13g2_nor2_1 _16402_ (.A(net7375),
    .B(_02821_),
    .Y(_02822_));
 sg13g2_a21oi_1 _16403_ (.A1(net6918),
    .A2(_02780_),
    .Y(_02823_),
    .B1(_02822_));
 sg13g2_o21ai_1 _16404_ (.B1(_02823_),
    .Y(_02824_),
    .A1(net6978),
    .A2(_02780_));
 sg13g2_mux2_1 _16405_ (.A0(_01578_),
    .A1(_00621_),
    .S(net7780),
    .X(_02825_));
 sg13g2_nor2_1 _16406_ (.A(_08527_),
    .B(_02825_),
    .Y(_02826_));
 sg13g2_mux2_1 _16407_ (.A0(_01507_),
    .A1(_01542_),
    .S(net7759),
    .X(_02827_));
 sg13g2_nor3_1 _16408_ (.A(net7585),
    .B(net7565),
    .C(_02827_),
    .Y(_02828_));
 sg13g2_mux2_1 _16409_ (.A0(_01437_),
    .A1(_01472_),
    .S(net7759),
    .X(_02829_));
 sg13g2_nor3_1 _16410_ (.A(net7584),
    .B(net7569),
    .C(_02829_),
    .Y(_02830_));
 sg13g2_mux2_1 _16411_ (.A0(_01366_),
    .A1(_01402_),
    .S(net7759),
    .X(_02831_));
 sg13g2_nor3_1 _16412_ (.A(net7584),
    .B(net7560),
    .C(_02831_),
    .Y(_02832_));
 sg13g2_nor4_1 _16413_ (.A(_02826_),
    .B(_02828_),
    .C(_02830_),
    .D(_02832_),
    .Y(_02833_));
 sg13g2_mux4_1 _16414_ (.S0(net7749),
    .A0(_01085_),
    .A1(_01120_),
    .A2(_01155_),
    .A3(_01190_),
    .S1(net7721),
    .X(_02834_));
 sg13g2_inv_1 _16415_ (.Y(_02835_),
    .A(_02834_));
 sg13g2_mux4_1 _16416_ (.S0(net7750),
    .A0(_01226_),
    .A1(_01261_),
    .A2(_01296_),
    .A3(_01331_),
    .S1(net7718),
    .X(_02836_));
 sg13g2_nor2_1 _16417_ (.A(net7586),
    .B(_02836_),
    .Y(_02837_));
 sg13g2_a21oi_1 _16418_ (.A1(net7433),
    .A2(_02835_),
    .Y(_02838_),
    .B1(_02837_));
 sg13g2_mux4_1 _16419_ (.S0(net7753),
    .A0(_00808_),
    .A1(_00840_),
    .A2(_00874_),
    .A3(_00909_),
    .S1(net7735),
    .X(_02839_));
 sg13g2_nand2_1 _16420_ (.Y(_02840_),
    .A(net7606),
    .B(_02839_));
 sg13g2_mux2_1 _16421_ (.A0(_00648_),
    .A1(_00776_),
    .S(net7701),
    .X(_02841_));
 sg13g2_a22oi_1 _16422_ (.Y(_02842_),
    .B1(_02841_),
    .B2(net7436),
    .A2(net7424),
    .A1(_01434_));
 sg13g2_a21oi_1 _16423_ (.A1(_01082_),
    .A2(net7422),
    .Y(_02843_),
    .B1(net7688));
 sg13g2_mux4_1 _16424_ (.S0(net7761),
    .A0(_00944_),
    .A1(_00979_),
    .A2(_01014_),
    .A3(_01050_),
    .S1(net7733),
    .X(_02844_));
 sg13g2_mux2_1 _16425_ (.A0(_00680_),
    .A1(_00712_),
    .S(net7780),
    .X(_02845_));
 sg13g2_a22oi_1 _16426_ (.Y(_02846_),
    .B1(_02845_),
    .B2(_09011_),
    .A2(_08313_),
    .A1(_00744_));
 sg13g2_o21ai_1 _16427_ (.B1(net7700),
    .Y(_02847_),
    .A1(_08946_),
    .A2(_02844_));
 sg13g2_a21o_1 _16428_ (.A2(_02846_),
    .A1(_08946_),
    .B1(_02847_),
    .X(_02848_));
 sg13g2_nand4_1 _16429_ (.B(_02842_),
    .C(_02843_),
    .A(_02840_),
    .Y(_02849_),
    .D(_02848_));
 sg13g2_inv_1 _16430_ (.Y(_02850_),
    .A(_02851_));
 sg13g2_nand3_1 _16431_ (.B(_02838_),
    .C(net7342),
    .A(_02833_),
    .Y(_02851_));
 sg13g2_and3_1 _16432_ (.X(_02852_),
    .A(net7677),
    .B(_08851_),
    .C(_13407_));
 sg13g2_a221oi_1 _16433_ (.B2(net7292),
    .C1(_02852_),
    .B1(_02850_),
    .A1(net7781),
    .Y(_02853_),
    .A2(net7267));
 sg13g2_nand2b_1 _16434_ (.Y(_02854_),
    .B(net8002),
    .A_N(net7980));
 sg13g2_o21ai_1 _16435_ (.B1(_02854_),
    .Y(_02855_),
    .A1(_01619_),
    .A2(_09260_));
 sg13g2_mux2_1 _16436_ (.A0(_01578_),
    .A1(_00621_),
    .S(net7861),
    .X(_02856_));
 sg13g2_nor2_1 _16437_ (.A(net7448),
    .B(_02856_),
    .Y(_02857_));
 sg13g2_mux2_1 _16438_ (.A0(_01507_),
    .A1(_01542_),
    .S(net7912),
    .X(_02858_));
 sg13g2_nor3_1 _16439_ (.A(net7505),
    .B(net7489),
    .C(_02858_),
    .Y(_02859_));
 sg13g2_mux2_1 _16440_ (.A0(_01014_),
    .A1(_01050_),
    .S(net7856),
    .X(_02860_));
 sg13g2_nor3_1 _16441_ (.A(net7538),
    .B(net7522),
    .C(_02860_),
    .Y(_02861_));
 sg13g2_mux2_1 _16442_ (.A0(_00944_),
    .A1(_00979_),
    .S(net7856),
    .X(_02862_));
 sg13g2_nor3_1 _16443_ (.A(net7538),
    .B(net7506),
    .C(_02862_),
    .Y(_02863_));
 sg13g2_nor4_1 _16444_ (.A(_02857_),
    .B(_02859_),
    .C(_02861_),
    .D(_02863_),
    .Y(_02864_));
 sg13g2_mux2_1 _16445_ (.A0(_00808_),
    .A1(_00840_),
    .S(net7856),
    .X(_02865_));
 sg13g2_nor3_1 _16446_ (.A(net7538),
    .B(net7467),
    .C(_02865_),
    .Y(_02866_));
 sg13g2_mux2_1 _16447_ (.A0(_00874_),
    .A1(_00909_),
    .S(net7856),
    .X(_02867_));
 sg13g2_nor3_1 _16448_ (.A(net7538),
    .B(net7458),
    .C(_02867_),
    .Y(_02868_));
 sg13g2_mux2_1 _16449_ (.A0(_01366_),
    .A1(_01402_),
    .S(net7912),
    .X(_02869_));
 sg13g2_nor3_1 _16450_ (.A(net7489),
    .B(net7467),
    .C(_02869_),
    .Y(_02870_));
 sg13g2_mux2_1 _16451_ (.A0(_01437_),
    .A1(_01472_),
    .S(net7912),
    .X(_02871_));
 sg13g2_nor3_1 _16452_ (.A(net7489),
    .B(net7458),
    .C(_02871_),
    .Y(_02872_));
 sg13g2_nor4_1 _16453_ (.A(_02866_),
    .B(_02868_),
    .C(_02870_),
    .D(_02872_),
    .Y(_02873_));
 sg13g2_mux2_1 _16454_ (.A0(_01434_),
    .A1(_00648_),
    .S(net7841),
    .X(_02874_));
 sg13g2_and2_1 _16455_ (.A(net7841),
    .B(_01082_),
    .X(_02875_));
 sg13g2_mux2_1 _16456_ (.A0(_00680_),
    .A1(_00712_),
    .S(net7841),
    .X(_02876_));
 sg13g2_mux2_1 _16457_ (.A0(_00744_),
    .A1(_00776_),
    .S(net7841),
    .X(_02877_));
 sg13g2_mux4_1 _16458_ (.S0(net7813),
    .A0(_02875_),
    .A1(_02876_),
    .A2(_02874_),
    .A3(_02877_),
    .S1(net7821),
    .X(_02878_));
 sg13g2_or2_1 _16459_ (.X(_02879_),
    .B(_02878_),
    .A(net7528));
 sg13g2_mux4_1 _16460_ (.S0(net7900),
    .A0(_01085_),
    .A1(_01120_),
    .A2(_01155_),
    .A3(_01190_),
    .S1(net7819),
    .X(_02880_));
 sg13g2_nor3_1 _16461_ (.A(net7809),
    .B(net7499),
    .C(_02880_),
    .Y(_02881_));
 sg13g2_mux4_1 _16462_ (.S0(net7897),
    .A0(_01226_),
    .A1(_01261_),
    .A2(_01296_),
    .A3(_01331_),
    .S1(net7818),
    .X(_02882_));
 sg13g2_nor2_1 _16463_ (.A(net7445),
    .B(_02882_),
    .Y(_02883_));
 sg13g2_nor2_1 _16464_ (.A(_02881_),
    .B(_02883_),
    .Y(_02884_));
 sg13g2_and4_1 _16465_ (.A(_02864_),
    .B(_02873_),
    .C(_02879_),
    .D(_02884_),
    .X(_02885_));
 sg13g2_nand4_1 _16466_ (.B(_02873_),
    .C(_02879_),
    .A(_02864_),
    .Y(_02886_),
    .D(_02884_));
 sg13g2_a221oi_1 _16467_ (.B2(net8008),
    .C1(_02855_),
    .B1(net7341),
    .A1(net7353),
    .Y(_02887_),
    .A2(net7261));
 sg13g2_nand2_1 _16468_ (.Y(_02888_),
    .A(net6978),
    .B(_02853_));
 sg13g2_o21ai_1 _16469_ (.B1(_02888_),
    .Y(_02889_),
    .A1(net6918),
    .A2(_02853_));
 sg13g2_o21ai_1 _16470_ (.B1(_02889_),
    .Y(_02890_),
    .A1(net7374),
    .A2(_02887_));
 sg13g2_mux2_1 _16471_ (.A0(_01508_),
    .A1(_01543_),
    .S(net7782),
    .X(_02891_));
 sg13g2_nor3_1 _16472_ (.A(net7576),
    .B(net7566),
    .C(_02891_),
    .Y(_02892_));
 sg13g2_mux2_1 _16473_ (.A0(_01579_),
    .A1(_00622_),
    .S(net7782),
    .X(_02893_));
 sg13g2_nor2_1 _16474_ (.A(net7554),
    .B(_02893_),
    .Y(_02894_));
 sg13g2_mux2_1 _16475_ (.A0(_01367_),
    .A1(_01403_),
    .S(net7782),
    .X(_02895_));
 sg13g2_nor3_1 _16476_ (.A(net7576),
    .B(net7557),
    .C(_02895_),
    .Y(_02896_));
 sg13g2_mux2_1 _16477_ (.A0(_01438_),
    .A1(_01473_),
    .S(net7782),
    .X(_02897_));
 sg13g2_nor3_1 _16478_ (.A(_08462_),
    .B(net7570),
    .C(_02897_),
    .Y(_02898_));
 sg13g2_or4_1 _16479_ (.A(_02892_),
    .B(_02894_),
    .C(_02896_),
    .D(_02898_),
    .X(_02899_));
 sg13g2_mux4_1 _16480_ (.S0(net7781),
    .A0(_01227_),
    .A1(_01262_),
    .A2(_01297_),
    .A3(_01332_),
    .S1(net7736),
    .X(_02900_));
 sg13g2_mux4_1 _16481_ (.S0(net7782),
    .A0(_01086_),
    .A1(_01121_),
    .A2(_01156_),
    .A3(_01191_),
    .S1(net7736),
    .X(_02901_));
 sg13g2_nand2b_1 _16482_ (.Y(_02902_),
    .B(net7717),
    .A_N(_02900_));
 sg13g2_o21ai_1 _16483_ (.B1(_02902_),
    .Y(_02903_),
    .A1(net7716),
    .A2(_02901_));
 sg13g2_a21o_1 _16484_ (.A2(_02903_),
    .A1(_08384_),
    .B1(_02899_),
    .X(_02904_));
 sg13g2_mux4_1 _16485_ (.S0(net7782),
    .A0(_00809_),
    .A1(_00841_),
    .A2(_00875_),
    .A3(_00910_),
    .S1(net7743),
    .X(_02905_));
 sg13g2_mux4_1 _16486_ (.S0(net7782),
    .A0(_00945_),
    .A1(_00980_),
    .A2(_01015_),
    .A3(_01051_),
    .S1(net7742),
    .X(_02906_));
 sg13g2_and2_1 _16487_ (.A(_02462_),
    .B(_02906_),
    .X(_02907_));
 sg13g2_and3_1 _16488_ (.X(_02908_),
    .A(_01093_),
    .B(_08305_),
    .C(net7597));
 sg13g2_nand2_1 _16489_ (.Y(_02909_),
    .A(net7717),
    .B(_00777_));
 sg13g2_nand2b_1 _16490_ (.Y(_02910_),
    .B(_00649_),
    .A_N(net7716));
 sg13g2_a21oi_1 _16491_ (.A1(_02909_),
    .A2(_02910_),
    .Y(_02911_),
    .B1(_08291_));
 sg13g2_and3_1 _16492_ (.X(_02912_),
    .A(_01445_),
    .B(_08305_),
    .C(net7596));
 sg13g2_nor4_1 _16493_ (.A(net7688),
    .B(_02908_),
    .C(_02911_),
    .D(_02912_),
    .Y(_02913_));
 sg13g2_mux2_1 _16494_ (.A0(_00681_),
    .A1(_00713_),
    .S(net7781),
    .X(_02914_));
 sg13g2_nor2b_1 _16495_ (.A(net7781),
    .B_N(_00745_),
    .Y(_02915_));
 sg13g2_mux2_1 _16496_ (.A0(_02914_),
    .A1(_02915_),
    .S(net7736),
    .X(_02916_));
 sg13g2_a221oi_1 _16497_ (.B2(_14476_),
    .C1(_02907_),
    .B1(_02916_),
    .A1(net7604),
    .Y(_02917_),
    .A2(_02905_));
 sg13g2_a221oi_1 _16498_ (.B2(_02917_),
    .C1(_02899_),
    .B1(_02913_),
    .A1(_08384_),
    .Y(_02918_),
    .A2(_02903_));
 sg13g2_a21o_1 _16499_ (.A2(_02917_),
    .A1(_02913_),
    .B1(_02904_),
    .X(_02919_));
 sg13g2_a221oi_1 _16500_ (.B2(net7292),
    .C1(_02852_),
    .B1(_02918_),
    .A1(net7736),
    .Y(_02920_),
    .A2(net7267));
 sg13g2_mux2_1 _16501_ (.A0(_01579_),
    .A1(_00622_),
    .S(net7840),
    .X(_02921_));
 sg13g2_nor2_1 _16502_ (.A(net7449),
    .B(_02921_),
    .Y(_02922_));
 sg13g2_mux2_1 _16503_ (.A0(_01508_),
    .A1(_01543_),
    .S(net7840),
    .X(_02923_));
 sg13g2_nor3_1 _16504_ (.A(net7510),
    .B(net7492),
    .C(_02923_),
    .Y(_02924_));
 sg13g2_mux2_1 _16505_ (.A0(_00809_),
    .A1(_00841_),
    .S(net7840),
    .X(_02925_));
 sg13g2_nor3_1 _16506_ (.A(net7536),
    .B(net7466),
    .C(_02925_),
    .Y(_02926_));
 sg13g2_mux2_1 _16507_ (.A0(_00875_),
    .A1(_00910_),
    .S(net7840),
    .X(_02927_));
 sg13g2_nor3_1 _16508_ (.A(net7536),
    .B(_10191_),
    .C(_02927_),
    .Y(_02928_));
 sg13g2_nor4_1 _16509_ (.A(_02922_),
    .B(_02924_),
    .C(_02926_),
    .D(_02928_),
    .Y(_02929_));
 sg13g2_mux2_1 _16510_ (.A0(_01015_),
    .A1(_01051_),
    .S(net7840),
    .X(_02930_));
 sg13g2_nor3_1 _16511_ (.A(net7536),
    .B(_09004_),
    .C(_02930_),
    .Y(_02931_));
 sg13g2_mux2_1 _16512_ (.A0(_00945_),
    .A1(_00980_),
    .S(net7840),
    .X(_02932_));
 sg13g2_nor3_1 _16513_ (.A(net7536),
    .B(net7510),
    .C(_02932_),
    .Y(_02933_));
 sg13g2_mux2_1 _16514_ (.A0(_01367_),
    .A1(_01403_),
    .S(net7840),
    .X(_02934_));
 sg13g2_nor3_1 _16515_ (.A(net7492),
    .B(net7466),
    .C(_02934_),
    .Y(_02935_));
 sg13g2_mux2_1 _16516_ (.A0(_01438_),
    .A1(_01473_),
    .S(net7840),
    .X(_02936_));
 sg13g2_nor3_1 _16517_ (.A(net7492),
    .B(_10191_),
    .C(_02936_),
    .Y(_02937_));
 sg13g2_nor4_1 _16518_ (.A(_02931_),
    .B(_02933_),
    .C(_02935_),
    .D(_02937_),
    .Y(_02938_));
 sg13g2_mux2_1 _16519_ (.A0(_01445_),
    .A1(_00649_),
    .S(net7839),
    .X(_02939_));
 sg13g2_and2_1 _16520_ (.A(net7839),
    .B(_01093_),
    .X(_02940_));
 sg13g2_mux2_1 _16521_ (.A0(_00681_),
    .A1(_00713_),
    .S(net7839),
    .X(_02941_));
 sg13g2_mux2_1 _16522_ (.A0(_00745_),
    .A1(_00777_),
    .S(net7839),
    .X(_02942_));
 sg13g2_mux4_1 _16523_ (.S0(net7812),
    .A0(_02940_),
    .A1(_02941_),
    .A2(_02939_),
    .A3(_02942_),
    .S1(net7821),
    .X(_02943_));
 sg13g2_or2_1 _16524_ (.X(_02944_),
    .B(_02943_),
    .A(_08974_));
 sg13g2_mux4_1 _16525_ (.S0(net7839),
    .A0(_01086_),
    .A1(_01121_),
    .A2(_01156_),
    .A3(_01191_),
    .S1(net7821),
    .X(_02945_));
 sg13g2_nor3_1 _16526_ (.A(net7812),
    .B(_09073_),
    .C(_02945_),
    .Y(_02946_));
 sg13g2_mux4_1 _16527_ (.S0(net7839),
    .A0(_01227_),
    .A1(_01262_),
    .A2(_01297_),
    .A3(_01332_),
    .S1(net7821),
    .X(_02947_));
 sg13g2_nor2_1 _16528_ (.A(_12187_),
    .B(_02947_),
    .Y(_02948_));
 sg13g2_nor2_1 _16529_ (.A(_02946_),
    .B(_02948_),
    .Y(_02949_));
 sg13g2_and4_1 _16530_ (.A(_02929_),
    .B(_02938_),
    .C(_02944_),
    .D(_02949_),
    .X(_02950_));
 sg13g2_nand4_1 _16531_ (.B(_02938_),
    .C(_02944_),
    .A(_02929_),
    .Y(_02951_),
    .D(_02949_));
 sg13g2_nand2b_1 _16532_ (.Y(_02952_),
    .B(net8002),
    .A_N(net7979));
 sg13g2_o21ai_1 _16533_ (.B1(_02952_),
    .Y(_02953_),
    .A1(_01620_),
    .A2(net7481));
 sg13g2_a221oi_1 _16534_ (.B2(net8004),
    .C1(_02953_),
    .B1(net7340),
    .A1(net7353),
    .Y(_02954_),
    .A2(_02919_));
 sg13g2_nand2_1 _16535_ (.Y(_02955_),
    .A(net6978),
    .B(_02920_));
 sg13g2_o21ai_1 _16536_ (.B1(_02955_),
    .Y(_02956_),
    .A1(net6918),
    .A2(_02920_));
 sg13g2_o21ai_1 _16537_ (.B1(_02956_),
    .Y(_02957_),
    .A1(net7374),
    .A2(_02954_));
 sg13g2_mux2_1 _16538_ (.A0(_01509_),
    .A1(_01545_),
    .S(net7754),
    .X(_02958_));
 sg13g2_nor3_1 _16539_ (.A(net7583),
    .B(net7565),
    .C(_02958_),
    .Y(_02959_));
 sg13g2_mux2_1 _16540_ (.A0(_01580_),
    .A1(_00623_),
    .S(net7754),
    .X(_02960_));
 sg13g2_nor2_1 _16541_ (.A(net7553),
    .B(_02960_),
    .Y(_02961_));
 sg13g2_mux2_1 _16542_ (.A0(_01369_),
    .A1(_01404_),
    .S(net7754),
    .X(_02962_));
 sg13g2_nor3_1 _16543_ (.A(net7583),
    .B(net7560),
    .C(_02962_),
    .Y(_02963_));
 sg13g2_mux2_1 _16544_ (.A0(_01439_),
    .A1(_01474_),
    .S(net7754),
    .X(_02964_));
 sg13g2_nor3_1 _16545_ (.A(net7583),
    .B(net7568),
    .C(_02964_),
    .Y(_02965_));
 sg13g2_or4_1 _16546_ (.A(_02959_),
    .B(_02961_),
    .C(_02963_),
    .D(_02965_),
    .X(_02966_));
 sg13g2_mux4_1 _16547_ (.S0(net7750),
    .A0(_01228_),
    .A1(_01263_),
    .A2(_01298_),
    .A3(_01333_),
    .S1(net7718),
    .X(_02967_));
 sg13g2_mux4_1 _16548_ (.S0(net7749),
    .A0(_01087_),
    .A1(_01122_),
    .A2(_01157_),
    .A3(_01193_),
    .S1(net7721),
    .X(_02968_));
 sg13g2_nand2b_1 _16549_ (.Y(_02969_),
    .B(net7702),
    .A_N(_02967_));
 sg13g2_o21ai_1 _16550_ (.B1(_02969_),
    .Y(_02970_),
    .A1(net7702),
    .A2(_02968_));
 sg13g2_a21o_1 _16551_ (.A2(_02970_),
    .A1(net7589),
    .B1(_02966_),
    .X(_02971_));
 sg13g2_mux4_1 _16552_ (.S0(net7753),
    .A0(_00810_),
    .A1(_00842_),
    .A2(_00876_),
    .A3(_00911_),
    .S1(net7719),
    .X(_02972_));
 sg13g2_mux4_1 _16553_ (.S0(net7752),
    .A0(_00946_),
    .A1(_00981_),
    .A2(_01017_),
    .A3(_01052_),
    .S1(net7719),
    .X(_02973_));
 sg13g2_and2_1 _16554_ (.A(net7640),
    .B(_02973_),
    .X(_02974_));
 sg13g2_and3_1 _16555_ (.X(_02975_),
    .A(_01104_),
    .B(net7599),
    .C(net7597));
 sg13g2_nand2_1 _16556_ (.Y(_02976_),
    .A(net7700),
    .B(_00778_));
 sg13g2_nand2b_1 _16557_ (.Y(_02977_),
    .B(_00650_),
    .A_N(net7700));
 sg13g2_a21oi_1 _16558_ (.A1(_02976_),
    .A2(_02977_),
    .Y(_02978_),
    .B1(net7601));
 sg13g2_and3_1 _16559_ (.X(_02979_),
    .A(_01456_),
    .B(net7599),
    .C(net7593));
 sg13g2_nor4_1 _16560_ (.A(net7689),
    .B(_02975_),
    .C(_02978_),
    .D(_02979_),
    .Y(_02980_));
 sg13g2_mux2_1 _16561_ (.A0(_00682_),
    .A1(_00714_),
    .S(net7760),
    .X(_02981_));
 sg13g2_nor2b_1 _16562_ (.A(net7760),
    .B_N(_00746_),
    .Y(_02982_));
 sg13g2_mux2_1 _16563_ (.A0(_02981_),
    .A1(_02982_),
    .S(net7733),
    .X(_02983_));
 sg13g2_a221oi_1 _16564_ (.B2(net7442),
    .C1(_02974_),
    .B1(_02983_),
    .A1(net7606),
    .Y(_02984_),
    .A2(_02972_));
 sg13g2_a221oi_1 _16565_ (.B2(_02984_),
    .C1(_02966_),
    .B1(_02980_),
    .A1(net7589),
    .Y(_02985_),
    .A2(_02970_));
 sg13g2_a21o_1 _16566_ (.A2(_02984_),
    .A1(_02980_),
    .B1(_02971_),
    .X(_02986_));
 sg13g2_a221oi_1 _16567_ (.B2(net7292),
    .C1(net7073),
    .B1(net7339),
    .A1(net7717),
    .Y(_02987_),
    .A2(net7267));
 sg13g2_mux2_1 _16568_ (.A0(_01580_),
    .A1(_00623_),
    .S(net7901),
    .X(_02988_));
 sg13g2_nor2_1 _16569_ (.A(net7448),
    .B(_02988_),
    .Y(_02989_));
 sg13g2_mux2_1 _16570_ (.A0(_01509_),
    .A1(_01545_),
    .S(net7902),
    .X(_02990_));
 sg13g2_nor3_1 _16571_ (.A(net7507),
    .B(net7488),
    .C(_02990_),
    .Y(_02991_));
 sg13g2_mux2_1 _16572_ (.A0(_01017_),
    .A1(_01052_),
    .S(net7901),
    .X(_02992_));
 sg13g2_nor3_1 _16573_ (.A(net7537),
    .B(net7523),
    .C(_02992_),
    .Y(_02993_));
 sg13g2_mux2_1 _16574_ (.A0(_00946_),
    .A1(_00981_),
    .S(net7902),
    .X(_02994_));
 sg13g2_nor3_1 _16575_ (.A(net7537),
    .B(net7507),
    .C(_02994_),
    .Y(_02995_));
 sg13g2_nor4_1 _16576_ (.A(_02989_),
    .B(_02991_),
    .C(_02993_),
    .D(_02995_),
    .Y(_02996_));
 sg13g2_mux2_1 _16577_ (.A0(_00810_),
    .A1(_00842_),
    .S(net7907),
    .X(_02997_));
 sg13g2_nor3_1 _16578_ (.A(net7537),
    .B(net7468),
    .C(_02997_),
    .Y(_02998_));
 sg13g2_mux2_1 _16579_ (.A0(_00876_),
    .A1(_00911_),
    .S(net7907),
    .X(_02999_));
 sg13g2_nor3_1 _16580_ (.A(net7537),
    .B(net7459),
    .C(_02999_),
    .Y(_03000_));
 sg13g2_mux2_1 _16581_ (.A0(_01369_),
    .A1(_01404_),
    .S(net7901),
    .X(_03001_));
 sg13g2_nor3_1 _16582_ (.A(net7488),
    .B(net7468),
    .C(_03001_),
    .Y(_03002_));
 sg13g2_mux2_1 _16583_ (.A0(_01439_),
    .A1(_01474_),
    .S(net7902),
    .X(_03003_));
 sg13g2_nor3_1 _16584_ (.A(net7488),
    .B(net7459),
    .C(_03003_),
    .Y(_03004_));
 sg13g2_nor4_1 _16585_ (.A(_02998_),
    .B(_03000_),
    .C(_03002_),
    .D(_03004_),
    .Y(_03005_));
 sg13g2_mux2_1 _16586_ (.A0(_01456_),
    .A1(_00650_),
    .S(net7837),
    .X(_03006_));
 sg13g2_and2_1 _16587_ (.A(net7837),
    .B(_01104_),
    .X(_03007_));
 sg13g2_mux2_1 _16588_ (.A0(_00682_),
    .A1(_00714_),
    .S(net7838),
    .X(_03008_));
 sg13g2_mux2_1 _16589_ (.A0(_00746_),
    .A1(_00778_),
    .S(net7837),
    .X(_03009_));
 sg13g2_mux4_1 _16590_ (.S0(net7810),
    .A0(_03007_),
    .A1(_03008_),
    .A2(_03006_),
    .A3(_03009_),
    .S1(net7823),
    .X(_03010_));
 sg13g2_or2_1 _16591_ (.X(_03011_),
    .B(_03010_),
    .A(net7528));
 sg13g2_mux4_1 _16592_ (.S0(net7899),
    .A0(_01087_),
    .A1(_01122_),
    .A2(_01157_),
    .A3(_01193_),
    .S1(net7819),
    .X(_03012_));
 sg13g2_nor3_1 _16593_ (.A(net7809),
    .B(net7499),
    .C(_03012_),
    .Y(_03013_));
 sg13g2_mux4_1 _16594_ (.S0(net7899),
    .A0(_01228_),
    .A1(_01263_),
    .A2(_01298_),
    .A3(_01333_),
    .S1(net7819),
    .X(_03014_));
 sg13g2_nor2_1 _16595_ (.A(net7444),
    .B(_03014_),
    .Y(_03015_));
 sg13g2_nor2_1 _16596_ (.A(_03013_),
    .B(_03015_),
    .Y(_03016_));
 sg13g2_and4_1 _16597_ (.A(_02996_),
    .B(_03005_),
    .C(_03011_),
    .D(_03016_),
    .X(_03017_));
 sg13g2_nand4_1 _16598_ (.B(_03005_),
    .C(_03011_),
    .A(_02996_),
    .Y(_03018_),
    .D(_03016_));
 sg13g2_nand2_1 _16599_ (.Y(_03019_),
    .A(_02081_),
    .B(net7999));
 sg13g2_o21ai_1 _16600_ (.B1(_03019_),
    .Y(_03020_),
    .A1(_01621_),
    .A2(net7478));
 sg13g2_a221oi_1 _16601_ (.B2(net8004),
    .C1(_03020_),
    .B1(net7338),
    .A1(net7353),
    .Y(_03021_),
    .A2(_02986_));
 sg13g2_nand2_1 _16602_ (.Y(_03022_),
    .A(net6978),
    .B(_02987_));
 sg13g2_o21ai_1 _16603_ (.B1(_03022_),
    .Y(_03023_),
    .A1(net6918),
    .A2(_02987_));
 sg13g2_o21ai_1 _16604_ (.B1(_03023_),
    .Y(_03024_),
    .A1(net7374),
    .A2(_03021_));
 sg13g2_mux2_1 _16605_ (.A0(_01440_),
    .A1(_01475_),
    .S(net7798),
    .X(_03025_));
 sg13g2_nor3_1 _16606_ (.A(net7576),
    .B(net7570),
    .C(_03025_),
    .Y(_03026_));
 sg13g2_mux2_1 _16607_ (.A0(_01370_),
    .A1(_01405_),
    .S(net7798),
    .X(_03027_));
 sg13g2_nor3_1 _16608_ (.A(net7576),
    .B(net7557),
    .C(_03027_),
    .Y(_03028_));
 sg13g2_mux2_1 _16609_ (.A0(_01510_),
    .A1(_01546_),
    .S(net7798),
    .X(_03029_));
 sg13g2_nor3_1 _16610_ (.A(net7576),
    .B(net7566),
    .C(_03029_),
    .Y(_03030_));
 sg13g2_mux2_1 _16611_ (.A0(_01581_),
    .A1(_00624_),
    .S(net7798),
    .X(_03031_));
 sg13g2_nor2_1 _16612_ (.A(net7554),
    .B(_03031_),
    .Y(_03032_));
 sg13g2_or4_1 _16613_ (.A(_03026_),
    .B(_03028_),
    .C(_03030_),
    .D(_03032_),
    .X(_03033_));
 sg13g2_mux4_1 _16614_ (.S0(net7789),
    .A0(_01229_),
    .A1(_01264_),
    .A2(_01299_),
    .A3(_01334_),
    .S1(net7739),
    .X(_03034_));
 sg13g2_mux4_1 _16615_ (.S0(net7789),
    .A0(_01088_),
    .A1(_01123_),
    .A2(_01158_),
    .A3(_01194_),
    .S1(net7737),
    .X(_03035_));
 sg13g2_nand2b_1 _16616_ (.Y(_03036_),
    .B(net7716),
    .A_N(_03034_));
 sg13g2_o21ai_1 _16617_ (.B1(_03036_),
    .Y(_03037_),
    .A1(net7716),
    .A2(_03035_));
 sg13g2_a21o_1 _16618_ (.A2(_03037_),
    .A1(_08384_),
    .B1(_03033_),
    .X(_03038_));
 sg13g2_mux4_1 _16619_ (.S0(net7798),
    .A0(_00811_),
    .A1(_00843_),
    .A2(_00877_),
    .A3(_00912_),
    .S1(net7739),
    .X(_03039_));
 sg13g2_mux4_1 _16620_ (.S0(net7803),
    .A0(_00947_),
    .A1(_00982_),
    .A2(_01018_),
    .A3(_01053_),
    .S1(net7739),
    .X(_03040_));
 sg13g2_and2_1 _16621_ (.A(_02462_),
    .B(_03040_),
    .X(_03041_));
 sg13g2_and3_1 _16622_ (.X(_03042_),
    .A(_01115_),
    .B(_08305_),
    .C(net7597));
 sg13g2_nand2_1 _16623_ (.Y(_03043_),
    .A(net7716),
    .B(_00779_));
 sg13g2_nand2b_1 _16624_ (.Y(_03044_),
    .B(_00651_),
    .A_N(net7716));
 sg13g2_a21oi_1 _16625_ (.A1(_03043_),
    .A2(_03044_),
    .Y(_03045_),
    .B1(_08291_));
 sg13g2_and3_1 _16626_ (.X(_03046_),
    .A(_01467_),
    .B(_08305_),
    .C(net7596));
 sg13g2_nor4_1 _16627_ (.A(net7688),
    .B(_03042_),
    .C(_03045_),
    .D(_03046_),
    .Y(_03047_));
 sg13g2_mux2_1 _16628_ (.A0(_00683_),
    .A1(_00715_),
    .S(net7782),
    .X(_03048_));
 sg13g2_nor2b_1 _16629_ (.A(net7804),
    .B_N(_00747_),
    .Y(_03049_));
 sg13g2_mux2_1 _16630_ (.A0(_03048_),
    .A1(_03049_),
    .S(net7739),
    .X(_03050_));
 sg13g2_a221oi_1 _16631_ (.B2(_14476_),
    .C1(_03041_),
    .B1(_03050_),
    .A1(net7604),
    .Y(_03051_),
    .A2(_03039_));
 sg13g2_a221oi_1 _16632_ (.B2(_03051_),
    .C1(_03033_),
    .B1(_03047_),
    .A1(_08384_),
    .Y(_03052_),
    .A2(_03037_));
 sg13g2_a21o_1 _16633_ (.A2(_03051_),
    .A1(_03047_),
    .B1(_03038_),
    .X(_03053_));
 sg13g2_a221oi_1 _16634_ (.B2(net7292),
    .C1(_02852_),
    .B1(net7337),
    .A1(net7692),
    .Y(_03054_),
    .A2(net7267));
 sg13g2_mux2_1 _16635_ (.A0(_01581_),
    .A1(_00624_),
    .S(net7853),
    .X(_03055_));
 sg13g2_nor2_1 _16636_ (.A(net7449),
    .B(_03055_),
    .Y(_03056_));
 sg13g2_mux2_1 _16637_ (.A0(_01510_),
    .A1(_01546_),
    .S(net7853),
    .X(_03057_));
 sg13g2_nor3_1 _16638_ (.A(net7510),
    .B(net7491),
    .C(_03057_),
    .Y(_03058_));
 sg13g2_mux2_1 _16639_ (.A0(_01018_),
    .A1(_01053_),
    .S(net7854),
    .X(_03059_));
 sg13g2_nor3_1 _16640_ (.A(net7536),
    .B(_09004_),
    .C(_03059_),
    .Y(_03060_));
 sg13g2_mux2_1 _16641_ (.A0(_00947_),
    .A1(_00982_),
    .S(net7853),
    .X(_03061_));
 sg13g2_nor3_1 _16642_ (.A(net7536),
    .B(net7510),
    .C(_03061_),
    .Y(_03062_));
 sg13g2_nor4_1 _16643_ (.A(_03056_),
    .B(_03058_),
    .C(_03060_),
    .D(_03062_),
    .Y(_03063_));
 sg13g2_mux2_1 _16644_ (.A0(_00811_),
    .A1(_00843_),
    .S(net7853),
    .X(_03064_));
 sg13g2_nor3_1 _16645_ (.A(net7536),
    .B(net7466),
    .C(_03064_),
    .Y(_03065_));
 sg13g2_mux2_1 _16646_ (.A0(_00877_),
    .A1(_00912_),
    .S(net7853),
    .X(_03066_));
 sg13g2_nor3_1 _16647_ (.A(net7536),
    .B(_10191_),
    .C(_03066_),
    .Y(_03067_));
 sg13g2_mux2_1 _16648_ (.A0(_01370_),
    .A1(_01405_),
    .S(net7853),
    .X(_03068_));
 sg13g2_nor3_1 _16649_ (.A(net7491),
    .B(net7466),
    .C(_03068_),
    .Y(_03069_));
 sg13g2_mux2_1 _16650_ (.A0(_01440_),
    .A1(_01475_),
    .S(net7853),
    .X(_03070_));
 sg13g2_nor3_1 _16651_ (.A(net7491),
    .B(_10191_),
    .C(_03070_),
    .Y(_03071_));
 sg13g2_nor4_1 _16652_ (.A(_03065_),
    .B(_03067_),
    .C(_03069_),
    .D(_03071_),
    .Y(_03072_));
 sg13g2_mux2_1 _16653_ (.A0(_01467_),
    .A1(_00651_),
    .S(net7844),
    .X(_03073_));
 sg13g2_and2_1 _16654_ (.A(net7844),
    .B(_01115_),
    .X(_03074_));
 sg13g2_mux2_1 _16655_ (.A0(_00683_),
    .A1(_00715_),
    .S(net7844),
    .X(_03075_));
 sg13g2_mux2_1 _16656_ (.A0(_00747_),
    .A1(_00779_),
    .S(net7844),
    .X(_03076_));
 sg13g2_mux4_1 _16657_ (.S0(net7811),
    .A0(_03074_),
    .A1(_03075_),
    .A2(_03073_),
    .A3(_03076_),
    .S1(net7823),
    .X(_03077_));
 sg13g2_or2_1 _16658_ (.X(_03078_),
    .B(_03077_),
    .A(_08974_));
 sg13g2_mux4_1 _16659_ (.S0(net7845),
    .A0(_01088_),
    .A1(_01123_),
    .A2(_01158_),
    .A3(_01194_),
    .S1(net7822),
    .X(_03079_));
 sg13g2_nor3_1 _16660_ (.A(net7811),
    .B(_09073_),
    .C(_03079_),
    .Y(_03080_));
 sg13g2_mux4_1 _16661_ (.S0(net7853),
    .A0(_01229_),
    .A1(_01264_),
    .A2(_01299_),
    .A3(_01334_),
    .S1(net7822),
    .X(_03081_));
 sg13g2_nor2_1 _16662_ (.A(_12187_),
    .B(_03081_),
    .Y(_03082_));
 sg13g2_nor2_1 _16663_ (.A(_03080_),
    .B(_03082_),
    .Y(_03083_));
 sg13g2_and4_1 _16664_ (.A(_03063_),
    .B(_03072_),
    .C(_03078_),
    .D(_03083_),
    .X(_03084_));
 sg13g2_nand4_1 _16665_ (.B(_03072_),
    .C(_03078_),
    .A(_03063_),
    .Y(_03085_),
    .D(_03083_));
 sg13g2_nand2b_1 _16666_ (.Y(_03086_),
    .B(net8002),
    .A_N(net7978));
 sg13g2_o21ai_1 _16667_ (.B1(_03086_),
    .Y(_03087_),
    .A1(_01622_),
    .A2(_09260_));
 sg13g2_a221oi_1 _16668_ (.B2(net8008),
    .C1(_03087_),
    .B1(net7336),
    .A1(net7353),
    .Y(_03088_),
    .A2(_03053_));
 sg13g2_nand2_1 _16669_ (.Y(_03089_),
    .A(net6978),
    .B(_03054_));
 sg13g2_o21ai_1 _16670_ (.B1(_03089_),
    .Y(_03090_),
    .A1(net6918),
    .A2(_03054_));
 sg13g2_o21ai_1 _16671_ (.B1(_03090_),
    .Y(_03091_),
    .A1(net7374),
    .A2(_03088_));
 sg13g2_mux2_1 _16672_ (.A0(_01512_),
    .A1(_01547_),
    .S(net7755),
    .X(_03092_));
 sg13g2_nor3_1 _16673_ (.A(net7580),
    .B(net7564),
    .C(_03092_),
    .Y(_03093_));
 sg13g2_mux2_1 _16674_ (.A0(_01371_),
    .A1(_01406_),
    .S(net7755),
    .X(_03094_));
 sg13g2_nor3_1 _16675_ (.A(net7580),
    .B(net7559),
    .C(_03094_),
    .Y(_03095_));
 sg13g2_mux2_1 _16676_ (.A0(_01582_),
    .A1(_00625_),
    .S(net7755),
    .X(_03096_));
 sg13g2_nor2_1 _16677_ (.A(net7553),
    .B(_03096_),
    .Y(_03097_));
 sg13g2_mux2_1 _16678_ (.A0(_01441_),
    .A1(_01476_),
    .S(net7755),
    .X(_03098_));
 sg13g2_nor3_1 _16679_ (.A(net7580),
    .B(net7567),
    .C(_03098_),
    .Y(_03099_));
 sg13g2_or4_1 _16680_ (.A(_03093_),
    .B(_03095_),
    .C(_03097_),
    .D(_03099_),
    .X(_03100_));
 sg13g2_mux4_1 _16681_ (.S0(net7751),
    .A0(_01230_),
    .A1(_01265_),
    .A2(_01300_),
    .A3(_01336_),
    .S1(net7720),
    .X(_03101_));
 sg13g2_mux4_1 _16682_ (.S0(net7750),
    .A0(_01089_),
    .A1(_01124_),
    .A2(_01160_),
    .A3(_01195_),
    .S1(net7718),
    .X(_03102_));
 sg13g2_nand2b_1 _16683_ (.Y(_03103_),
    .B(net7698),
    .A_N(_03101_));
 sg13g2_o21ai_1 _16684_ (.B1(_03103_),
    .Y(_03104_),
    .A1(net7698),
    .A2(_03102_));
 sg13g2_a21oi_1 _16685_ (.A1(net7589),
    .A2(_03104_),
    .Y(_03105_),
    .B1(_03100_));
 sg13g2_mux4_1 _16686_ (.S0(net7764),
    .A0(_00812_),
    .A1(_00844_),
    .A2(_00878_),
    .A3(_00913_),
    .S1(net7722),
    .X(_03106_));
 sg13g2_and2_1 _16687_ (.A(_08255_),
    .B(_03106_),
    .X(_03107_));
 sg13g2_nand2_1 _16688_ (.Y(_03108_),
    .A(net7705),
    .B(_00780_));
 sg13g2_nand2b_1 _16689_ (.Y(_03109_),
    .B(_00652_),
    .A_N(net7705));
 sg13g2_a21oi_1 _16690_ (.A1(_03108_),
    .A2(_03109_),
    .Y(_03110_),
    .B1(net7601));
 sg13g2_nand3b_1 _16691_ (.B(net7764),
    .C(_01126_),
    .Y(_03111_),
    .A_N(net7722));
 sg13g2_nand3b_1 _16692_ (.B(_01478_),
    .C(net7722),
    .Y(_03112_),
    .A_N(net7764));
 sg13g2_a21oi_1 _16693_ (.A1(_03111_),
    .A2(_03112_),
    .Y(_03113_),
    .B1(_08306_));
 sg13g2_nor4_1 _16694_ (.A(net7687),
    .B(_03107_),
    .C(_03110_),
    .D(_03113_),
    .Y(_03114_));
 sg13g2_mux4_1 _16695_ (.S0(net7759),
    .A0(_00948_),
    .A1(_00984_),
    .A2(_01019_),
    .A3(_01054_),
    .S1(net7730),
    .X(_03115_));
 sg13g2_nand2b_1 _16696_ (.Y(_03116_),
    .B(net7692),
    .A_N(_03115_));
 sg13g2_mux2_1 _16697_ (.A0(_00684_),
    .A1(_00716_),
    .S(net7753),
    .X(_03117_));
 sg13g2_a221oi_1 _16698_ (.B2(net7519),
    .C1(net7692),
    .B1(_03117_),
    .A1(_00748_),
    .Y(_03118_),
    .A2(net7593));
 sg13g2_nand3b_1 _16699_ (.B(net7701),
    .C(_03116_),
    .Y(_03119_),
    .A_N(_03118_));
 sg13g2_nand2_1 _16700_ (.Y(_03120_),
    .A(_03114_),
    .B(_03119_));
 sg13g2_a221oi_1 _16701_ (.B2(_03119_),
    .C1(_03100_),
    .B1(_03114_),
    .A1(net7589),
    .Y(_03121_),
    .A2(_03104_));
 sg13g2_nand2_1 _16702_ (.Y(_03122_),
    .A(_03105_),
    .B(_03120_));
 sg13g2_a221oi_1 _16703_ (.B2(net7292),
    .C1(net7073),
    .B1(net7335),
    .A1(net7688),
    .Y(_03123_),
    .A2(net7267));
 sg13g2_mux2_1 _16704_ (.A0(_00684_),
    .A1(_00716_),
    .S(net7861),
    .X(_03124_));
 sg13g2_nor2_1 _16705_ (.A(net7505),
    .B(_03124_),
    .Y(_03125_));
 sg13g2_mux2_1 _16706_ (.A0(_00748_),
    .A1(_00780_),
    .S(net7857),
    .X(_03126_));
 sg13g2_nor2_1 _16707_ (.A(net7522),
    .B(_03126_),
    .Y(_03127_));
 sg13g2_mux2_1 _16708_ (.A0(_01478_),
    .A1(_00652_),
    .S(net7857),
    .X(_03128_));
 sg13g2_a221oi_1 _16709_ (.B2(net7829),
    .C1(net7810),
    .B1(_03128_),
    .A1(_01126_),
    .Y(_03129_),
    .A2(_08988_));
 sg13g2_nor4_1 _16710_ (.A(net7528),
    .B(_03125_),
    .C(_03127_),
    .D(_03129_),
    .Y(_03130_));
 sg13g2_mux2_1 _16711_ (.A0(_01300_),
    .A1(_01336_),
    .S(net7896),
    .X(_03131_));
 sg13g2_nor2_1 _16712_ (.A(net7523),
    .B(_03131_),
    .Y(_03132_));
 sg13g2_mux2_1 _16713_ (.A0(_01089_),
    .A1(_01124_),
    .S(net7896),
    .X(_03133_));
 sg13g2_nor2_1 _16714_ (.A(net7468),
    .B(_03133_),
    .Y(_03134_));
 sg13g2_mux2_1 _16715_ (.A0(_01160_),
    .A1(_01195_),
    .S(net7896),
    .X(_03135_));
 sg13g2_nor2_1 _16716_ (.A(net7459),
    .B(_03135_),
    .Y(_03136_));
 sg13g2_mux2_1 _16717_ (.A0(_01230_),
    .A1(_01265_),
    .S(net7896),
    .X(_03137_));
 sg13g2_o21ai_1 _16718_ (.B1(net7503),
    .Y(_03138_),
    .A1(net7507),
    .A2(_03137_));
 sg13g2_nor4_1 _16719_ (.A(_03132_),
    .B(_03134_),
    .C(_03136_),
    .D(_03138_),
    .Y(_03139_));
 sg13g2_mux2_1 _16720_ (.A0(_01582_),
    .A1(_00625_),
    .S(net7909),
    .X(_03140_));
 sg13g2_nand2_1 _16721_ (.Y(_03141_),
    .A(_10980_),
    .B(_03140_));
 sg13g2_mux2_1 _16722_ (.A0(_01512_),
    .A1(_01547_),
    .S(net7903),
    .X(_03142_));
 sg13g2_nand3_1 _16723_ (.B(net7498),
    .C(_03142_),
    .A(net7511),
    .Y(_03143_));
 sg13g2_mux2_1 _16724_ (.A0(_01441_),
    .A1(_01476_),
    .S(net7909),
    .X(_03144_));
 sg13g2_nand3_1 _16725_ (.B(net7464),
    .C(_03144_),
    .A(net7498),
    .Y(_03145_));
 sg13g2_mux2_1 _16726_ (.A0(_01371_),
    .A1(_01406_),
    .S(net7909),
    .X(_03146_));
 sg13g2_nand3_1 _16727_ (.B(net7473),
    .C(_03146_),
    .A(net7498),
    .Y(_03147_));
 sg13g2_mux2_1 _16728_ (.A0(_00878_),
    .A1(_00913_),
    .S(net7911),
    .X(_03148_));
 sg13g2_nand3_1 _16729_ (.B(net7464),
    .C(_03148_),
    .A(net7541),
    .Y(_03149_));
 sg13g2_mux2_1 _16730_ (.A0(_00812_),
    .A1(_00844_),
    .S(net7911),
    .X(_03150_));
 sg13g2_nand3_1 _16731_ (.B(net7473),
    .C(_03150_),
    .A(net7541),
    .Y(_03151_));
 sg13g2_mux2_1 _16732_ (.A0(_00948_),
    .A1(_00984_),
    .S(net7912),
    .X(_03152_));
 sg13g2_nand3_1 _16733_ (.B(net7511),
    .C(_03152_),
    .A(net7542),
    .Y(_03153_));
 sg13g2_mux2_1 _16734_ (.A0(_01019_),
    .A1(_01054_),
    .S(net7911),
    .X(_03154_));
 sg13g2_nand3_1 _16735_ (.B(_09001_),
    .C(_03154_),
    .A(net7541),
    .Y(_03155_));
 sg13g2_nand4_1 _16736_ (.B(_03145_),
    .C(_03147_),
    .A(_03141_),
    .Y(_03156_),
    .D(_03153_));
 sg13g2_nand4_1 _16737_ (.B(_03149_),
    .C(_03151_),
    .A(_03143_),
    .Y(_03157_),
    .D(_03155_));
 sg13g2_nor4_1 _16738_ (.A(_03130_),
    .B(_03139_),
    .C(_03156_),
    .D(_03157_),
    .Y(_03158_));
 sg13g2_or4_1 _16739_ (.A(_03130_),
    .B(_03139_),
    .C(_03156_),
    .D(_03157_),
    .X(_03159_));
 sg13g2_nand2b_1 _16740_ (.Y(_03160_),
    .B(net7998),
    .A_N(_01658_));
 sg13g2_o21ai_1 _16741_ (.B1(_03160_),
    .Y(_03161_),
    .A1(_01623_),
    .A2(_09260_));
 sg13g2_a221oi_1 _16742_ (.B2(net8007),
    .C1(_03161_),
    .B1(net7334),
    .A1(_09275_),
    .Y(_03162_),
    .A2(_03122_));
 sg13g2_nand2_1 _16743_ (.Y(_03163_),
    .A(net6979),
    .B(net7030));
 sg13g2_o21ai_1 _16744_ (.B1(_03163_),
    .Y(_03164_),
    .A1(net6919),
    .A2(net7030));
 sg13g2_o21ai_1 _16745_ (.B1(_03164_),
    .Y(_03165_),
    .A1(net7375),
    .A2(_03162_));
 sg13g2_mux2_1 _16746_ (.A0(_01442_),
    .A1(_01477_),
    .S(net7785),
    .X(_03166_));
 sg13g2_nor3_1 _16747_ (.A(_08462_),
    .B(net7570),
    .C(_03166_),
    .Y(_03167_));
 sg13g2_mux2_1 _16748_ (.A0(_01583_),
    .A1(_00626_),
    .S(net7787),
    .X(_03168_));
 sg13g2_nor2_1 _16749_ (.A(net7554),
    .B(_03168_),
    .Y(_03169_));
 sg13g2_mux2_1 _16750_ (.A0(_01513_),
    .A1(_01548_),
    .S(net7785),
    .X(_03170_));
 sg13g2_nor3_1 _16751_ (.A(_08462_),
    .B(net7566),
    .C(_03170_),
    .Y(_03171_));
 sg13g2_mux2_1 _16752_ (.A0(_01372_),
    .A1(_01407_),
    .S(net7785),
    .X(_03172_));
 sg13g2_nor3_1 _16753_ (.A(_08462_),
    .B(net7557),
    .C(_03172_),
    .Y(_03173_));
 sg13g2_nor4_1 _16754_ (.A(_03167_),
    .B(_03169_),
    .C(_03171_),
    .D(_03173_),
    .Y(_03174_));
 sg13g2_mux4_1 _16755_ (.S0(net7779),
    .A0(_01231_),
    .A1(_01266_),
    .A2(_01301_),
    .A3(_01337_),
    .S1(net7729),
    .X(_03175_));
 sg13g2_nor2_1 _16756_ (.A(net7587),
    .B(_03175_),
    .Y(_03176_));
 sg13g2_mux4_1 _16757_ (.S0(net7779),
    .A0(_01090_),
    .A1(_01125_),
    .A2(_01161_),
    .A3(_01196_),
    .S1(net7729),
    .X(_03177_));
 sg13g2_inv_1 _16758_ (.Y(_03178_),
    .A(_03177_));
 sg13g2_a21oi_1 _16759_ (.A1(net7434),
    .A2(_03178_),
    .Y(_03179_),
    .B1(_03176_));
 sg13g2_mux4_1 _16760_ (.S0(net7787),
    .A0(_00813_),
    .A1(_00845_),
    .A2(_00879_),
    .A3(_00914_),
    .S1(net7742),
    .X(_03180_));
 sg13g2_nand2_1 _16761_ (.Y(_03181_),
    .A(net7603),
    .B(_03180_));
 sg13g2_mux2_1 _16762_ (.A0(_00653_),
    .A1(_00781_),
    .S(net7704),
    .X(_03182_));
 sg13g2_a22oi_1 _16763_ (.Y(_03183_),
    .B1(_03182_),
    .B2(net7435),
    .A2(net7424),
    .A1(_01489_));
 sg13g2_a21oi_1 _16764_ (.A1(_01137_),
    .A2(net7423),
    .Y(_03184_),
    .B1(net7686));
 sg13g2_mux4_1 _16765_ (.S0(net7788),
    .A0(_00949_),
    .A1(_00985_),
    .A2(_01020_),
    .A3(_01055_),
    .S1(net7742),
    .X(_03185_));
 sg13g2_mux2_1 _16766_ (.A0(_00685_),
    .A1(_00717_),
    .S(net7788),
    .X(_03186_));
 sg13g2_a22oi_1 _16767_ (.Y(_03187_),
    .B1(_03186_),
    .B2(net7518),
    .A2(net7594),
    .A1(_00749_));
 sg13g2_o21ai_1 _16768_ (.B1(net7704),
    .Y(_03188_),
    .A1(net7534),
    .A2(_03185_));
 sg13g2_a21o_1 _16769_ (.A2(_03187_),
    .A1(net7534),
    .B1(_03188_),
    .X(_03189_));
 sg13g2_nand4_1 _16770_ (.B(_03183_),
    .C(_03184_),
    .A(_03181_),
    .Y(_03190_),
    .D(_03189_));
 sg13g2_inv_1 _16771_ (.Y(_03191_),
    .A(_03192_));
 sg13g2_nand3_1 _16772_ (.B(_03179_),
    .C(_03190_),
    .A(_03174_),
    .Y(_03192_));
 sg13g2_a221oi_1 _16773_ (.B2(net7292),
    .C1(net7073),
    .B1(_03191_),
    .A1(net7684),
    .Y(_03193_),
    .A2(net7268));
 sg13g2_nand2b_1 _16774_ (.Y(_03194_),
    .B(net8002),
    .A_N(_01659_));
 sg13g2_o21ai_1 _16775_ (.B1(_03194_),
    .Y(_03195_),
    .A1(_01624_),
    .A2(net7481));
 sg13g2_mux2_1 _16776_ (.A0(_01583_),
    .A1(_00626_),
    .S(net7860),
    .X(_03196_));
 sg13g2_nor2_1 _16777_ (.A(net7449),
    .B(_03196_),
    .Y(_03197_));
 sg13g2_mux2_1 _16778_ (.A0(_01513_),
    .A1(_01548_),
    .S(net7894),
    .X(_03198_));
 sg13g2_nor3_1 _16779_ (.A(net7510),
    .B(net7492),
    .C(_03198_),
    .Y(_03199_));
 sg13g2_mux2_1 _16780_ (.A0(_01020_),
    .A1(_01055_),
    .S(net7859),
    .X(_03200_));
 sg13g2_nor3_1 _16781_ (.A(net7535),
    .B(_09004_),
    .C(_03200_),
    .Y(_03201_));
 sg13g2_mux2_1 _16782_ (.A0(_00949_),
    .A1(_00985_),
    .S(net7859),
    .X(_03202_));
 sg13g2_nor3_1 _16783_ (.A(net7535),
    .B(net7510),
    .C(_03202_),
    .Y(_03203_));
 sg13g2_nor4_1 _16784_ (.A(_03197_),
    .B(_03199_),
    .C(_03201_),
    .D(_03203_),
    .Y(_03204_));
 sg13g2_mux2_1 _16785_ (.A0(_00813_),
    .A1(_00845_),
    .S(net7859),
    .X(_03205_));
 sg13g2_nor3_1 _16786_ (.A(net7535),
    .B(net7465),
    .C(_03205_),
    .Y(_03206_));
 sg13g2_mux2_1 _16787_ (.A0(_00879_),
    .A1(_00914_),
    .S(net7859),
    .X(_03207_));
 sg13g2_nor3_1 _16788_ (.A(net7535),
    .B(net7461),
    .C(_03207_),
    .Y(_03208_));
 sg13g2_mux2_1 _16789_ (.A0(_01372_),
    .A1(_01407_),
    .S(net7895),
    .X(_03209_));
 sg13g2_nor3_1 _16790_ (.A(net7491),
    .B(net7465),
    .C(_03209_),
    .Y(_03210_));
 sg13g2_mux2_1 _16791_ (.A0(_01442_),
    .A1(_01477_),
    .S(net7895),
    .X(_03211_));
 sg13g2_nor3_1 _16792_ (.A(net7491),
    .B(net7461),
    .C(_03211_),
    .Y(_03212_));
 sg13g2_nor4_1 _16793_ (.A(_03206_),
    .B(_03208_),
    .C(_03210_),
    .D(_03212_),
    .Y(_03213_));
 sg13g2_mux2_1 _16794_ (.A0(_01489_),
    .A1(_00653_),
    .S(net7859),
    .X(_03214_));
 sg13g2_and2_1 _16795_ (.A(net7859),
    .B(_01137_),
    .X(_03215_));
 sg13g2_mux2_1 _16796_ (.A0(_00685_),
    .A1(_00717_),
    .S(net7859),
    .X(_03216_));
 sg13g2_mux2_1 _16797_ (.A0(_00749_),
    .A1(_00781_),
    .S(net7859),
    .X(_03217_));
 sg13g2_mux4_1 _16798_ (.S0(net7812),
    .A0(_03215_),
    .A1(_03216_),
    .A2(_03214_),
    .A3(_03217_),
    .S1(net7834),
    .X(_03218_));
 sg13g2_or2_1 _16799_ (.X(_03219_),
    .B(_03218_),
    .A(net7529));
 sg13g2_mux4_1 _16800_ (.S0(net7895),
    .A0(_01090_),
    .A1(_01125_),
    .A2(_01161_),
    .A3(_01196_),
    .S1(net7834),
    .X(_03220_));
 sg13g2_nor3_1 _16801_ (.A(net7816),
    .B(net7500),
    .C(_03220_),
    .Y(_03221_));
 sg13g2_mux4_1 _16802_ (.S0(net7867),
    .A0(_01231_),
    .A1(_01266_),
    .A2(_01301_),
    .A3(_01337_),
    .S1(net7834),
    .X(_03222_));
 sg13g2_nor2_1 _16803_ (.A(net7443),
    .B(_03222_),
    .Y(_03223_));
 sg13g2_nor2_1 _16804_ (.A(_03221_),
    .B(_03223_),
    .Y(_03224_));
 sg13g2_and4_1 _16805_ (.A(_03204_),
    .B(_03213_),
    .C(_03219_),
    .D(_03224_),
    .X(_03225_));
 sg13g2_nand4_1 _16806_ (.B(_03213_),
    .C(_03219_),
    .A(_03204_),
    .Y(_03226_),
    .D(_03224_));
 sg13g2_a221oi_1 _16807_ (.B2(net8008),
    .C1(_03195_),
    .B1(net7333),
    .A1(net7353),
    .Y(_03227_),
    .A2(_03192_));
 sg13g2_nand2_1 _16808_ (.Y(_03228_),
    .A(net6979),
    .B(_03193_));
 sg13g2_o21ai_1 _16809_ (.B1(_03228_),
    .Y(_03229_),
    .A1(net6919),
    .A2(_03193_));
 sg13g2_o21ai_1 _16810_ (.B1(_03229_),
    .Y(_03230_),
    .A1(net7374),
    .A2(_03227_));
 sg13g2_mux2_1 _16811_ (.A0(_01373_),
    .A1(_01408_),
    .S(net7758),
    .X(_03231_));
 sg13g2_nor3_1 _16812_ (.A(net7580),
    .B(net7559),
    .C(_03231_),
    .Y(_03232_));
 sg13g2_mux2_1 _16813_ (.A0(_01584_),
    .A1(_00627_),
    .S(net7758),
    .X(_03233_));
 sg13g2_nor2_1 _16814_ (.A(net7551),
    .B(_03233_),
    .Y(_03234_));
 sg13g2_mux2_1 _16815_ (.A0(_01514_),
    .A1(_01549_),
    .S(net7758),
    .X(_03235_));
 sg13g2_nor3_1 _16816_ (.A(net7580),
    .B(net7565),
    .C(_03235_),
    .Y(_03236_));
 sg13g2_mux2_1 _16817_ (.A0(_01443_),
    .A1(_01479_),
    .S(net7758),
    .X(_03237_));
 sg13g2_nor3_1 _16818_ (.A(net7580),
    .B(net7567),
    .C(_03237_),
    .Y(_03238_));
 sg13g2_nor4_1 _16819_ (.A(_03232_),
    .B(_03234_),
    .C(_03236_),
    .D(_03238_),
    .Y(_03239_));
 sg13g2_mux4_1 _16820_ (.S0(net7752),
    .A0(_01232_),
    .A1(_01267_),
    .A2(_01303_),
    .A3(_01338_),
    .S1(net7719),
    .X(_03240_));
 sg13g2_nor2_1 _16821_ (.A(net7586),
    .B(_03240_),
    .Y(_03241_));
 sg13g2_mux4_1 _16822_ (.S0(net7752),
    .A0(_01091_),
    .A1(_01127_),
    .A2(_01162_),
    .A3(_01197_),
    .S1(net7719),
    .X(_03242_));
 sg13g2_inv_1 _16823_ (.Y(_03243_),
    .A(_03242_));
 sg13g2_a21oi_1 _16824_ (.A1(net7433),
    .A2(_03243_),
    .Y(_03244_),
    .B1(_03241_));
 sg13g2_mux4_1 _16825_ (.S0(net7764),
    .A0(_00814_),
    .A1(_00846_),
    .A2(_00880_),
    .A3(_00915_),
    .S1(net7722),
    .X(_03245_));
 sg13g2_nand2_1 _16826_ (.Y(_03246_),
    .A(net7605),
    .B(_03245_));
 sg13g2_mux2_1 _16827_ (.A0(_00654_),
    .A1(_00782_),
    .S(_01900_),
    .X(_03247_));
 sg13g2_a22oi_1 _16828_ (.Y(_03248_),
    .B1(_03247_),
    .B2(net7436),
    .A2(net7424),
    .A1(_01500_));
 sg13g2_a21oi_1 _16829_ (.A1(_01148_),
    .A2(net7422),
    .Y(_03249_),
    .B1(net7687));
 sg13g2_mux4_1 _16830_ (.S0(net7764),
    .A0(_00951_),
    .A1(_00986_),
    .A2(_01021_),
    .A3(_01056_),
    .S1(net7722),
    .X(_03250_));
 sg13g2_mux2_1 _16831_ (.A0(_00686_),
    .A1(_00718_),
    .S(net7764),
    .X(_03251_));
 sg13g2_a22oi_1 _16832_ (.Y(_03252_),
    .B1(_03251_),
    .B2(net7519),
    .A2(net7593),
    .A1(_00750_));
 sg13g2_o21ai_1 _16833_ (.B1(_01900_),
    .Y(_03253_),
    .A1(net7532),
    .A2(_03250_));
 sg13g2_a21o_1 _16834_ (.A2(_03252_),
    .A1(net7532),
    .B1(_03253_),
    .X(_03254_));
 sg13g2_nand4_1 _16835_ (.B(_03248_),
    .C(_03249_),
    .A(_03246_),
    .Y(_03255_),
    .D(_03254_));
 sg13g2_and3_1 _16836_ (.X(_03256_),
    .A(_03239_),
    .B(_03244_),
    .C(_03255_));
 sg13g2_a221oi_1 _16837_ (.B2(_08639_),
    .C1(_02852_),
    .B1(_03256_),
    .A1(net7683),
    .Y(_03257_),
    .A2(net7268));
 sg13g2_mux2_1 _16838_ (.A0(_01500_),
    .A1(_00654_),
    .S(net7857),
    .X(_03258_));
 sg13g2_a22oi_1 _16839_ (.Y(_03259_),
    .B1(_03258_),
    .B2(net7829),
    .A2(_08988_),
    .A1(_01148_));
 sg13g2_nand2b_1 _16840_ (.Y(_03260_),
    .B(net7861),
    .A_N(_00718_));
 sg13g2_o21ai_1 _16841_ (.B1(_03260_),
    .Y(_03261_),
    .A1(net7861),
    .A2(_00686_));
 sg13g2_mux2_1 _16842_ (.A0(_00750_),
    .A1(_00782_),
    .S(net7857),
    .X(_03262_));
 sg13g2_o21ai_1 _16843_ (.B1(_08973_),
    .Y(_03263_),
    .A1(net7522),
    .A2(_03262_));
 sg13g2_a221oi_1 _16844_ (.B2(_09026_),
    .C1(_03263_),
    .B1(_03261_),
    .A1(net7485),
    .Y(_03264_),
    .A2(_03259_));
 sg13g2_mux2_1 _16845_ (.A0(_01303_),
    .A1(_01338_),
    .S(net7900),
    .X(_03265_));
 sg13g2_nor2_1 _16846_ (.A(net7523),
    .B(_03265_),
    .Y(_03266_));
 sg13g2_mux2_1 _16847_ (.A0(_01091_),
    .A1(_01127_),
    .S(net7898),
    .X(_03267_));
 sg13g2_nor2_1 _16848_ (.A(net7470),
    .B(_03267_),
    .Y(_03268_));
 sg13g2_mux2_1 _16849_ (.A0(_01162_),
    .A1(_01197_),
    .S(net7898),
    .X(_03269_));
 sg13g2_nor2_1 _16850_ (.A(net7460),
    .B(_03269_),
    .Y(_03270_));
 sg13g2_mux2_1 _16851_ (.A0(_01232_),
    .A1(_01267_),
    .S(net7898),
    .X(_03271_));
 sg13g2_o21ai_1 _16852_ (.B1(net7503),
    .Y(_03272_),
    .A1(net7507),
    .A2(_03271_));
 sg13g2_nor4_1 _16853_ (.A(_03266_),
    .B(_03268_),
    .C(_03270_),
    .D(_03272_),
    .Y(_03273_));
 sg13g2_mux2_1 _16854_ (.A0(_01584_),
    .A1(_00627_),
    .S(net7909),
    .X(_03274_));
 sg13g2_nand2_1 _16855_ (.Y(_03275_),
    .A(_10980_),
    .B(_03274_));
 sg13g2_mux2_1 _16856_ (.A0(_01514_),
    .A1(_01549_),
    .S(net7909),
    .X(_03276_));
 sg13g2_nand3_1 _16857_ (.B(net7498),
    .C(_03276_),
    .A(net7511),
    .Y(_03277_));
 sg13g2_mux2_1 _16858_ (.A0(_01443_),
    .A1(_01479_),
    .S(net7909),
    .X(_03278_));
 sg13g2_nand3_1 _16859_ (.B(net7464),
    .C(_03278_),
    .A(net7498),
    .Y(_03279_));
 sg13g2_mux2_1 _16860_ (.A0(_01373_),
    .A1(_01408_),
    .S(net7909),
    .X(_03280_));
 sg13g2_nand3_1 _16861_ (.B(net7473),
    .C(_03280_),
    .A(net7498),
    .Y(_03281_));
 sg13g2_mux2_1 _16862_ (.A0(_00880_),
    .A1(_00915_),
    .S(net7910),
    .X(_03282_));
 sg13g2_nand3_1 _16863_ (.B(net7464),
    .C(_03282_),
    .A(net7541),
    .Y(_03283_));
 sg13g2_mux2_1 _16864_ (.A0(_00814_),
    .A1(_00846_),
    .S(net7910),
    .X(_03284_));
 sg13g2_nand3_1 _16865_ (.B(net7473),
    .C(_03284_),
    .A(net7541),
    .Y(_03285_));
 sg13g2_mux2_1 _16866_ (.A0(_00951_),
    .A1(_00986_),
    .S(net7911),
    .X(_03286_));
 sg13g2_nand3_1 _16867_ (.B(net7511),
    .C(_03286_),
    .A(net7542),
    .Y(_03287_));
 sg13g2_mux2_1 _16868_ (.A0(_01021_),
    .A1(_01056_),
    .S(net7910),
    .X(_03288_));
 sg13g2_nand3_1 _16869_ (.B(_09001_),
    .C(_03288_),
    .A(net7541),
    .Y(_03289_));
 sg13g2_nand4_1 _16870_ (.B(_03279_),
    .C(_03281_),
    .A(_03275_),
    .Y(_03290_),
    .D(_03287_));
 sg13g2_nand4_1 _16871_ (.B(_03283_),
    .C(_03285_),
    .A(_03277_),
    .Y(_03291_),
    .D(_03289_));
 sg13g2_nor4_1 _16872_ (.A(_03264_),
    .B(_03273_),
    .C(_03290_),
    .D(_03291_),
    .Y(_03292_));
 sg13g2_or4_1 _16873_ (.A(_03264_),
    .B(_03273_),
    .C(_03290_),
    .D(_03291_),
    .X(_03293_));
 sg13g2_nand2b_1 _16874_ (.Y(_03294_),
    .B(net7998),
    .A_N(_01661_));
 sg13g2_o21ai_1 _16875_ (.B1(_03294_),
    .Y(_03295_),
    .A1(_01625_),
    .A2(_09260_));
 sg13g2_a21oi_1 _16876_ (.A1(_00541_),
    .A2(net7332),
    .Y(_03296_),
    .B1(_03295_));
 sg13g2_o21ai_1 _16877_ (.B1(_03296_),
    .Y(_03297_),
    .A1(_09277_),
    .A2(_03256_));
 sg13g2_nand2_1 _16878_ (.Y(_03298_),
    .A(net7384),
    .B(_03297_));
 sg13g2_nand2_1 _16879_ (.Y(_03299_),
    .A(_08228_),
    .B(_03257_));
 sg13g2_o21ai_1 _16880_ (.B1(_03299_),
    .Y(_03300_),
    .A1(net6917),
    .A2(_03257_));
 sg13g2_nand2_1 _16881_ (.Y(_03301_),
    .A(_03298_),
    .B(_03300_));
 sg13g2_mux2_1 _16882_ (.A0(_01374_),
    .A1(_01409_),
    .S(net7783),
    .X(_03302_));
 sg13g2_nor3_1 _16883_ (.A(net7574),
    .B(net7558),
    .C(_03302_),
    .Y(_03303_));
 sg13g2_mux2_1 _16884_ (.A0(_01585_),
    .A1(_00628_),
    .S(net7783),
    .X(_03304_));
 sg13g2_nor2_1 _16885_ (.A(net7556),
    .B(_03304_),
    .Y(_03305_));
 sg13g2_mux2_1 _16886_ (.A0(_01515_),
    .A1(_01550_),
    .S(net7783),
    .X(_03306_));
 sg13g2_nor3_1 _16887_ (.A(net7574),
    .B(net7562),
    .C(_03306_),
    .Y(_03307_));
 sg13g2_mux2_1 _16888_ (.A0(_01444_),
    .A1(_01480_),
    .S(net7783),
    .X(_03308_));
 sg13g2_nor3_1 _16889_ (.A(net7572),
    .B(net7571),
    .C(_03308_),
    .Y(_03309_));
 sg13g2_nor4_1 _16890_ (.A(_03303_),
    .B(_03305_),
    .C(_03307_),
    .D(_03309_),
    .Y(_03310_));
 sg13g2_mux4_1 _16891_ (.S0(net7786),
    .A0(_01233_),
    .A1(_01268_),
    .A2(_01304_),
    .A3(_01339_),
    .S1(net7727),
    .X(_03311_));
 sg13g2_nor2_1 _16892_ (.A(net7588),
    .B(_03311_),
    .Y(_03312_));
 sg13g2_mux4_1 _16893_ (.S0(net7786),
    .A0(_01092_),
    .A1(_01128_),
    .A2(_01163_),
    .A3(_01198_),
    .S1(net7727),
    .X(_03313_));
 sg13g2_inv_1 _16894_ (.Y(_03314_),
    .A(_03313_));
 sg13g2_a21oi_1 _16895_ (.A1(_08387_),
    .A2(_03314_),
    .Y(_03315_),
    .B1(_03312_));
 sg13g2_mux4_1 _16896_ (.S0(net7783),
    .A0(_00815_),
    .A1(_00847_),
    .A2(_00881_),
    .A3(_00916_),
    .S1(net7745),
    .X(_03316_));
 sg13g2_nand2_1 _16897_ (.Y(_03317_),
    .A(net7602),
    .B(_03316_));
 sg13g2_mux2_1 _16898_ (.A0(_00655_),
    .A1(_00783_),
    .S(net7711),
    .X(_03318_));
 sg13g2_a22oi_1 _16899_ (.Y(_03319_),
    .B1(_03318_),
    .B2(net7435),
    .A2(_10449_),
    .A1(_01511_));
 sg13g2_a21oi_1 _16900_ (.A1(_01159_),
    .A2(net7423),
    .Y(_03320_),
    .B1(net7691));
 sg13g2_mux4_1 _16901_ (.S0(net7784),
    .A0(_00952_),
    .A1(_00987_),
    .A2(_01022_),
    .A3(_01057_),
    .S1(net7745),
    .X(_03321_));
 sg13g2_mux2_1 _16902_ (.A0(_00687_),
    .A1(_00719_),
    .S(net7799),
    .X(_03322_));
 sg13g2_a22oi_1 _16903_ (.Y(_03323_),
    .B1(_03322_),
    .B2(net7516),
    .A2(net7595),
    .A1(_00751_));
 sg13g2_o21ai_1 _16904_ (.B1(net7711),
    .Y(_03324_),
    .A1(net7533),
    .A2(_03321_));
 sg13g2_a21o_1 _16905_ (.A2(_03323_),
    .A1(net7533),
    .B1(_03324_),
    .X(_03325_));
 sg13g2_nand4_1 _16906_ (.B(_03319_),
    .C(_03320_),
    .A(_03317_),
    .Y(_03326_),
    .D(_03325_));
 sg13g2_and3_1 _16907_ (.X(_03327_),
    .A(_03310_),
    .B(_03315_),
    .C(_03326_));
 sg13g2_a221oi_1 _16908_ (.B2(_08639_),
    .C1(net7073),
    .B1(_03327_),
    .A1(net7682),
    .Y(_03328_),
    .A2(net7268));
 sg13g2_nor2b_1 _16909_ (.A(net6979),
    .B_N(_03328_),
    .Y(_03329_));
 sg13g2_nand2b_1 _16910_ (.Y(_03330_),
    .B(_01585_),
    .A_N(net7874));
 sg13g2_nand2_1 _16911_ (.Y(_03331_),
    .A(net7874),
    .B(_00628_));
 sg13g2_nand3_1 _16912_ (.B(_03330_),
    .C(_03331_),
    .A(net7450),
    .Y(_03332_));
 sg13g2_nand2_1 _16913_ (.Y(_03333_),
    .A(net7874),
    .B(_01550_));
 sg13g2_nand2b_1 _16914_ (.Y(_03334_),
    .B(_01515_),
    .A_N(net7874));
 sg13g2_nand4_1 _16915_ (.B(net7493),
    .C(_03333_),
    .A(net7514),
    .Y(_03335_),
    .D(_03334_));
 sg13g2_nand2_1 _16916_ (.Y(_03336_),
    .A(net7873),
    .B(_01057_));
 sg13g2_nand2b_1 _16917_ (.Y(_03337_),
    .B(_01022_),
    .A_N(net7873));
 sg13g2_nand4_1 _16918_ (.B(net7526),
    .C(_03336_),
    .A(net7543),
    .Y(_03338_),
    .D(_03337_));
 sg13g2_nand2_1 _16919_ (.Y(_03339_),
    .A(net7873),
    .B(_00987_));
 sg13g2_nand2b_1 _16920_ (.Y(_03340_),
    .B(_00952_),
    .A_N(net7873));
 sg13g2_nand4_1 _16921_ (.B(net7514),
    .C(_03339_),
    .A(net7543),
    .Y(_03341_),
    .D(_03340_));
 sg13g2_nand2_1 _16922_ (.Y(_03342_),
    .A(net7873),
    .B(_00847_));
 sg13g2_nand2b_1 _16923_ (.Y(_03343_),
    .B(_00815_),
    .A_N(net7873));
 sg13g2_nand4_1 _16924_ (.B(net7472),
    .C(_03342_),
    .A(net7543),
    .Y(_03344_),
    .D(_03343_));
 sg13g2_nand2_1 _16925_ (.Y(_03345_),
    .A(net7873),
    .B(_00916_));
 sg13g2_nand2b_1 _16926_ (.Y(_03346_),
    .B(_00881_),
    .A_N(net7873));
 sg13g2_nand4_1 _16927_ (.B(net7463),
    .C(_03345_),
    .A(net7543),
    .Y(_03347_),
    .D(_03346_));
 sg13g2_nand2_1 _16928_ (.Y(_03348_),
    .A(net7874),
    .B(_01409_));
 sg13g2_nand2b_1 _16929_ (.Y(_03349_),
    .B(_01374_),
    .A_N(net7874));
 sg13g2_nand4_1 _16930_ (.B(net7472),
    .C(_03348_),
    .A(net7493),
    .Y(_03350_),
    .D(_03349_));
 sg13g2_nand2_1 _16931_ (.Y(_03351_),
    .A(net7874),
    .B(_01480_));
 sg13g2_nand2b_1 _16932_ (.Y(_03352_),
    .B(_01444_),
    .A_N(net7874));
 sg13g2_nand4_1 _16933_ (.B(net7463),
    .C(_03351_),
    .A(net7493),
    .Y(_03353_),
    .D(_03352_));
 sg13g2_nand4_1 _16934_ (.B(_03344_),
    .C(_03350_),
    .A(_03338_),
    .Y(_03354_),
    .D(_03353_));
 sg13g2_nand4_1 _16935_ (.B(_03335_),
    .C(_03341_),
    .A(_03332_),
    .Y(_03355_),
    .D(_03347_));
 sg13g2_mux2_1 _16936_ (.A0(_01511_),
    .A1(_00655_),
    .S(net7893),
    .X(_03356_));
 sg13g2_and2_1 _16937_ (.A(net7893),
    .B(_01159_),
    .X(_03357_));
 sg13g2_mux2_1 _16938_ (.A0(_00687_),
    .A1(_00719_),
    .S(net7893),
    .X(_03358_));
 sg13g2_mux2_1 _16939_ (.A0(_00751_),
    .A1(_00783_),
    .S(net7893),
    .X(_03359_));
 sg13g2_mux4_1 _16940_ (.S0(net7815),
    .A0(_03357_),
    .A1(_03358_),
    .A2(_03356_),
    .A3(_03359_),
    .S1(net7833),
    .X(_03360_));
 sg13g2_nor2_1 _16941_ (.A(net7529),
    .B(_03360_),
    .Y(_03361_));
 sg13g2_mux4_1 _16942_ (.S0(net7872),
    .A0(_01092_),
    .A1(_01128_),
    .A2(_01163_),
    .A3(_01198_),
    .S1(net7833),
    .X(_03362_));
 sg13g2_mux4_1 _16943_ (.S0(net7872),
    .A0(_01233_),
    .A1(_01268_),
    .A2(_01304_),
    .A3(_01339_),
    .S1(net7833),
    .X(_03363_));
 sg13g2_or2_1 _16944_ (.X(_03364_),
    .B(_03363_),
    .A(net7443));
 sg13g2_o21ai_1 _16945_ (.B1(_03364_),
    .Y(_03365_),
    .A1(net7421),
    .A2(_03362_));
 sg13g2_nor4_1 _16946_ (.A(_03354_),
    .B(_03355_),
    .C(_03361_),
    .D(_03365_),
    .Y(_03366_));
 sg13g2_or4_1 _16947_ (.A(_03354_),
    .B(_03355_),
    .C(_03361_),
    .D(_03365_),
    .X(_03367_));
 sg13g2_nand2b_1 _16948_ (.Y(_03368_),
    .B(net7999),
    .A_N(_01662_));
 sg13g2_o21ai_1 _16949_ (.B1(_03368_),
    .Y(_03369_),
    .A1(_01626_),
    .A2(net7478));
 sg13g2_a21oi_1 _16950_ (.A1(net8004),
    .A2(_03367_),
    .Y(_03370_),
    .B1(_03369_));
 sg13g2_o21ai_1 _16951_ (.B1(_03370_),
    .Y(_03371_),
    .A1(_09277_),
    .A2(_03327_));
 sg13g2_a21oi_1 _16952_ (.A1(net7377),
    .A2(_03371_),
    .Y(_03372_),
    .B1(_03329_));
 sg13g2_o21ai_1 _16953_ (.B1(_03372_),
    .Y(_03373_),
    .A1(_08254_),
    .A2(_03328_));
 sg13g2_mux2_1 _16954_ (.A0(_01375_),
    .A1(_01410_),
    .S(net7802),
    .X(_03374_));
 sg13g2_nor3_1 _16955_ (.A(net7572),
    .B(net7558),
    .C(_03374_),
    .Y(_03375_));
 sg13g2_mux2_1 _16956_ (.A0(_01516_),
    .A1(_01551_),
    .S(net7802),
    .X(_03376_));
 sg13g2_nor3_1 _16957_ (.A(net7572),
    .B(net7562),
    .C(_03376_),
    .Y(_03377_));
 sg13g2_mux2_1 _16958_ (.A0(_01446_),
    .A1(_01481_),
    .S(net7802),
    .X(_03378_));
 sg13g2_nor3_1 _16959_ (.A(net7572),
    .B(net7571),
    .C(_03378_),
    .Y(_03379_));
 sg13g2_mux2_1 _16960_ (.A0(_01586_),
    .A1(_00630_),
    .S(net7799),
    .X(_03380_));
 sg13g2_nor2_1 _16961_ (.A(net7555),
    .B(_03380_),
    .Y(_03381_));
 sg13g2_or4_1 _16962_ (.A(_03375_),
    .B(_03377_),
    .C(_03379_),
    .D(_03381_),
    .X(_03382_));
 sg13g2_mux4_1 _16963_ (.S0(net7801),
    .A0(_01234_),
    .A1(_01270_),
    .A2(_01305_),
    .A3(_01340_),
    .S1(net7746),
    .X(_03383_));
 sg13g2_mux4_1 _16964_ (.S0(net7802),
    .A0(_01094_),
    .A1(_01129_),
    .A2(_01164_),
    .A3(_01199_),
    .S1(net7741),
    .X(_03384_));
 sg13g2_nand2b_1 _16965_ (.Y(_03385_),
    .B(net7709),
    .A_N(_03383_));
 sg13g2_o21ai_1 _16966_ (.B1(_03385_),
    .Y(_03386_),
    .A1(net7710),
    .A2(_03384_));
 sg13g2_a21oi_1 _16967_ (.A1(net7591),
    .A2(_03386_),
    .Y(_03387_),
    .B1(_03382_));
 sg13g2_mux4_1 _16968_ (.S0(net7794),
    .A0(_00816_),
    .A1(_00848_),
    .A2(_00882_),
    .A3(_00918_),
    .S1(net7741),
    .X(_03388_));
 sg13g2_and2_1 _16969_ (.A(net7604),
    .B(_03388_),
    .X(_03389_));
 sg13g2_nand2_1 _16970_ (.Y(_03390_),
    .A(net7707),
    .B(_00784_));
 sg13g2_nand2b_1 _16971_ (.Y(_03391_),
    .B(_00656_),
    .A_N(net7707));
 sg13g2_a21oi_1 _16972_ (.A1(_03390_),
    .A2(_03391_),
    .Y(_03392_),
    .B1(net7600));
 sg13g2_nand3b_1 _16973_ (.B(net7794),
    .C(_01170_),
    .Y(_03393_),
    .A_N(net7738));
 sg13g2_nand3b_1 _16974_ (.B(_01522_),
    .C(net7738),
    .Y(_03394_),
    .A_N(net7794));
 sg13g2_a21oi_1 _16975_ (.A1(_03393_),
    .A2(_03394_),
    .Y(_03395_),
    .B1(net7598));
 sg13g2_nor4_1 _16976_ (.A(net7690),
    .B(_03389_),
    .C(_03392_),
    .D(_03395_),
    .Y(_03396_));
 sg13g2_mux4_1 _16977_ (.S0(net7792),
    .A0(_00953_),
    .A1(_00988_),
    .A2(_01023_),
    .A3(_01058_),
    .S1(net7741),
    .X(_03397_));
 sg13g2_nand2b_1 _16978_ (.Y(_03398_),
    .B(net7694),
    .A_N(_03397_));
 sg13g2_mux2_1 _16979_ (.A0(_00688_),
    .A1(_00720_),
    .S(net7796),
    .X(_03399_));
 sg13g2_a221oi_1 _16980_ (.B2(net7516),
    .C1(net7694),
    .B1(_03399_),
    .A1(_00752_),
    .Y(_03400_),
    .A2(net7595));
 sg13g2_nand3b_1 _16981_ (.B(net7707),
    .C(_03398_),
    .Y(_03401_),
    .A_N(_03400_));
 sg13g2_nand2_1 _16982_ (.Y(_03402_),
    .A(_03396_),
    .B(_03401_));
 sg13g2_a221oi_1 _16983_ (.B2(_03401_),
    .C1(_03382_),
    .B1(_03396_),
    .A1(net7591),
    .Y(_03403_),
    .A2(_03386_));
 sg13g2_nand2_1 _16984_ (.Y(_03404_),
    .A(_03387_),
    .B(_03402_));
 sg13g2_a21oi_1 _16985_ (.A1(net7681),
    .A2(net7268),
    .Y(_03405_),
    .B1(_02852_));
 sg13g2_o21ai_1 _16986_ (.B1(_03405_),
    .Y(_03406_),
    .A1(net7291),
    .A2(_03404_));
 sg13g2_mux2_1 _16987_ (.A0(_01586_),
    .A1(_00630_),
    .S(net7886),
    .X(_03407_));
 sg13g2_nor2_1 _16988_ (.A(net7449),
    .B(_03407_),
    .Y(_03408_));
 sg13g2_mux2_1 _16989_ (.A0(_01516_),
    .A1(_01551_),
    .S(net7890),
    .X(_03409_));
 sg13g2_nor3_1 _16990_ (.A(net7509),
    .B(net7491),
    .C(_03409_),
    .Y(_03410_));
 sg13g2_mux2_1 _16991_ (.A0(_00816_),
    .A1(_00848_),
    .S(net7883),
    .X(_03411_));
 sg13g2_nor3_1 _16992_ (.A(net7535),
    .B(net7465),
    .C(_03411_),
    .Y(_03412_));
 sg13g2_mux2_1 _16993_ (.A0(_00882_),
    .A1(_00918_),
    .S(net7883),
    .X(_03413_));
 sg13g2_nor3_1 _16994_ (.A(net7535),
    .B(net7461),
    .C(_03413_),
    .Y(_03414_));
 sg13g2_nor4_1 _16995_ (.A(_03408_),
    .B(_03410_),
    .C(_03412_),
    .D(_03414_),
    .Y(_03415_));
 sg13g2_mux2_1 _16996_ (.A0(_01023_),
    .A1(_01058_),
    .S(net7884),
    .X(_03416_));
 sg13g2_nor3_1 _16997_ (.A(net7535),
    .B(net7521),
    .C(_03416_),
    .Y(_03417_));
 sg13g2_mux2_1 _16998_ (.A0(_00953_),
    .A1(_00988_),
    .S(net7884),
    .X(_03418_));
 sg13g2_nor3_1 _16999_ (.A(net7535),
    .B(net7509),
    .C(_03418_),
    .Y(_03419_));
 sg13g2_mux2_1 _17000_ (.A0(_01375_),
    .A1(_01410_),
    .S(net7890),
    .X(_03420_));
 sg13g2_nor3_1 _17001_ (.A(net7491),
    .B(net7465),
    .C(_03420_),
    .Y(_03421_));
 sg13g2_mux2_1 _17002_ (.A0(_01446_),
    .A1(_01481_),
    .S(net7890),
    .X(_03422_));
 sg13g2_nor3_1 _17003_ (.A(net7491),
    .B(net7461),
    .C(_03422_),
    .Y(_03423_));
 sg13g2_nor4_1 _17004_ (.A(_03417_),
    .B(_03419_),
    .C(_03421_),
    .D(_03423_),
    .Y(_03424_));
 sg13g2_mux2_1 _17005_ (.A0(_01522_),
    .A1(_00656_),
    .S(net7847),
    .X(_03425_));
 sg13g2_and2_1 _17006_ (.A(net7847),
    .B(_01170_),
    .X(_03426_));
 sg13g2_mux2_1 _17007_ (.A0(_00688_),
    .A1(_00720_),
    .S(net7850),
    .X(_03427_));
 sg13g2_mux2_1 _17008_ (.A0(_00752_),
    .A1(_00784_),
    .S(net7850),
    .X(_03428_));
 sg13g2_mux4_1 _17009_ (.S0(net7811),
    .A0(_03426_),
    .A1(_03427_),
    .A2(_03425_),
    .A3(_03428_),
    .S1(net7826),
    .X(_03429_));
 sg13g2_or2_1 _17010_ (.X(_03430_),
    .B(_03429_),
    .A(net7529));
 sg13g2_mux4_1 _17011_ (.S0(net7886),
    .A0(_01094_),
    .A1(_01129_),
    .A2(_01164_),
    .A3(_01199_),
    .S1(net7824),
    .X(_03431_));
 sg13g2_nor3_1 _17012_ (.A(net7815),
    .B(_09073_),
    .C(_03431_),
    .Y(_03432_));
 sg13g2_mux4_1 _17013_ (.S0(net7888),
    .A0(_01234_),
    .A1(_01270_),
    .A2(_01305_),
    .A3(_01340_),
    .S1(net7824),
    .X(_03433_));
 sg13g2_nor2_1 _17014_ (.A(net7443),
    .B(_03433_),
    .Y(_03434_));
 sg13g2_nor2_1 _17015_ (.A(_03432_),
    .B(_03434_),
    .Y(_03435_));
 sg13g2_and4_1 _17016_ (.A(_03415_),
    .B(_03424_),
    .C(_03430_),
    .D(_03435_),
    .X(_03436_));
 sg13g2_nand4_1 _17017_ (.B(_03424_),
    .C(_03430_),
    .A(_03415_),
    .Y(_03437_),
    .D(_03435_));
 sg13g2_nand2b_1 _17018_ (.Y(_03438_),
    .B(net7999),
    .A_N(_01663_));
 sg13g2_o21ai_1 _17019_ (.B1(_03438_),
    .Y(_03439_),
    .A1(_01627_),
    .A2(net7478));
 sg13g2_a221oi_1 _17020_ (.B2(net8004),
    .C1(_03439_),
    .B1(net7331),
    .A1(net7352),
    .Y(_03440_),
    .A2(net7260));
 sg13g2_mux2_1 _17021_ (.A0(net6981),
    .A1(_08254_),
    .S(_03406_),
    .X(_03441_));
 sg13g2_o21ai_1 _17022_ (.B1(_03441_),
    .Y(_03442_),
    .A1(net7375),
    .A2(_03440_));
 sg13g2_mux2_1 _17023_ (.A0(_01376_),
    .A1(_01411_),
    .S(net7755),
    .X(_03443_));
 sg13g2_nor3_1 _17024_ (.A(net7581),
    .B(net7560),
    .C(_03443_),
    .Y(_03444_));
 sg13g2_mux2_1 _17025_ (.A0(_01517_),
    .A1(_01552_),
    .S(net7756),
    .X(_03445_));
 sg13g2_nor3_1 _17026_ (.A(net7581),
    .B(net7564),
    .C(_03445_),
    .Y(_03446_));
 sg13g2_mux2_1 _17027_ (.A0(_01447_),
    .A1(_01482_),
    .S(net7755),
    .X(_03447_));
 sg13g2_nor3_1 _17028_ (.A(net7581),
    .B(net7568),
    .C(_03447_),
    .Y(_03448_));
 sg13g2_mux2_1 _17029_ (.A0(_01587_),
    .A1(_00631_),
    .S(net7756),
    .X(_03449_));
 sg13g2_nor2_1 _17030_ (.A(net7552),
    .B(_03449_),
    .Y(_03450_));
 sg13g2_or4_1 _17031_ (.A(_03444_),
    .B(_03446_),
    .C(_03448_),
    .D(_03450_),
    .X(_03451_));
 sg13g2_mux4_1 _17032_ (.S0(net7750),
    .A0(_01235_),
    .A1(_01271_),
    .A2(_01306_),
    .A3(_01341_),
    .S1(net7718),
    .X(_03452_));
 sg13g2_mux4_1 _17033_ (.S0(net7749),
    .A0(_01095_),
    .A1(_01130_),
    .A2(_01165_),
    .A3(_01200_),
    .S1(net7721),
    .X(_03453_));
 sg13g2_nand2b_1 _17034_ (.Y(_03454_),
    .B(net7702),
    .A_N(_03452_));
 sg13g2_o21ai_1 _17035_ (.B1(_03454_),
    .Y(_03455_),
    .A1(net7702),
    .A2(_03453_));
 sg13g2_a21oi_1 _17036_ (.A1(net7589),
    .A2(_03455_),
    .Y(_03456_),
    .B1(_03451_));
 sg13g2_mux4_1 _17037_ (.S0(net7762),
    .A0(_00817_),
    .A1(_00849_),
    .A2(_00883_),
    .A3(_00919_),
    .S1(net7730),
    .X(_03457_));
 sg13g2_and2_1 _17038_ (.A(net7606),
    .B(_03457_),
    .X(_03458_));
 sg13g2_nand2_1 _17039_ (.Y(_03459_),
    .A(net7700),
    .B(_00785_));
 sg13g2_nand2b_1 _17040_ (.Y(_03460_),
    .B(_00657_),
    .A_N(net7700));
 sg13g2_a21oi_1 _17041_ (.A1(_03459_),
    .A2(_03460_),
    .Y(_03461_),
    .B1(net7601));
 sg13g2_nand3b_1 _17042_ (.B(net7760),
    .C(_01181_),
    .Y(_03462_),
    .A_N(net7733));
 sg13g2_nand3b_1 _17043_ (.B(_01533_),
    .C(net7733),
    .Y(_03463_),
    .A_N(net7760));
 sg13g2_a21oi_1 _17044_ (.A1(_03462_),
    .A2(_03463_),
    .Y(_03464_),
    .B1(_08306_));
 sg13g2_nor4_1 _17045_ (.A(net7689),
    .B(_03458_),
    .C(_03461_),
    .D(_03464_),
    .Y(_03465_));
 sg13g2_mux4_1 _17046_ (.S0(net7752),
    .A0(_00954_),
    .A1(_00989_),
    .A2(_01024_),
    .A3(_01059_),
    .S1(net7719),
    .X(_03466_));
 sg13g2_nand2b_1 _17047_ (.Y(_03467_),
    .B(net7692),
    .A_N(_03466_));
 sg13g2_mux2_1 _17048_ (.A0(_00689_),
    .A1(_00721_),
    .S(net7760),
    .X(_03468_));
 sg13g2_a221oi_1 _17049_ (.B2(_09011_),
    .C1(net7692),
    .B1(_03468_),
    .A1(_00753_),
    .Y(_03469_),
    .A2(net7593));
 sg13g2_nand3b_1 _17050_ (.B(net7701),
    .C(_03467_),
    .Y(_03470_),
    .A_N(_03469_));
 sg13g2_nand2_1 _17051_ (.Y(_03471_),
    .A(_03465_),
    .B(_03470_));
 sg13g2_a221oi_1 _17052_ (.B2(_03470_),
    .C1(_03451_),
    .B1(_03465_),
    .A1(net7589),
    .Y(_03472_),
    .A2(_03455_));
 sg13g2_nand2_1 _17053_ (.Y(_03473_),
    .A(_03456_),
    .B(_03471_));
 sg13g2_a221oi_1 _17054_ (.B2(_08639_),
    .C1(net7073),
    .B1(net7330),
    .A1(_01907_),
    .Y(_03474_),
    .A2(net7268));
 sg13g2_mux2_1 _17055_ (.A0(_01587_),
    .A1(_00631_),
    .S(net7904),
    .X(_03475_));
 sg13g2_nor2_1 _17056_ (.A(net7448),
    .B(_03475_),
    .Y(_03476_));
 sg13g2_mux2_1 _17057_ (.A0(_01517_),
    .A1(_01552_),
    .S(net7904),
    .X(_03477_));
 sg13g2_nor3_1 _17058_ (.A(net7508),
    .B(net7488),
    .C(_03477_),
    .Y(_03478_));
 sg13g2_mux2_1 _17059_ (.A0(_01024_),
    .A1(_01059_),
    .S(net7901),
    .X(_03479_));
 sg13g2_nor3_1 _17060_ (.A(net7537),
    .B(net7522),
    .C(_03479_),
    .Y(_03480_));
 sg13g2_mux2_1 _17061_ (.A0(_00954_),
    .A1(_00989_),
    .S(net7901),
    .X(_03481_));
 sg13g2_nor3_1 _17062_ (.A(net7537),
    .B(net7506),
    .C(_03481_),
    .Y(_03482_));
 sg13g2_nor4_1 _17063_ (.A(_03476_),
    .B(_03478_),
    .C(_03480_),
    .D(_03482_),
    .Y(_03483_));
 sg13g2_mux2_1 _17064_ (.A0(_00817_),
    .A1(_00849_),
    .S(net7907),
    .X(_03484_));
 sg13g2_nor3_1 _17065_ (.A(net7539),
    .B(net7469),
    .C(_03484_),
    .Y(_03485_));
 sg13g2_mux2_1 _17066_ (.A0(_00883_),
    .A1(_00919_),
    .S(net7907),
    .X(_03486_));
 sg13g2_nor3_1 _17067_ (.A(net7539),
    .B(net7458),
    .C(_03486_),
    .Y(_03487_));
 sg13g2_mux2_1 _17068_ (.A0(_01376_),
    .A1(_01411_),
    .S(net7903),
    .X(_03488_));
 sg13g2_nor3_1 _17069_ (.A(net7488),
    .B(net7469),
    .C(_03488_),
    .Y(_03489_));
 sg13g2_mux2_1 _17070_ (.A0(_01447_),
    .A1(_01482_),
    .S(net7903),
    .X(_03490_));
 sg13g2_nor3_1 _17071_ (.A(net7489),
    .B(net7459),
    .C(_03490_),
    .Y(_03491_));
 sg13g2_nor4_1 _17072_ (.A(_03485_),
    .B(_03487_),
    .C(_03489_),
    .D(_03491_),
    .Y(_03492_));
 sg13g2_mux2_1 _17073_ (.A0(_01533_),
    .A1(_00657_),
    .S(net7836),
    .X(_03493_));
 sg13g2_and2_1 _17074_ (.A(net7836),
    .B(_01181_),
    .X(_03494_));
 sg13g2_mux2_1 _17075_ (.A0(_00689_),
    .A1(_00721_),
    .S(net7838),
    .X(_03495_));
 sg13g2_mux2_1 _17076_ (.A0(_00753_),
    .A1(_00785_),
    .S(net7836),
    .X(_03496_));
 sg13g2_mux4_1 _17077_ (.S0(net7810),
    .A0(_03494_),
    .A1(_03495_),
    .A2(_03493_),
    .A3(_03496_),
    .S1(net7820),
    .X(_03497_));
 sg13g2_or2_1 _17078_ (.X(_03498_),
    .B(_03497_),
    .A(net7528));
 sg13g2_mux4_1 _17079_ (.S0(net7899),
    .A0(_01095_),
    .A1(_01130_),
    .A2(_01165_),
    .A3(_01200_),
    .S1(net7818),
    .X(_03499_));
 sg13g2_nor3_1 _17080_ (.A(net7809),
    .B(net7499),
    .C(_03499_),
    .Y(_03500_));
 sg13g2_mux4_1 _17081_ (.S0(net7899),
    .A0(_01235_),
    .A1(_01271_),
    .A2(_01306_),
    .A3(_01341_),
    .S1(net7819),
    .X(_03501_));
 sg13g2_nor2_1 _17082_ (.A(net7444),
    .B(_03501_),
    .Y(_03502_));
 sg13g2_nor2_1 _17083_ (.A(_03500_),
    .B(_03502_),
    .Y(_03503_));
 sg13g2_and4_1 _17084_ (.A(_03483_),
    .B(_03492_),
    .C(_03498_),
    .D(_03503_),
    .X(_03504_));
 sg13g2_nand4_1 _17085_ (.B(_03492_),
    .C(_03498_),
    .A(_03483_),
    .Y(_03505_),
    .D(_03503_));
 sg13g2_nand2b_1 _17086_ (.Y(_03506_),
    .B(net7993),
    .A_N(_01664_));
 sg13g2_o21ai_1 _17087_ (.B1(_03506_),
    .Y(_03507_),
    .A1(_01628_),
    .A2(net7481));
 sg13g2_a221oi_1 _17088_ (.B2(net8008),
    .C1(_03507_),
    .B1(net7329),
    .A1(net7353),
    .Y(_03508_),
    .A2(_03473_));
 sg13g2_nand2_1 _17089_ (.Y(_03509_),
    .A(net6978),
    .B(_03474_));
 sg13g2_o21ai_1 _17090_ (.B1(_03509_),
    .Y(_03510_),
    .A1(net6918),
    .A2(_03474_));
 sg13g2_o21ai_1 _17091_ (.B1(_03510_),
    .Y(_03511_),
    .A1(net7374),
    .A2(_03508_));
 sg13g2_mux2_1 _17092_ (.A0(_01589_),
    .A1(_00632_),
    .S(net7800),
    .X(_03512_));
 sg13g2_nor2_1 _17093_ (.A(net7550),
    .B(_03512_),
    .Y(_03513_));
 sg13g2_mux2_1 _17094_ (.A0(_01377_),
    .A1(_01413_),
    .S(net7800),
    .X(_03514_));
 sg13g2_nor3_1 _17095_ (.A(net7575),
    .B(net7557),
    .C(_03514_),
    .Y(_03515_));
 sg13g2_mux2_1 _17096_ (.A0(_01448_),
    .A1(_01483_),
    .S(net7800),
    .X(_03516_));
 sg13g2_nor3_1 _17097_ (.A(net7575),
    .B(net7570),
    .C(_03516_),
    .Y(_03517_));
 sg13g2_mux2_1 _17098_ (.A0(_01518_),
    .A1(_01553_),
    .S(net7800),
    .X(_03518_));
 sg13g2_nor3_1 _17099_ (.A(net7575),
    .B(net7566),
    .C(_03518_),
    .Y(_03519_));
 sg13g2_nor4_1 _17100_ (.A(_03513_),
    .B(_03515_),
    .C(_03517_),
    .D(_03519_),
    .Y(_03520_));
 sg13g2_mux4_1 _17101_ (.S0(net7785),
    .A0(_01237_),
    .A1(_01272_),
    .A2(_01307_),
    .A3(_01342_),
    .S1(net7743),
    .X(_03521_));
 sg13g2_nor2_1 _17102_ (.A(net7587),
    .B(_03521_),
    .Y(_03522_));
 sg13g2_mux4_1 _17103_ (.S0(net7785),
    .A0(_01096_),
    .A1(_01131_),
    .A2(_01166_),
    .A3(_01201_),
    .S1(net7742),
    .X(_03523_));
 sg13g2_inv_1 _17104_ (.Y(_03524_),
    .A(_03523_));
 sg13g2_a21oi_1 _17105_ (.A1(net7434),
    .A2(_03524_),
    .Y(_03525_),
    .B1(_03522_));
 sg13g2_mux4_1 _17106_ (.S0(net7798),
    .A0(_00818_),
    .A1(_00850_),
    .A2(_00885_),
    .A3(_00920_),
    .S1(net7740),
    .X(_03526_));
 sg13g2_nand2_1 _17107_ (.Y(_03527_),
    .A(net7603),
    .B(_03526_));
 sg13g2_mux2_1 _17108_ (.A0(_00658_),
    .A1(_00786_),
    .S(net7704),
    .X(_03528_));
 sg13g2_a22oi_1 _17109_ (.Y(_03529_),
    .B1(_03528_),
    .B2(net7435),
    .A2(net7423),
    .A1(_01192_));
 sg13g2_a21oi_1 _17110_ (.A1(_01544_),
    .A2(_10449_),
    .Y(_03530_),
    .B1(net7691));
 sg13g2_mux4_1 _17111_ (.S0(net7800),
    .A0(_00955_),
    .A1(_00990_),
    .A2(_01025_),
    .A3(_01061_),
    .S1(net7740),
    .X(_03531_));
 sg13g2_nand2b_1 _17112_ (.Y(_03532_),
    .B(net7694),
    .A_N(_03531_));
 sg13g2_mux2_1 _17113_ (.A0(_00690_),
    .A1(_00722_),
    .S(net7800),
    .X(_03533_));
 sg13g2_a221oi_1 _17114_ (.B2(net7517),
    .C1(net7694),
    .B1(_03533_),
    .A1(_00754_),
    .Y(_03534_),
    .A2(net7596));
 sg13g2_nand3b_1 _17115_ (.B(net7704),
    .C(_03532_),
    .Y(_03535_),
    .A_N(_03534_));
 sg13g2_nand4_1 _17116_ (.B(_03529_),
    .C(_03530_),
    .A(_03527_),
    .Y(_03536_),
    .D(_03535_));
 sg13g2_inv_1 _17117_ (.Y(_03537_),
    .A(net7259));
 sg13g2_nand3_1 _17118_ (.B(_03525_),
    .C(_03536_),
    .A(_03520_),
    .Y(_03538_));
 sg13g2_a221oi_1 _17119_ (.B2(net7292),
    .C1(net7073),
    .B1(_03537_),
    .A1(_01909_),
    .Y(_03539_),
    .A2(net7268));
 sg13g2_mux2_1 _17120_ (.A0(_01544_),
    .A1(_00658_),
    .S(net7881),
    .X(_03540_));
 sg13g2_a22oi_1 _17121_ (.Y(_03541_),
    .B1(_03540_),
    .B2(net7824),
    .A2(net7527),
    .A1(_01192_));
 sg13g2_nand2b_1 _17122_ (.Y(_03542_),
    .B(net7881),
    .A_N(_00722_));
 sg13g2_o21ai_1 _17123_ (.B1(_03542_),
    .Y(_03543_),
    .A1(net7881),
    .A2(_00690_));
 sg13g2_mux2_1 _17124_ (.A0(_00754_),
    .A1(_00786_),
    .S(net7881),
    .X(_03544_));
 sg13g2_o21ai_1 _17125_ (.B1(net7530),
    .Y(_03545_),
    .A1(net7521),
    .A2(_03544_));
 sg13g2_a221oi_1 _17126_ (.B2(_09026_),
    .C1(_03545_),
    .B1(_03543_),
    .A1(net7483),
    .Y(_03546_),
    .A2(_03541_));
 sg13g2_mux2_1 _17127_ (.A0(_01307_),
    .A1(_01342_),
    .S(net7893),
    .X(_03547_));
 sg13g2_nor2_1 _17128_ (.A(net7521),
    .B(_03547_),
    .Y(_03548_));
 sg13g2_mux2_1 _17129_ (.A0(_01096_),
    .A1(_01131_),
    .S(net7894),
    .X(_03549_));
 sg13g2_nor2_1 _17130_ (.A(net7465),
    .B(_03549_),
    .Y(_03550_));
 sg13g2_mux2_1 _17131_ (.A0(_01166_),
    .A1(_01201_),
    .S(net7882),
    .X(_03551_));
 sg13g2_nor2_1 _17132_ (.A(net7461),
    .B(_03551_),
    .Y(_03552_));
 sg13g2_mux2_1 _17133_ (.A0(_01237_),
    .A1(_01272_),
    .S(net7894),
    .X(_03553_));
 sg13g2_o21ai_1 _17134_ (.B1(net7501),
    .Y(_03554_),
    .A1(net7509),
    .A2(_03553_));
 sg13g2_nor4_1 _17135_ (.A(_03548_),
    .B(_03550_),
    .C(_03552_),
    .D(_03554_),
    .Y(_03555_));
 sg13g2_mux2_1 _17136_ (.A0(_01589_),
    .A1(_00632_),
    .S(net7882),
    .X(_03556_));
 sg13g2_nand2_1 _17137_ (.Y(_03557_),
    .A(net7450),
    .B(_03556_));
 sg13g2_mux2_1 _17138_ (.A0(_01518_),
    .A1(_01553_),
    .S(net7881),
    .X(_03558_));
 sg13g2_nand3_1 _17139_ (.B(net7496),
    .C(_03558_),
    .A(_09026_),
    .Y(_03559_));
 sg13g2_mux2_1 _17140_ (.A0(_01448_),
    .A1(_01483_),
    .S(net7882),
    .X(_03560_));
 sg13g2_nand3_1 _17141_ (.B(net7462),
    .C(_03560_),
    .A(net7496),
    .Y(_03561_));
 sg13g2_mux2_1 _17142_ (.A0(_01377_),
    .A1(_01413_),
    .S(net7882),
    .X(_03562_));
 sg13g2_nand3_1 _17143_ (.B(net7471),
    .C(_03562_),
    .A(net7496),
    .Y(_03563_));
 sg13g2_mux2_1 _17144_ (.A0(_00885_),
    .A1(_00920_),
    .S(net7881),
    .X(_03564_));
 sg13g2_nand3_1 _17145_ (.B(net7462),
    .C(_03564_),
    .A(net7547),
    .Y(_03565_));
 sg13g2_mux2_1 _17146_ (.A0(_00818_),
    .A1(_00850_),
    .S(net7881),
    .X(_03566_));
 sg13g2_nand3_1 _17147_ (.B(net7471),
    .C(_03566_),
    .A(net7547),
    .Y(_03567_));
 sg13g2_mux2_1 _17148_ (.A0(_00955_),
    .A1(_00990_),
    .S(net7882),
    .X(_03568_));
 sg13g2_nand3_1 _17149_ (.B(_09026_),
    .C(_03568_),
    .A(net7547),
    .Y(_03569_));
 sg13g2_mux2_1 _17150_ (.A0(_01025_),
    .A1(_01061_),
    .S(net7881),
    .X(_03570_));
 sg13g2_nand3_1 _17151_ (.B(net7525),
    .C(_03570_),
    .A(net7547),
    .Y(_03571_));
 sg13g2_nand4_1 _17152_ (.B(_03561_),
    .C(_03563_),
    .A(_03557_),
    .Y(_03572_),
    .D(_03569_));
 sg13g2_nand4_1 _17153_ (.B(_03565_),
    .C(_03567_),
    .A(_03559_),
    .Y(_03573_),
    .D(_03571_));
 sg13g2_nor4_1 _17154_ (.A(_03546_),
    .B(_03555_),
    .C(_03572_),
    .D(_03573_),
    .Y(_03574_));
 sg13g2_or4_1 _17155_ (.A(_03546_),
    .B(_03555_),
    .C(_03572_),
    .D(_03573_),
    .X(_03575_));
 sg13g2_nand2b_1 _17156_ (.Y(_03576_),
    .B(net8002),
    .A_N(_01665_));
 sg13g2_o21ai_1 _17157_ (.B1(_03576_),
    .Y(_03577_),
    .A1(_01630_),
    .A2(net7481));
 sg13g2_a221oi_1 _17158_ (.B2(net8008),
    .C1(_03577_),
    .B1(net7328),
    .A1(net7353),
    .Y(_03578_),
    .A2(net7259));
 sg13g2_nand2_1 _17159_ (.Y(_03579_),
    .A(net6979),
    .B(_03539_));
 sg13g2_o21ai_1 _17160_ (.B1(_03579_),
    .Y(_03580_),
    .A1(net6919),
    .A2(_03539_));
 sg13g2_o21ai_1 _17161_ (.B1(_03580_),
    .Y(_03581_),
    .A1(net7374),
    .A2(_03578_));
 sg13g2_mux4_1 _17162_ (.S0(net7790),
    .A0(_00819_),
    .A1(_00851_),
    .A2(_00886_),
    .A3(_00921_),
    .S1(net7740),
    .X(_03582_));
 sg13g2_nand2_1 _17163_ (.Y(_03583_),
    .A(net7604),
    .B(_03582_));
 sg13g2_a21oi_1 _17164_ (.A1(_01203_),
    .A2(net7423),
    .Y(_03584_),
    .B1(net7691));
 sg13g2_mux2_1 _17165_ (.A0(_00659_),
    .A1(_00787_),
    .S(net7704),
    .X(_03585_));
 sg13g2_a22oi_1 _17166_ (.Y(_03586_),
    .B1(_03585_),
    .B2(_08288_),
    .A2(_10449_),
    .A1(_01555_));
 sg13g2_mux4_1 _17167_ (.S0(net7797),
    .A0(_00956_),
    .A1(_00991_),
    .A2(_01026_),
    .A3(_01062_),
    .S1(net7739),
    .X(_03587_));
 sg13g2_mux2_1 _17168_ (.A0(_00691_),
    .A1(_00723_),
    .S(net7804),
    .X(_03588_));
 sg13g2_a22oi_1 _17169_ (.Y(_03589_),
    .B1(_03588_),
    .B2(net7517),
    .A2(net7596),
    .A1(_00755_));
 sg13g2_o21ai_1 _17170_ (.B1(net7704),
    .Y(_03590_),
    .A1(net7531),
    .A2(_03587_));
 sg13g2_a21o_1 _17171_ (.A2(_03589_),
    .A1(net7531),
    .B1(_03590_),
    .X(_03591_));
 sg13g2_nand4_1 _17172_ (.B(_03584_),
    .C(_03586_),
    .A(_03583_),
    .Y(_03592_),
    .D(_03591_));
 sg13g2_mux2_1 _17173_ (.A0(_01590_),
    .A1(_00633_),
    .S(net7790),
    .X(_03593_));
 sg13g2_nor2_1 _17174_ (.A(net7550),
    .B(_03593_),
    .Y(_03594_));
 sg13g2_mux2_1 _17175_ (.A0(_01449_),
    .A1(_01484_),
    .S(net7790),
    .X(_03595_));
 sg13g2_nor3_1 _17176_ (.A(net7575),
    .B(net7570),
    .C(_03595_),
    .Y(_03596_));
 sg13g2_mux2_1 _17177_ (.A0(_01519_),
    .A1(_01554_),
    .S(net7790),
    .X(_03597_));
 sg13g2_nor3_1 _17178_ (.A(net7575),
    .B(net7566),
    .C(_03597_),
    .Y(_03598_));
 sg13g2_mux2_1 _17179_ (.A0(_01378_),
    .A1(_01414_),
    .S(net7790),
    .X(_03599_));
 sg13g2_nor3_1 _17180_ (.A(net7575),
    .B(net7557),
    .C(_03599_),
    .Y(_03600_));
 sg13g2_nor4_1 _17181_ (.A(_03594_),
    .B(_03596_),
    .C(_03598_),
    .D(_03600_),
    .Y(_03601_));
 sg13g2_mux4_1 _17182_ (.S0(net7790),
    .A0(_01097_),
    .A1(_01132_),
    .A2(_01167_),
    .A3(_01202_),
    .S1(net7737),
    .X(_03602_));
 sg13g2_inv_1 _17183_ (.Y(_03603_),
    .A(_03602_));
 sg13g2_mux4_1 _17184_ (.S0(net7790),
    .A0(_01238_),
    .A1(_01273_),
    .A2(_01308_),
    .A3(_01343_),
    .S1(net7737),
    .X(_03604_));
 sg13g2_nor2_1 _17185_ (.A(net7587),
    .B(_03604_),
    .Y(_03605_));
 sg13g2_a21oi_1 _17186_ (.A1(net7434),
    .A2(_03603_),
    .Y(_03606_),
    .B1(_03605_));
 sg13g2_and2_1 _17187_ (.A(_03601_),
    .B(_03606_),
    .X(_03607_));
 sg13g2_nand2_1 _17188_ (.Y(_03608_),
    .A(_03592_),
    .B(_03607_));
 sg13g2_o21ai_1 _17189_ (.B1(_08819_),
    .Y(_03609_),
    .A1(_08777_),
    .A2(_08797_));
 sg13g2_nand2_1 _17190_ (.Y(_03610_),
    .A(net7677),
    .B(_03609_));
 sg13g2_mux2_1 _17191_ (.A0(_03608_),
    .A1(_03610_),
    .S(net7291),
    .X(_03611_));
 sg13g2_nand2b_1 _17192_ (.Y(_03612_),
    .B(net7999),
    .A_N(net7977));
 sg13g2_o21ai_1 _17193_ (.B1(_03612_),
    .Y(_03613_),
    .A1(_01631_),
    .A2(net7481));
 sg13g2_mux4_1 _17194_ (.S0(net7855),
    .A0(_01238_),
    .A1(_01273_),
    .A2(_01308_),
    .A3(_01343_),
    .S1(net7826),
    .X(_03614_));
 sg13g2_mux4_1 _17195_ (.S0(net7855),
    .A0(_01097_),
    .A1(_01132_),
    .A2(_01167_),
    .A3(_01202_),
    .S1(net7826),
    .X(_03615_));
 sg13g2_mux2_1 _17196_ (.A0(_03614_),
    .A1(_03615_),
    .S(net7483),
    .X(_03616_));
 sg13g2_mux4_1 _17197_ (.S0(net7852),
    .A0(_01378_),
    .A1(_01414_),
    .A2(_01449_),
    .A3(_01484_),
    .S1(net7826),
    .X(_03617_));
 sg13g2_mux4_1 _17198_ (.S0(net7855),
    .A0(_01519_),
    .A1(_01554_),
    .A2(_01590_),
    .A3(_00633_),
    .S1(net7827),
    .X(_03618_));
 sg13g2_mux4_1 _17199_ (.S0(net7854),
    .A0(_00819_),
    .A1(_00851_),
    .A2(_00886_),
    .A3(_00921_),
    .S1(net7827),
    .X(_03619_));
 sg13g2_mux4_1 _17200_ (.S0(net7852),
    .A0(_00956_),
    .A1(_00991_),
    .A2(_01026_),
    .A3(_01062_),
    .S1(net7826),
    .X(_03620_));
 sg13g2_mux2_1 _17201_ (.A0(_00691_),
    .A1(_00723_),
    .S(net7854),
    .X(_03621_));
 sg13g2_mux2_1 _17202_ (.A0(_00755_),
    .A1(_00787_),
    .S(net7854),
    .X(_03622_));
 sg13g2_mux2_1 _17203_ (.A0(_01555_),
    .A1(_00659_),
    .S(net7854),
    .X(_03623_));
 sg13g2_and2_1 _17204_ (.A(net7854),
    .B(_01203_),
    .X(_03624_));
 sg13g2_mux4_1 _17205_ (.S0(net7825),
    .A0(_03621_),
    .A1(_03622_),
    .A2(_03624_),
    .A3(_03623_),
    .S1(net7483),
    .X(_03625_));
 sg13g2_mux2_1 _17206_ (.A0(_03617_),
    .A1(_03618_),
    .S(net7811),
    .X(_03626_));
 sg13g2_mux2_1 _17207_ (.A0(_03619_),
    .A1(_03620_),
    .S(net7811),
    .X(_03627_));
 sg13g2_inv_1 _17208_ (.Y(_03628_),
    .A(_03629_));
 sg13g2_mux4_1 _17209_ (.S0(net7807),
    .A0(_03625_),
    .A1(_03627_),
    .A2(_03616_),
    .A3(_03626_),
    .S1(net7805),
    .X(_03629_));
 sg13g2_a221oi_1 _17210_ (.B2(_00541_),
    .C1(_03613_),
    .B1(_03628_),
    .A1(_09275_),
    .Y(_03630_),
    .A2(_03608_));
 sg13g2_mux2_1 _17211_ (.A0(_08254_),
    .A1(_08228_),
    .S(_03611_),
    .X(_03631_));
 sg13g2_o21ai_1 _17212_ (.B1(_03631_),
    .Y(_03632_),
    .A1(net7374),
    .A2(_03630_));
 sg13g2_a21oi_1 _17213_ (.A1(_01914_),
    .A2(_07925_),
    .Y(_03633_),
    .B1(net7609));
 sg13g2_nand2b_1 _17214_ (.Y(_03634_),
    .B(net7674),
    .A_N(_03633_));
 sg13g2_nand3b_1 _17215_ (.B(net7676),
    .C(_01908_),
    .Y(_03635_),
    .A_N(_01912_));
 sg13g2_a21oi_1 _17216_ (.A1(_07954_),
    .A2(_03635_),
    .Y(_03636_),
    .B1(net7673));
 sg13g2_o21ai_1 _17217_ (.B1(_08533_),
    .Y(_03637_),
    .A1(net7609),
    .A2(_03636_));
 sg13g2_nor3_1 _17218_ (.A(_07590_),
    .B(_07948_),
    .C(_07954_),
    .Y(_03638_));
 sg13g2_and2_1 _17219_ (.A(net7920),
    .B(_03638_),
    .X(_03639_));
 sg13g2_or4_1 _17220_ (.A(_09244_),
    .B(_07590_),
    .C(_07948_),
    .D(_07954_),
    .X(_03640_));
 sg13g2_nand4_1 _17221_ (.B(_07895_),
    .C(net7432),
    .A(net7610),
    .Y(_03641_),
    .D(_03640_));
 sg13g2_a21oi_1 _17222_ (.A1(_03634_),
    .A2(_03637_),
    .Y(_03642_),
    .B1(_03641_));
 sg13g2_o21ai_1 _17223_ (.B1(_07590_),
    .Y(_03643_),
    .A1(net7607),
    .A2(_07872_));
 sg13g2_a21o_1 _17224_ (.A2(_03643_),
    .A1(_07881_),
    .B1(_07964_),
    .X(_03644_));
 sg13g2_a22oi_1 _17225_ (.Y(_03645_),
    .B1(_03644_),
    .B2(net7679),
    .A2(_08673_),
    .A1(_08622_));
 sg13g2_nand2_1 _17226_ (.Y(_03646_),
    .A(_03642_),
    .B(_03645_));
 sg13g2_and3_1 _17227_ (.X(_03647_),
    .A(net7838),
    .B(net7432),
    .C(_03639_));
 sg13g2_a21oi_1 _17228_ (.A1(_01949_),
    .A2(net7360),
    .Y(_03648_),
    .B1(_03647_));
 sg13g2_o21ai_1 _17229_ (.B1(_03648_),
    .Y(_03649_),
    .A1(_09252_),
    .A2(_03646_));
 sg13g2_nand2_1 _17230_ (.Y(_03650_),
    .A(net7364),
    .B(net7072));
 sg13g2_nand3_1 _17231_ (.B(net7384),
    .C(net7428),
    .A(_01632_),
    .Y(_03651_));
 sg13g2_nand2_1 _17232_ (.Y(_03652_),
    .A(_03650_),
    .B(_03651_));
 sg13g2_nor2b_1 _17233_ (.A(_03645_),
    .B_N(_03642_),
    .Y(_03653_));
 sg13g2_and3_1 _17234_ (.X(_03654_),
    .A(net7820),
    .B(net7432),
    .C(_03639_));
 sg13g2_a221oi_1 _17235_ (.B2(_01928_),
    .C1(_03654_),
    .B1(_03653_),
    .A1(_01960_),
    .Y(_03655_),
    .A2(net7362));
 sg13g2_nor2_1 _17236_ (.A(_10370_),
    .B(_03646_),
    .Y(_03656_));
 sg13g2_nor2b_1 _17237_ (.A(_03656_),
    .B_N(_03655_),
    .Y(_03657_));
 sg13g2_a21oi_1 _17238_ (.A1(_01633_),
    .A2(net7428),
    .Y(_03658_),
    .B1(net7376));
 sg13g2_a21oi_1 _17239_ (.A1(net7364),
    .A2(_03657_),
    .Y(_03659_),
    .B1(_03658_));
 sg13g2_nor3_1 _17240_ (.A(net7483),
    .B(net7360),
    .C(_03640_),
    .Y(_03660_));
 sg13g2_a221oi_1 _17241_ (.B2(_01939_),
    .C1(_03660_),
    .B1(_03653_),
    .A1(_01971_),
    .Y(_03661_),
    .A2(net7360));
 sg13g2_o21ai_1 _17242_ (.B1(_03661_),
    .Y(_03662_),
    .A1(net7283),
    .A2(_03646_));
 sg13g2_nand2_1 _17243_ (.Y(_03663_),
    .A(_08250_),
    .B(_03662_));
 sg13g2_nand3_1 _17244_ (.B(net7384),
    .C(net7428),
    .A(_01634_),
    .Y(_03664_));
 sg13g2_nand2_1 _17245_ (.Y(_03665_),
    .A(_03663_),
    .B(_03664_));
 sg13g2_and3_1 _17246_ (.X(_03666_),
    .A(net7807),
    .B(net7432),
    .C(_03639_));
 sg13g2_a221oi_1 _17247_ (.B2(_01942_),
    .C1(_03666_),
    .B1(_03653_),
    .A1(_01974_),
    .Y(_03667_),
    .A2(net7362));
 sg13g2_o21ai_1 _17248_ (.B1(_03667_),
    .Y(_03668_),
    .A1(net7282),
    .A2(net7256));
 sg13g2_nand2_1 _17249_ (.Y(_03669_),
    .A(_08250_),
    .B(_03668_));
 sg13g2_nand3_1 _17250_ (.B(net7384),
    .C(net7429),
    .A(_01635_),
    .Y(_03670_));
 sg13g2_nand2_1 _17251_ (.Y(_03671_),
    .A(_03669_),
    .B(_03670_));
 sg13g2_and3_1 _17252_ (.X(_03672_),
    .A(net7805),
    .B(net7432),
    .C(_03639_));
 sg13g2_a221oi_1 _17253_ (.B2(_01943_),
    .C1(_03672_),
    .B1(_03653_),
    .A1(_01975_),
    .Y(_03673_),
    .A2(net7362));
 sg13g2_o21ai_1 _17254_ (.B1(_03673_),
    .Y(_03674_),
    .A1(_13358_),
    .A2(net7256));
 sg13g2_nand2_1 _17255_ (.Y(_03675_),
    .A(net7366),
    .B(_03674_));
 sg13g2_nand3_1 _17256_ (.B(net7383),
    .C(net7428),
    .A(_01636_),
    .Y(_03676_));
 sg13g2_nand2_1 _17257_ (.Y(_03677_),
    .A(_03675_),
    .B(_03676_));
 sg13g2_a22oi_1 _17258_ (.Y(_03678_),
    .B1(net7252),
    .B2(_01944_),
    .A2(net7356),
    .A1(_01976_));
 sg13g2_o21ai_1 _17259_ (.B1(_03678_),
    .Y(_03679_),
    .A1(net7275),
    .A2(net7256));
 sg13g2_nand2_1 _17260_ (.Y(_03680_),
    .A(net7366),
    .B(_03679_));
 sg13g2_nand3_1 _17261_ (.B(net7379),
    .C(net7429),
    .A(_01637_),
    .Y(_03681_));
 sg13g2_nand2_1 _17262_ (.Y(_03682_),
    .A(_03680_),
    .B(_03681_));
 sg13g2_a22oi_1 _17263_ (.Y(_03683_),
    .B1(net7252),
    .B2(_01945_),
    .A2(net7356),
    .A1(_01977_));
 sg13g2_o21ai_1 _17264_ (.B1(_03683_),
    .Y(_03684_),
    .A1(net7273),
    .A2(net7255));
 sg13g2_nand2_1 _17265_ (.Y(_03685_),
    .A(net7366),
    .B(_03684_));
 sg13g2_nand3_1 _17266_ (.B(net7383),
    .C(net7426),
    .A(_01639_),
    .Y(_03686_));
 sg13g2_nand2_1 _17267_ (.Y(_03687_),
    .A(_03685_),
    .B(_03686_));
 sg13g2_a22oi_1 _17268_ (.Y(_03688_),
    .B1(net7252),
    .B2(_01946_),
    .A2(net7356),
    .A1(_01978_));
 sg13g2_o21ai_1 _17269_ (.B1(_03688_),
    .Y(_03689_),
    .A1(_15563_),
    .A2(net7256));
 sg13g2_nand2_1 _17270_ (.Y(_03690_),
    .A(net7365),
    .B(_03689_));
 sg13g2_nand3_1 _17271_ (.B(net7379),
    .C(net7429),
    .A(_01640_),
    .Y(_03691_));
 sg13g2_nand2_1 _17272_ (.Y(_03692_),
    .A(_03690_),
    .B(_03691_));
 sg13g2_nor2_1 _17273_ (.A(_02067_),
    .B(net7256),
    .Y(_03693_));
 sg13g2_a221oi_1 _17274_ (.B2(_01947_),
    .C1(_03693_),
    .B1(net7251),
    .A1(_01979_),
    .Y(_03694_),
    .A2(net7359));
 sg13g2_inv_1 _17275_ (.Y(_03695_),
    .A(net7022));
 sg13g2_a21oi_1 _17276_ (.A1(_01641_),
    .A2(net7428),
    .Y(_03696_),
    .B1(net7376));
 sg13g2_a21oi_1 _17277_ (.A1(net7364),
    .A2(_03694_),
    .Y(_03697_),
    .B1(_03696_));
 sg13g2_a22oi_1 _17278_ (.Y(_03698_),
    .B1(net7251),
    .B2(_01948_),
    .A2(net7355),
    .A1(_01980_));
 sg13g2_o21ai_1 _17279_ (.B1(_03698_),
    .Y(_03699_),
    .A1(net7349),
    .A2(net7255));
 sg13g2_nand2_1 _17280_ (.Y(_03700_),
    .A(net7366),
    .B(_03699_));
 sg13g2_nand3_1 _17281_ (.B(net7380),
    .C(net7429),
    .A(_01642_),
    .Y(_03701_));
 sg13g2_nand2_1 _17282_ (.Y(_03702_),
    .A(_03700_),
    .B(_03701_));
 sg13g2_a22oi_1 _17283_ (.Y(_03703_),
    .B1(_03653_),
    .B2(_01918_),
    .A2(net7355),
    .A1(_01950_));
 sg13g2_o21ai_1 _17284_ (.B1(_03703_),
    .Y(_03704_),
    .A1(_02206_),
    .A2(net7258));
 sg13g2_nand2_1 _17285_ (.Y(_03705_),
    .A(_08250_),
    .B(net7020));
 sg13g2_nand3_1 _17286_ (.B(net7384),
    .C(net7428),
    .A(_01643_),
    .Y(_03706_));
 sg13g2_nand2_1 _17287_ (.Y(_03707_),
    .A(_03705_),
    .B(_03706_));
 sg13g2_a22oi_1 _17288_ (.Y(_03708_),
    .B1(net7252),
    .B2(_01919_),
    .A2(net7356),
    .A1(_01951_));
 sg13g2_o21ai_1 _17289_ (.B1(_03708_),
    .Y(_03709_),
    .A1(_02283_),
    .A2(net7255));
 sg13g2_nand2_1 _17290_ (.Y(_03710_),
    .A(net7365),
    .B(_03709_));
 sg13g2_nand3_1 _17291_ (.B(net7380),
    .C(net7429),
    .A(_01644_),
    .Y(_03711_));
 sg13g2_nand2_1 _17292_ (.Y(_03712_),
    .A(_03710_),
    .B(_03711_));
 sg13g2_a22oi_1 _17293_ (.Y(_03713_),
    .B1(net7251),
    .B2(_01920_),
    .A2(net7355),
    .A1(_01952_));
 sg13g2_o21ai_1 _17294_ (.B1(_03713_),
    .Y(_03714_),
    .A1(_02361_),
    .A2(net7255));
 sg13g2_nand2_1 _17295_ (.Y(_03715_),
    .A(net7365),
    .B(_03714_));
 sg13g2_nand3_1 _17296_ (.B(net7380),
    .C(net7428),
    .A(_01645_),
    .Y(_03716_));
 sg13g2_nand2_1 _17297_ (.Y(_03717_),
    .A(_03715_),
    .B(_03716_));
 sg13g2_a22oi_1 _17298_ (.Y(_03718_),
    .B1(net7251),
    .B2(_01921_),
    .A2(net7355),
    .A1(_01953_));
 sg13g2_o21ai_1 _17299_ (.B1(_03718_),
    .Y(_03719_),
    .A1(_02439_),
    .A2(net7255));
 sg13g2_nand2_1 _17300_ (.Y(_03720_),
    .A(net7365),
    .B(_03719_));
 sg13g2_nand3_1 _17301_ (.B(net7383),
    .C(net7429),
    .A(_01646_),
    .Y(_03721_));
 sg13g2_nand2_1 _17302_ (.Y(_03722_),
    .A(_03720_),
    .B(_03721_));
 sg13g2_a22oi_1 _17303_ (.Y(_03723_),
    .B1(net7251),
    .B2(_01922_),
    .A2(net7359),
    .A1(_01954_));
 sg13g2_o21ai_1 _17304_ (.B1(_03723_),
    .Y(_03724_),
    .A1(_02503_),
    .A2(net7255));
 sg13g2_nand2_1 _17305_ (.Y(_03725_),
    .A(net7365),
    .B(net7016));
 sg13g2_nand3_1 _17306_ (.B(net7380),
    .C(net7428),
    .A(_01647_),
    .Y(_03726_));
 sg13g2_nand2_1 _17307_ (.Y(_03727_),
    .A(_03725_),
    .B(_03726_));
 sg13g2_a22oi_1 _17308_ (.Y(_03728_),
    .B1(net7251),
    .B2(_01923_),
    .A2(net7359),
    .A1(_01955_));
 sg13g2_inv_1 _17309_ (.Y(_03729_),
    .A(_03730_));
 sg13g2_o21ai_1 _17310_ (.B1(_03728_),
    .Y(_03730_),
    .A1(_02549_),
    .A2(net7256));
 sg13g2_a21oi_1 _17311_ (.A1(_01648_),
    .A2(net7425),
    .Y(_03731_),
    .B1(net7371));
 sg13g2_a21oi_1 _17312_ (.A1(net7372),
    .A2(_03729_),
    .Y(_03732_),
    .B1(_03731_));
 sg13g2_a22oi_1 _17313_ (.Y(_03733_),
    .B1(net7252),
    .B2(_01924_),
    .A2(net7356),
    .A1(_01956_));
 sg13g2_inv_1 _17314_ (.Y(_03734_),
    .A(_03735_));
 sg13g2_o21ai_1 _17315_ (.B1(_03733_),
    .Y(_03735_),
    .A1(_02615_),
    .A2(net7255));
 sg13g2_a21oi_1 _17316_ (.A1(_01650_),
    .A2(net7427),
    .Y(_03736_),
    .B1(net7371));
 sg13g2_a21oi_1 _17317_ (.A1(net7373),
    .A2(_03734_),
    .Y(_03737_),
    .B1(_03736_));
 sg13g2_a22oi_1 _17318_ (.Y(_03738_),
    .B1(net7252),
    .B2(_01925_),
    .A2(net7356),
    .A1(_01957_));
 sg13g2_o21ai_1 _17319_ (.B1(_03738_),
    .Y(_03739_),
    .A1(net7344),
    .A2(net7257));
 sg13g2_nand2_1 _17320_ (.Y(_03740_),
    .A(net7373),
    .B(_03739_));
 sg13g2_nand3_1 _17321_ (.B(net7381),
    .C(net7426),
    .A(_01651_),
    .Y(_03741_));
 sg13g2_nand2_1 _17322_ (.Y(_03742_),
    .A(_03740_),
    .B(_03741_));
 sg13g2_a22oi_1 _17323_ (.Y(_03743_),
    .B1(net7252),
    .B2(_01926_),
    .A2(net7356),
    .A1(_01958_));
 sg13g2_o21ai_1 _17324_ (.B1(_03743_),
    .Y(_03744_),
    .A1(net7343),
    .A2(net7257));
 sg13g2_nand2_1 _17325_ (.Y(_03745_),
    .A(net7372),
    .B(_03744_));
 sg13g2_nand3_1 _17326_ (.B(net7383),
    .C(net7426),
    .A(_01652_),
    .Y(_03746_));
 sg13g2_nand2_1 _17327_ (.Y(_03747_),
    .A(_03745_),
    .B(_03746_));
 sg13g2_a22oi_1 _17328_ (.Y(_03748_),
    .B1(net7254),
    .B2(_01927_),
    .A2(net7358),
    .A1(_01959_));
 sg13g2_o21ai_1 _17329_ (.B1(_03748_),
    .Y(_03749_),
    .A1(_02818_),
    .A2(net7257));
 sg13g2_nand2_1 _17330_ (.Y(_03750_),
    .A(net7372),
    .B(net7012));
 sg13g2_nand3_1 _17331_ (.B(net7381),
    .C(net7426),
    .A(_01653_),
    .Y(_03751_));
 sg13g2_nand2_1 _17332_ (.Y(_03752_),
    .A(_03750_),
    .B(_03751_));
 sg13g2_nor2_1 _17333_ (.A(_02886_),
    .B(net7258),
    .Y(_03753_));
 sg13g2_a221oi_1 _17334_ (.B2(_01929_),
    .C1(_03753_),
    .B1(net7254),
    .A1(_01961_),
    .Y(_03754_),
    .A2(net7358));
 sg13g2_inv_1 _17335_ (.Y(_03755_),
    .A(_03754_));
 sg13g2_a21oi_1 _17336_ (.A1(net7980),
    .A2(net7425),
    .Y(_03756_),
    .B1(net7369));
 sg13g2_a21oi_1 _17337_ (.A1(net7372),
    .A2(_03754_),
    .Y(_03757_),
    .B1(_03756_));
 sg13g2_nor2_1 _17338_ (.A(_02951_),
    .B(net7258),
    .Y(_03758_));
 sg13g2_a221oi_1 _17339_ (.B2(_01930_),
    .C1(_03758_),
    .B1(net7253),
    .A1(_01962_),
    .Y(_03759_),
    .A2(net7357));
 sg13g2_inv_1 _17340_ (.Y(_03760_),
    .A(_03759_));
 sg13g2_a21oi_1 _17341_ (.A1(net7979),
    .A2(net7425),
    .Y(_03761_),
    .B1(net7369));
 sg13g2_a21oi_1 _17342_ (.A1(net7369),
    .A2(_03759_),
    .Y(_03762_),
    .B1(_03761_));
 sg13g2_nor2_1 _17343_ (.A(_03018_),
    .B(net7258),
    .Y(_03763_));
 sg13g2_a221oi_1 _17344_ (.B2(_01931_),
    .C1(_03763_),
    .B1(net7253),
    .A1(_01963_),
    .Y(_03764_),
    .A2(net7357));
 sg13g2_inv_1 _17345_ (.Y(_03765_),
    .A(_03764_));
 sg13g2_a21oi_1 _17346_ (.A1(_01656_),
    .A2(net7425),
    .Y(_03766_),
    .B1(net7368));
 sg13g2_a21oi_1 _17347_ (.A1(net7368),
    .A2(_03764_),
    .Y(_03767_),
    .B1(_03766_));
 sg13g2_a22oi_1 _17348_ (.Y(_03768_),
    .B1(net7253),
    .B2(_01932_),
    .A2(net7357),
    .A1(_01964_));
 sg13g2_o21ai_1 _17349_ (.B1(_03768_),
    .Y(_03769_),
    .A1(_03085_),
    .A2(net7257));
 sg13g2_nand2_1 _17350_ (.Y(_03770_),
    .A(net7371),
    .B(_03769_));
 sg13g2_nand3_1 _17351_ (.B(net7381),
    .C(net7427),
    .A(net7978),
    .Y(_03771_));
 sg13g2_nand2_1 _17352_ (.Y(_03772_),
    .A(_03770_),
    .B(_03771_));
 sg13g2_a22oi_1 _17353_ (.Y(_03773_),
    .B1(net7253),
    .B2(_01933_),
    .A2(net7357),
    .A1(_01965_));
 sg13g2_o21ai_1 _17354_ (.B1(_03773_),
    .Y(_03774_),
    .A1(net7334),
    .A2(net7257));
 sg13g2_nand2_1 _17355_ (.Y(_03775_),
    .A(net7367),
    .B(net7010));
 sg13g2_nand3_1 _17356_ (.B(net7381),
    .C(net7425),
    .A(_01658_),
    .Y(_03776_));
 sg13g2_nand2_1 _17357_ (.Y(_03777_),
    .A(_03775_),
    .B(_03776_));
 sg13g2_nor2_1 _17358_ (.A(net7333),
    .B(net7258),
    .Y(_03778_));
 sg13g2_a221oi_1 _17359_ (.B2(_01934_),
    .C1(_03778_),
    .B1(net7253),
    .A1(_01966_),
    .Y(_03779_),
    .A2(net7357));
 sg13g2_inv_1 _17360_ (.Y(_03780_),
    .A(net7009));
 sg13g2_a21oi_1 _17361_ (.A1(_01659_),
    .A2(net7425),
    .Y(_03781_),
    .B1(net7369));
 sg13g2_a21oi_1 _17362_ (.A1(net7369),
    .A2(_03779_),
    .Y(_03782_),
    .B1(_03781_));
 sg13g2_nor2_1 _17363_ (.A(net7332),
    .B(net7258),
    .Y(_03783_));
 sg13g2_a221oi_1 _17364_ (.B2(_01935_),
    .C1(_03783_),
    .B1(net7253),
    .A1(_01967_),
    .Y(_03784_),
    .A2(net7357));
 sg13g2_inv_1 _17365_ (.Y(_03785_),
    .A(_03784_));
 sg13g2_a21oi_1 _17366_ (.A1(_01661_),
    .A2(net7425),
    .Y(_03786_),
    .B1(net7369));
 sg13g2_a21oi_1 _17367_ (.A1(net7369),
    .A2(_03784_),
    .Y(_03787_),
    .B1(_03786_));
 sg13g2_a22oi_1 _17368_ (.Y(_03788_),
    .B1(net7253),
    .B2(_01936_),
    .A2(net7357),
    .A1(_01968_));
 sg13g2_o21ai_1 _17369_ (.B1(_03788_),
    .Y(_03789_),
    .A1(_03367_),
    .A2(net7257));
 sg13g2_nand2_1 _17370_ (.Y(_03790_),
    .A(net7372),
    .B(_03789_));
 sg13g2_nand3_1 _17371_ (.B(net7381),
    .C(net7427),
    .A(_01662_),
    .Y(_03791_));
 sg13g2_nand2_1 _17372_ (.Y(_03792_),
    .A(_03790_),
    .B(_03791_));
 sg13g2_nor2_1 _17373_ (.A(net7331),
    .B(net7257),
    .Y(_03793_));
 sg13g2_a22oi_1 _17374_ (.Y(_03794_),
    .B1(net7253),
    .B2(_01937_),
    .A2(net7357),
    .A1(_01969_));
 sg13g2_nor2b_1 _17375_ (.A(_03793_),
    .B_N(_03794_),
    .Y(_03795_));
 sg13g2_nand2b_1 _17376_ (.Y(_03796_),
    .B(_03794_),
    .A_N(_03793_));
 sg13g2_a21oi_1 _17377_ (.A1(_01663_),
    .A2(net7425),
    .Y(_03797_),
    .B1(net7368));
 sg13g2_a21oi_1 _17378_ (.A1(net7367),
    .A2(_03795_),
    .Y(_03798_),
    .B1(_03797_));
 sg13g2_a22oi_1 _17379_ (.Y(_03799_),
    .B1(net7254),
    .B2(_01938_),
    .A2(net7358),
    .A1(_01970_));
 sg13g2_o21ai_1 _17380_ (.B1(_03799_),
    .Y(_03800_),
    .A1(_03505_),
    .A2(net7257));
 sg13g2_nand2_1 _17381_ (.Y(_03801_),
    .A(net7372),
    .B(_03800_));
 sg13g2_nand3_1 _17382_ (.B(net7381),
    .C(net7427),
    .A(_01664_),
    .Y(_03802_));
 sg13g2_nand2_1 _17383_ (.Y(_03803_),
    .A(_03801_),
    .B(_03802_));
 sg13g2_a22oi_1 _17384_ (.Y(_03804_),
    .B1(net7252),
    .B2(_01940_),
    .A2(net7356),
    .A1(_01972_));
 sg13g2_o21ai_1 _17385_ (.B1(_03804_),
    .Y(_03805_),
    .A1(net7328),
    .A2(net7256));
 sg13g2_nand2_1 _17386_ (.Y(_03806_),
    .A(net7373),
    .B(net7006));
 sg13g2_nand3_1 _17387_ (.B(net7381),
    .C(net7427),
    .A(_01665_),
    .Y(_03807_));
 sg13g2_nand2_1 _17388_ (.Y(_03808_),
    .A(_03806_),
    .B(_03807_));
 sg13g2_nand3_1 _17389_ (.B(_03642_),
    .C(_03645_),
    .A(_03629_),
    .Y(_03809_));
 sg13g2_a22oi_1 _17390_ (.Y(_03810_),
    .B1(net7251),
    .B2(_01941_),
    .A2(net7355),
    .A1(_01973_));
 sg13g2_and2_1 _17391_ (.A(_03809_),
    .B(_03810_),
    .X(_03811_));
 sg13g2_nand2_1 _17392_ (.Y(_03812_),
    .A(_03809_),
    .B(_03810_));
 sg13g2_a21oi_1 _17393_ (.A1(net7977),
    .A2(net7427),
    .Y(_03813_),
    .B1(net7370));
 sg13g2_a21oi_1 _17394_ (.A1(net7370),
    .A2(_03811_),
    .Y(_03814_),
    .B1(_03813_));
 sg13g2_or2_1 _17395_ (.X(_03815_),
    .B(_00537_),
    .A(net8016));
 sg13g2_nand3b_1 _17396_ (.B(_07792_),
    .C(_07812_),
    .Y(_03816_),
    .A_N(_08238_));
 sg13g2_a21o_1 _17397_ (.A2(_03816_),
    .A1(_00536_),
    .B1(net7637),
    .X(_03817_));
 sg13g2_nor2_1 _17398_ (.A(_05195_),
    .B(_03816_),
    .Y(_03818_));
 sg13g2_nor3_1 _17399_ (.A(_05195_),
    .B(net7607),
    .C(net7376),
    .Y(_03819_));
 sg13g2_a22oi_1 _17400_ (.Y(_03820_),
    .B1(net7319),
    .B2(_01632_),
    .A2(net7327),
    .A1(_01650_));
 sg13g2_nor2_1 _17401_ (.A(_00538_),
    .B(_00536_),
    .Y(_03821_));
 sg13g2_or2_1 _17402_ (.X(_03822_),
    .B(_00536_),
    .A(net8016));
 sg13g2_nand2b_1 _17403_ (.Y(_03823_),
    .B(_00004_),
    .A_N(_00537_));
 sg13g2_nand2_1 _17404_ (.Y(_03824_),
    .A(net7284),
    .B(_03823_));
 sg13g2_a22oi_1 _17405_ (.Y(_03825_),
    .B1(_03823_),
    .B2(net7284),
    .A2(_03822_),
    .A1(_02616_));
 sg13g2_o21ai_1 _17406_ (.B1(_03824_),
    .Y(_03826_),
    .A1(net7346),
    .A2(_03821_));
 sg13g2_nand2_1 _17407_ (.Y(_03827_),
    .A(_05195_),
    .B(_00004_));
 sg13g2_and4_1 _17408_ (.A(_08420_),
    .B(_08460_),
    .C(_08557_),
    .D(net7441),
    .X(_03828_));
 sg13g2_a22oi_1 _17409_ (.Y(_03829_),
    .B1(_03828_),
    .B2(_08381_),
    .A2(net7639),
    .A1(_02584_));
 sg13g2_nor3_1 _17410_ (.A(_03820_),
    .B(net7248),
    .C(net7242),
    .Y(_03830_));
 sg13g2_o21ai_1 _17411_ (.B1(_03820_),
    .Y(_03831_),
    .A1(net7250),
    .A2(net7246));
 sg13g2_nor2b_1 _17412_ (.A(_03830_),
    .B_N(_03831_),
    .Y(_03832_));
 sg13g2_nand2b_1 _17413_ (.Y(_03833_),
    .B(_03822_),
    .A_N(net7344));
 sg13g2_nand3_1 _17414_ (.B(_10351_),
    .C(net7634),
    .A(_10200_),
    .Y(_03834_));
 sg13g2_and2_1 _17415_ (.A(_03833_),
    .B(_03834_),
    .X(_03835_));
 sg13g2_nand2_1 _17416_ (.Y(_03836_),
    .A(_03833_),
    .B(net7241));
 sg13g2_a21oi_1 _17417_ (.A1(_03833_),
    .A2(_03834_),
    .Y(_03837_),
    .B1(net7245));
 sg13g2_and3_1 _17418_ (.X(_03838_),
    .A(_09816_),
    .B(_09900_),
    .C(net7441));
 sg13g2_a22oi_1 _17419_ (.Y(_03839_),
    .B1(_03838_),
    .B2(_09684_),
    .A2(net7639),
    .A1(net7345));
 sg13g2_or2_1 _17420_ (.X(_03840_),
    .B(net7234),
    .A(net7248));
 sg13g2_xnor2_1 _17421_ (.Y(_03841_),
    .A(_03837_),
    .B(_03840_));
 sg13g2_a22oi_1 _17422_ (.Y(_03842_),
    .B1(net7319),
    .B2(_01633_),
    .A2(net7327),
    .A1(_01651_));
 sg13g2_xor2_1 _17423_ (.B(_03842_),
    .A(_03830_),
    .X(_03843_));
 sg13g2_xnor2_1 _17424_ (.Y(_03844_),
    .A(_03841_),
    .B(_03843_));
 sg13g2_nor2_1 _17425_ (.A(net7069),
    .B(net7234),
    .Y(_03845_));
 sg13g2_a22oi_1 _17426_ (.Y(_03846_),
    .B1(net7632),
    .B2(_11150_),
    .A2(net7635),
    .A1(_02745_));
 sg13g2_a22oi_1 _17427_ (.Y(_03847_),
    .B1(net7319),
    .B2(_01634_),
    .A2(net7327),
    .A1(_01652_));
 sg13g2_o21ai_1 _17428_ (.B1(_03847_),
    .Y(_03848_),
    .A1(net7242),
    .A2(net7229));
 sg13g2_nor3_1 _17429_ (.A(net7242),
    .B(net7229),
    .C(_03847_),
    .Y(_03849_));
 sg13g2_or3_1 _17430_ (.A(net7242),
    .B(net7229),
    .C(_03847_),
    .X(_03850_));
 sg13g2_nand2_1 _17431_ (.Y(_03851_),
    .A(_03848_),
    .B(_03850_));
 sg13g2_xor2_1 _17432_ (.B(_03851_),
    .A(_03845_),
    .X(_03852_));
 sg13g2_or3_1 _17433_ (.A(net7245),
    .B(net7069),
    .C(_03840_),
    .X(_03853_));
 sg13g2_nor2_1 _17434_ (.A(_03842_),
    .B(_03853_),
    .Y(_03854_));
 sg13g2_nor2b_1 _17435_ (.A(_03837_),
    .B_N(_03840_),
    .Y(_03855_));
 sg13g2_a22oi_1 _17436_ (.Y(_03856_),
    .B1(_03855_),
    .B2(_03842_),
    .A2(_03854_),
    .A1(_03830_));
 sg13g2_o21ai_1 _17437_ (.B1(_03853_),
    .Y(_03857_),
    .A1(_03842_),
    .A2(_03855_));
 sg13g2_o21ai_1 _17438_ (.B1(_03856_),
    .Y(_03858_),
    .A1(_03830_),
    .A2(_03857_));
 sg13g2_xor2_1 _17439_ (.B(_03858_),
    .A(_03852_),
    .X(_03859_));
 sg13g2_and4_1 _17440_ (.A(_10612_),
    .B(_10646_),
    .C(_10733_),
    .D(net7441),
    .X(_03860_));
 sg13g2_and3_1 _17441_ (.X(_03861_),
    .A(_02697_),
    .B(_02702_),
    .C(net7639));
 sg13g2_a22oi_1 _17442_ (.Y(_03862_),
    .B1(_03861_),
    .B2(_02712_),
    .A2(_03860_),
    .A1(_10581_));
 sg13g2_inv_1 _17443_ (.Y(_03863_),
    .A(_03862_));
 sg13g2_nor2_1 _17444_ (.A(net7248),
    .B(net7226),
    .Y(_03864_));
 sg13g2_xor2_1 _17445_ (.B(_03864_),
    .A(_03859_),
    .X(_03865_));
 sg13g2_nand2_1 _17446_ (.Y(_03866_),
    .A(_03859_),
    .B(_03864_));
 sg13g2_nor2_1 _17447_ (.A(net7234),
    .B(net7229),
    .Y(_03867_));
 sg13g2_a22oi_1 _17448_ (.Y(_03868_),
    .B1(net7319),
    .B2(_01635_),
    .A2(net7327),
    .A1(_01653_));
 sg13g2_a22oi_1 _17449_ (.Y(_03869_),
    .B1(net7632),
    .B2(_12225_),
    .A2(net7635),
    .A1(_02817_));
 sg13g2_nor3_1 _17450_ (.A(net7242),
    .B(_03868_),
    .C(net7221),
    .Y(_03870_));
 sg13g2_o21ai_1 _17451_ (.B1(_03868_),
    .Y(_03871_),
    .A1(net7242),
    .A2(net7221));
 sg13g2_nor2b_1 _17452_ (.A(_03870_),
    .B_N(_03871_),
    .Y(_03872_));
 sg13g2_xnor2_1 _17453_ (.Y(_03873_),
    .A(_03867_),
    .B(_03872_));
 sg13g2_o21ai_1 _17454_ (.B1(_03848_),
    .Y(_03874_),
    .A1(_03849_),
    .A2(_03857_));
 sg13g2_nor2b_1 _17455_ (.A(_03845_),
    .B_N(_03874_),
    .Y(_03875_));
 sg13g2_nand3_1 _17456_ (.B(_03849_),
    .C(_03857_),
    .A(_03845_),
    .Y(_03876_));
 sg13g2_o21ai_1 _17457_ (.B1(_03876_),
    .Y(_03877_),
    .A1(_03848_),
    .A2(_03857_));
 sg13g2_nor2_1 _17458_ (.A(_03875_),
    .B(_03877_),
    .Y(_03878_));
 sg13g2_xnor2_1 _17459_ (.Y(_03879_),
    .A(_03873_),
    .B(_03878_));
 sg13g2_o21ai_1 _17460_ (.B1(net7441),
    .Y(_03880_),
    .A1(_08389_),
    .A2(_11474_));
 sg13g2_nor3_1 _17461_ (.A(_11524_),
    .B(_11648_),
    .C(_03880_),
    .Y(_03881_));
 sg13g2_and3_1 _17462_ (.X(_03882_),
    .A(_02762_),
    .B(_02767_),
    .C(net7639));
 sg13g2_a22oi_1 _17463_ (.Y(_03883_),
    .B1(_03882_),
    .B2(_02777_),
    .A2(_03881_),
    .A1(_11432_));
 sg13g2_nor2_1 _17464_ (.A(net7248),
    .B(net7218),
    .Y(_03884_));
 sg13g2_nor2_1 _17465_ (.A(net7069),
    .B(net7226),
    .Y(_03885_));
 sg13g2_xnor2_1 _17466_ (.Y(_03886_),
    .A(_03884_),
    .B(_03885_));
 sg13g2_mux2_1 _17467_ (.A0(_03855_),
    .A1(_03841_),
    .S(_03842_),
    .X(_03887_));
 sg13g2_mux2_1 _17468_ (.A0(_03887_),
    .A1(_03854_),
    .S(_03852_),
    .X(_03888_));
 sg13g2_nand2_1 _17469_ (.Y(_03889_),
    .A(_03830_),
    .B(_03888_));
 sg13g2_nor2_1 _17470_ (.A(_03886_),
    .B(_03889_),
    .Y(_03890_));
 sg13g2_and2_1 _17471_ (.A(_03886_),
    .B(_03889_),
    .X(_03891_));
 sg13g2_inv_1 _17472_ (.Y(_03892_),
    .A(_03891_));
 sg13g2_nor2_1 _17473_ (.A(_03890_),
    .B(_03891_),
    .Y(_03893_));
 sg13g2_xnor2_1 _17474_ (.Y(_03894_),
    .A(_03879_),
    .B(_03893_));
 sg13g2_nor2_1 _17475_ (.A(_03866_),
    .B(_03894_),
    .Y(_03895_));
 sg13g2_xor2_1 _17476_ (.B(_03894_),
    .A(_03866_),
    .X(_03896_));
 sg13g2_mux2_1 _17477_ (.A0(_03848_),
    .A1(_03850_),
    .S(_03873_),
    .X(_03897_));
 sg13g2_nor2b_1 _17478_ (.A(_03897_),
    .B_N(_03845_),
    .Y(_03898_));
 sg13g2_nor3_1 _17479_ (.A(_03845_),
    .B(_03851_),
    .C(_03873_),
    .Y(_03899_));
 sg13g2_o21ai_1 _17480_ (.B1(_03857_),
    .Y(_03900_),
    .A1(_03898_),
    .A2(_03899_));
 sg13g2_or2_1 _17481_ (.X(_03901_),
    .B(net7226),
    .A(net7229));
 sg13g2_nor2_1 _17482_ (.A(net7069),
    .B(net7218),
    .Y(_03902_));
 sg13g2_and3_1 _17483_ (.X(_03903_),
    .A(_02833_),
    .B(_02838_),
    .C(net7639));
 sg13g2_a22oi_1 _17484_ (.Y(_03904_),
    .B1(_03903_),
    .B2(net7342),
    .A2(net7440),
    .A1(_12788_));
 sg13g2_nor2_1 _17485_ (.A(net7248),
    .B(net7213),
    .Y(_03905_));
 sg13g2_xnor2_1 _17486_ (.Y(_03906_),
    .A(_03901_),
    .B(_03905_));
 sg13g2_xnor2_1 _17487_ (.Y(_03907_),
    .A(_03902_),
    .B(_03906_));
 sg13g2_a22oi_1 _17488_ (.Y(_03908_),
    .B1(net7634),
    .B2(_13356_),
    .A2(net7636),
    .A1(_02885_));
 sg13g2_nor2_1 _17489_ (.A(net7242),
    .B(net7211),
    .Y(_03909_));
 sg13g2_a22oi_1 _17490_ (.Y(_03910_),
    .B1(net7319),
    .B2(_01636_),
    .A2(net7327),
    .A1(net7980));
 sg13g2_nor2_1 _17491_ (.A(net7234),
    .B(net7221),
    .Y(_03911_));
 sg13g2_o21ai_1 _17492_ (.B1(_03910_),
    .Y(_03912_),
    .A1(net7234),
    .A2(net7221));
 sg13g2_nor3_1 _17493_ (.A(net7234),
    .B(net7221),
    .C(_03910_),
    .Y(_03913_));
 sg13g2_xor2_1 _17494_ (.B(_03911_),
    .A(_03910_),
    .X(_03914_));
 sg13g2_xnor2_1 _17495_ (.Y(_03915_),
    .A(_03909_),
    .B(_03914_));
 sg13g2_a21oi_1 _17496_ (.A1(_03867_),
    .A2(_03871_),
    .Y(_03916_),
    .B1(_03870_));
 sg13g2_nand2_1 _17497_ (.Y(_03917_),
    .A(_03864_),
    .B(_03902_));
 sg13g2_nor2_1 _17498_ (.A(_03916_),
    .B(_03917_),
    .Y(_03918_));
 sg13g2_nand2_1 _17499_ (.Y(_03919_),
    .A(_03916_),
    .B(_03917_));
 sg13g2_xor2_1 _17500_ (.B(_03917_),
    .A(_03916_),
    .X(_03920_));
 sg13g2_xnor2_1 _17501_ (.Y(_03921_),
    .A(_03915_),
    .B(_03920_));
 sg13g2_a21oi_1 _17502_ (.A1(_03845_),
    .A2(_03848_),
    .Y(_03922_),
    .B1(_03849_));
 sg13g2_nor2_1 _17503_ (.A(_03873_),
    .B(_03922_),
    .Y(_03923_));
 sg13g2_nand2b_1 _17504_ (.Y(_03924_),
    .B(_03923_),
    .A_N(_03921_));
 sg13g2_xor2_1 _17505_ (.B(_03923_),
    .A(_03921_),
    .X(_03925_));
 sg13g2_nand2_1 _17506_ (.Y(_03926_),
    .A(_03907_),
    .B(_03925_));
 sg13g2_xnor2_1 _17507_ (.Y(_03927_),
    .A(_03907_),
    .B(_03925_));
 sg13g2_xnor2_1 _17508_ (.Y(_03928_),
    .A(_03900_),
    .B(_03927_));
 sg13g2_a21oi_1 _17509_ (.A1(_03879_),
    .A2(_03892_),
    .Y(_03929_),
    .B1(_03890_));
 sg13g2_xor2_1 _17510_ (.B(_03929_),
    .A(_03928_),
    .X(_03930_));
 sg13g2_a22oi_1 _17511_ (.Y(_03931_),
    .B1(net7633),
    .B2(_14253_),
    .A2(net7636),
    .A1(_02950_));
 sg13g2_nor2_1 _17512_ (.A(net7246),
    .B(net7209),
    .Y(_03932_));
 sg13g2_a22oi_1 _17513_ (.Y(_03933_),
    .B1(net7319),
    .B2(_01637_),
    .A2(net7326),
    .A1(net7979));
 sg13g2_nor3_1 _17514_ (.A(net7239),
    .B(net7211),
    .C(_03933_),
    .Y(_03934_));
 sg13g2_o21ai_1 _17515_ (.B1(_03933_),
    .Y(_03935_),
    .A1(net7239),
    .A2(net7211));
 sg13g2_nor2b_1 _17516_ (.A(_03934_),
    .B_N(_03935_),
    .Y(_03936_));
 sg13g2_xnor2_1 _17517_ (.Y(_03937_),
    .A(_03932_),
    .B(_03936_));
 sg13g2_nor3_1 _17518_ (.A(net7069),
    .B(net7218),
    .C(_03901_),
    .Y(_03938_));
 sg13g2_o21ai_1 _17519_ (.B1(_03901_),
    .Y(_03939_),
    .A1(net7069),
    .A2(net7218));
 sg13g2_a21oi_1 _17520_ (.A1(_03905_),
    .A2(_03939_),
    .Y(_03940_),
    .B1(_03938_));
 sg13g2_a21oi_1 _17521_ (.A1(_03909_),
    .A2(_03912_),
    .Y(_03941_),
    .B1(_03913_));
 sg13g2_xnor2_1 _17522_ (.Y(_03942_),
    .A(_03940_),
    .B(_03941_));
 sg13g2_xnor2_1 _17523_ (.Y(_03943_),
    .A(_03937_),
    .B(_03942_));
 sg13g2_a21oi_1 _17524_ (.A1(_03915_),
    .A2(_03919_),
    .Y(_03944_),
    .B1(_03918_));
 sg13g2_xnor2_1 _17525_ (.Y(_03945_),
    .A(_03943_),
    .B(_03944_));
 sg13g2_a21oi_1 _17526_ (.A1(_03833_),
    .A2(_03834_),
    .Y(_03946_),
    .B1(net7213));
 sg13g2_nor2_1 _17527_ (.A(net7229),
    .B(net7217),
    .Y(_03947_));
 sg13g2_nor2_1 _17528_ (.A(net7226),
    .B(net7221),
    .Y(_03948_));
 sg13g2_xnor2_1 _17529_ (.Y(_03949_),
    .A(_03947_),
    .B(_03948_));
 sg13g2_xnor2_1 _17530_ (.Y(_03950_),
    .A(_03946_),
    .B(_03949_));
 sg13g2_and4_1 _17531_ (.A(_13629_),
    .B(_13681_),
    .C(_13783_),
    .D(net7440),
    .X(_03951_));
 sg13g2_a22oi_1 _17532_ (.Y(_03952_),
    .B1(_03951_),
    .B2(_13580_),
    .A2(net7638),
    .A1(_02918_));
 sg13g2_nor2_1 _17533_ (.A(net7247),
    .B(net7205),
    .Y(_03953_));
 sg13g2_xnor2_1 _17534_ (.Y(_03954_),
    .A(_03950_),
    .B(_03953_));
 sg13g2_and2_1 _17535_ (.A(_03924_),
    .B(_03954_),
    .X(_03955_));
 sg13g2_xnor2_1 _17536_ (.Y(_03956_),
    .A(_03924_),
    .B(_03954_));
 sg13g2_xnor2_1 _17537_ (.Y(_03957_),
    .A(_03945_),
    .B(_03956_));
 sg13g2_o21ai_1 _17538_ (.B1(_03900_),
    .Y(_03958_),
    .A1(_03907_),
    .A2(_03925_));
 sg13g2_nand2_1 _17539_ (.Y(_03959_),
    .A(_03926_),
    .B(_03958_));
 sg13g2_nor2_1 _17540_ (.A(_03957_),
    .B(_03959_),
    .Y(_03960_));
 sg13g2_xor2_1 _17541_ (.B(_03959_),
    .A(_03957_),
    .X(_03961_));
 sg13g2_inv_1 _17542_ (.Y(_03962_),
    .A(_03963_));
 sg13g2_o21ai_1 _17543_ (.B1(_03945_),
    .Y(_03963_),
    .A1(_03924_),
    .A2(_03954_));
 sg13g2_nor2_1 _17544_ (.A(net7226),
    .B(net7211),
    .Y(_03964_));
 sg13g2_nor2_1 _17545_ (.A(net7221),
    .B(net7217),
    .Y(_03965_));
 sg13g2_nor2_1 _17546_ (.A(net7229),
    .B(net7213),
    .Y(_03966_));
 sg13g2_xnor2_1 _17547_ (.Y(_03967_),
    .A(_03964_),
    .B(_03966_));
 sg13g2_xnor2_1 _17548_ (.Y(_03968_),
    .A(_03965_),
    .B(_03967_));
 sg13g2_nor2_1 _17549_ (.A(net7069),
    .B(net7205),
    .Y(_03969_));
 sg13g2_a22oi_1 _17550_ (.Y(_03970_),
    .B1(net7440),
    .B2(_14722_),
    .A2(net7638),
    .A1(net7339));
 sg13g2_inv_1 _17551_ (.Y(_03971_),
    .A(_03970_));
 sg13g2_o21ai_1 _17552_ (.B1(net7071),
    .Y(_03972_),
    .A1(_03950_),
    .A2(_03971_));
 sg13g2_nand2_1 _17553_ (.Y(_03973_),
    .A(_03969_),
    .B(_03972_));
 sg13g2_nor2_1 _17554_ (.A(net7205),
    .B(_03971_),
    .Y(_03974_));
 sg13g2_mux2_1 _17555_ (.A0(_03971_),
    .A1(_03974_),
    .S(_03950_),
    .X(_03975_));
 sg13g2_a21o_1 _17556_ (.A2(_03950_),
    .A1(_03836_),
    .B1(net7205),
    .X(_03976_));
 sg13g2_a22oi_1 _17557_ (.Y(_03977_),
    .B1(_03976_),
    .B2(_03971_),
    .A2(_03975_),
    .A1(net7070));
 sg13g2_o21ai_1 _17558_ (.B1(_03973_),
    .Y(_03978_),
    .A1(net7247),
    .A2(_03977_));
 sg13g2_xor2_1 _17559_ (.B(_03978_),
    .A(_03968_),
    .X(_03979_));
 sg13g2_nor2_1 _17560_ (.A(_03943_),
    .B(_03944_),
    .Y(_03980_));
 sg13g2_a22oi_1 _17561_ (.Y(_03981_),
    .B1(net7632),
    .B2(_15075_),
    .A2(net7635),
    .A1(_03017_));
 sg13g2_nor2_1 _17562_ (.A(net7246),
    .B(net7199),
    .Y(_03982_));
 sg13g2_a22oi_1 _17563_ (.Y(_03983_),
    .B1(net7319),
    .B2(_01639_),
    .A2(net7326),
    .A1(_01656_));
 sg13g2_o21ai_1 _17564_ (.B1(_03983_),
    .Y(_03984_),
    .A1(net7239),
    .A2(net7209));
 sg13g2_nor3_1 _17565_ (.A(net7235),
    .B(net7209),
    .C(_03983_),
    .Y(_03985_));
 sg13g2_or3_1 _17566_ (.A(net7239),
    .B(net7209),
    .C(_03983_),
    .X(_03986_));
 sg13g2_nand2_1 _17567_ (.Y(_03987_),
    .A(_03984_),
    .B(_03986_));
 sg13g2_xnor2_1 _17568_ (.Y(_03988_),
    .A(_03982_),
    .B(_03987_));
 sg13g2_a21oi_1 _17569_ (.A1(_03932_),
    .A2(_03935_),
    .Y(_03989_),
    .B1(_03934_));
 sg13g2_nand2_1 _17570_ (.Y(_03990_),
    .A(_03947_),
    .B(_03948_));
 sg13g2_o21ai_1 _17571_ (.B1(_03946_),
    .Y(_03991_),
    .A1(_03947_),
    .A2(_03948_));
 sg13g2_nand2_1 _17572_ (.Y(_03992_),
    .A(_03990_),
    .B(_03991_));
 sg13g2_xor2_1 _17573_ (.B(_03992_),
    .A(_03988_),
    .X(_03993_));
 sg13g2_xnor2_1 _17574_ (.Y(_03994_),
    .A(_03989_),
    .B(_03993_));
 sg13g2_a21oi_1 _17575_ (.A1(_03940_),
    .A2(_03941_),
    .Y(_03995_),
    .B1(_03937_));
 sg13g2_nor2_1 _17576_ (.A(_03940_),
    .B(_03941_),
    .Y(_03996_));
 sg13g2_nor2_1 _17577_ (.A(_03995_),
    .B(_03996_),
    .Y(_03997_));
 sg13g2_xnor2_1 _17578_ (.Y(_03998_),
    .A(_03994_),
    .B(_03997_));
 sg13g2_xor2_1 _17579_ (.B(_03998_),
    .A(_03980_),
    .X(_03999_));
 sg13g2_xnor2_1 _17580_ (.Y(_04000_),
    .A(_03979_),
    .B(_03999_));
 sg13g2_nor3_1 _17581_ (.A(_03955_),
    .B(_03962_),
    .C(_04000_),
    .Y(_04001_));
 sg13g2_o21ai_1 _17582_ (.B1(_04000_),
    .Y(_04002_),
    .A1(_03955_),
    .A2(_03962_));
 sg13g2_nor2b_1 _17583_ (.A(_04001_),
    .B_N(_04002_),
    .Y(_04003_));
 sg13g2_a21o_1 _17584_ (.A2(_03998_),
    .A1(_03980_),
    .B1(_03979_),
    .X(_04004_));
 sg13g2_o21ai_1 _17585_ (.B1(_04004_),
    .Y(_04005_),
    .A1(_03980_),
    .A2(_03998_));
 sg13g2_nor2_1 _17586_ (.A(net7247),
    .B(_03970_),
    .Y(_04006_));
 sg13g2_xor2_1 _17587_ (.B(_04006_),
    .A(_03969_),
    .X(_04007_));
 sg13g2_and2_1 _17588_ (.A(_03968_),
    .B(_04007_),
    .X(_04008_));
 sg13g2_nand2_1 _17589_ (.Y(_04009_),
    .A(_03968_),
    .B(_04007_));
 sg13g2_nor2_1 _17590_ (.A(net7225),
    .B(net7209),
    .Y(_04010_));
 sg13g2_nor2_1 _17591_ (.A(net7217),
    .B(net7211),
    .Y(_04011_));
 sg13g2_nor2_1 _17592_ (.A(net7221),
    .B(net7213),
    .Y(_04012_));
 sg13g2_xnor2_1 _17593_ (.Y(_04013_),
    .A(_04011_),
    .B(_04012_));
 sg13g2_xnor2_1 _17594_ (.Y(_04014_),
    .A(_04010_),
    .B(_04013_));
 sg13g2_a21oi_1 _17595_ (.A1(_03833_),
    .A2(net7241),
    .Y(_04015_),
    .B1(net7201));
 sg13g2_nor2_1 _17596_ (.A(net7230),
    .B(net7208),
    .Y(_04016_));
 sg13g2_and2_1 _17597_ (.A(net7068),
    .B(_04016_),
    .X(_04017_));
 sg13g2_nand2_1 _17598_ (.Y(_04018_),
    .A(net7068),
    .B(_04016_));
 sg13g2_and2_1 _17599_ (.A(net7272),
    .B(_03827_),
    .X(_04019_));
 sg13g2_and2_1 _17600_ (.A(net7337),
    .B(net7637),
    .X(_04020_));
 sg13g2_a22oi_1 _17601_ (.Y(_04021_),
    .B1(_03827_),
    .B2(_15458_),
    .A2(net7637),
    .A1(_03052_));
 sg13g2_inv_1 _17602_ (.Y(_04022_),
    .A(_04021_));
 sg13g2_and2_1 _17603_ (.A(net7208),
    .B(net7068),
    .X(_04023_));
 sg13g2_a21oi_1 _17604_ (.A1(net7207),
    .A2(net7068),
    .Y(_04024_),
    .B1(_04016_));
 sg13g2_nand2_1 _17605_ (.Y(_04025_),
    .A(_03826_),
    .B(_04022_));
 sg13g2_nor2_1 _17606_ (.A(_04024_),
    .B(_04025_),
    .Y(_04026_));
 sg13g2_nor3_1 _17607_ (.A(net7247),
    .B(net7208),
    .C(net7197),
    .Y(_04027_));
 sg13g2_a21o_1 _17608_ (.A2(net7068),
    .A1(net7247),
    .B1(_04027_),
    .X(_04028_));
 sg13g2_mux2_1 _17609_ (.A0(_04016_),
    .A1(net7208),
    .S(net7068),
    .X(_04029_));
 sg13g2_a22oi_1 _17610_ (.Y(_04030_),
    .B1(_04029_),
    .B2(net7247),
    .A2(_04028_),
    .A1(net7230));
 sg13g2_nand2b_1 _17611_ (.Y(_04031_),
    .B(net7205),
    .A_N(_04021_));
 sg13g2_or4_1 _17612_ (.A(net7229),
    .B(_03952_),
    .C(_04019_),
    .D(_04020_),
    .X(_04032_));
 sg13g2_o21ai_1 _17613_ (.B1(_04032_),
    .Y(_04033_),
    .A1(net7068),
    .A2(_04031_));
 sg13g2_a22oi_1 _17614_ (.Y(_04034_),
    .B1(_04033_),
    .B2(net7071),
    .A2(_04023_),
    .A1(net7197));
 sg13g2_nand3_1 _17615_ (.B(_04030_),
    .C(_04034_),
    .A(_04014_),
    .Y(_04035_));
 sg13g2_a21o_1 _17616_ (.A2(_04034_),
    .A1(_04030_),
    .B1(_04014_),
    .X(_04036_));
 sg13g2_nand2_1 _17617_ (.Y(_04037_),
    .A(_04035_),
    .B(_04036_));
 sg13g2_a21oi_1 _17618_ (.A1(_04035_),
    .A2(_04036_),
    .Y(_04038_),
    .B1(_04009_));
 sg13g2_a21o_1 _17619_ (.A2(_04036_),
    .A1(_04035_),
    .B1(_04009_),
    .X(_04039_));
 sg13g2_xnor2_1 _17620_ (.Y(_04040_),
    .A(_04008_),
    .B(_04037_));
 sg13g2_a22oi_1 _17621_ (.Y(_04041_),
    .B1(net7634),
    .B2(_15562_),
    .A2(net7636),
    .A1(_03084_));
 sg13g2_nor2_1 _17622_ (.A(net7244),
    .B(net7191),
    .Y(_04042_));
 sg13g2_a22oi_1 _17623_ (.Y(_04043_),
    .B1(_03819_),
    .B2(_01640_),
    .A2(_03817_),
    .A1(net7978));
 sg13g2_o21ai_1 _17624_ (.B1(_04043_),
    .Y(_04044_),
    .A1(net7235),
    .A2(net7198));
 sg13g2_nor3_1 _17625_ (.A(net7235),
    .B(net7198),
    .C(_04043_),
    .Y(_04045_));
 sg13g2_or3_1 _17626_ (.A(net7235),
    .B(net7198),
    .C(_04043_),
    .X(_04046_));
 sg13g2_nand2_1 _17627_ (.Y(_04047_),
    .A(_04044_),
    .B(_04046_));
 sg13g2_xnor2_1 _17628_ (.Y(_04048_),
    .A(_04042_),
    .B(_04047_));
 sg13g2_xor2_1 _17629_ (.B(_04047_),
    .A(_04042_),
    .X(_04049_));
 sg13g2_a21o_1 _17630_ (.A2(_03984_),
    .A1(_03982_),
    .B1(_03985_),
    .X(_04050_));
 sg13g2_a21oi_1 _17631_ (.A1(_03982_),
    .A2(_03984_),
    .Y(_04051_),
    .B1(_03985_));
 sg13g2_nand2_1 _17632_ (.Y(_04052_),
    .A(_03964_),
    .B(_03965_));
 sg13g2_o21ai_1 _17633_ (.B1(_03966_),
    .Y(_04053_),
    .A1(_03964_),
    .A2(_03965_));
 sg13g2_a21oi_1 _17634_ (.A1(_04052_),
    .A2(_04053_),
    .Y(_04054_),
    .B1(_04050_));
 sg13g2_a21o_1 _17635_ (.A2(_04053_),
    .A1(_04052_),
    .B1(_04050_),
    .X(_04055_));
 sg13g2_and3_1 _17636_ (.X(_04056_),
    .A(_04050_),
    .B(_04052_),
    .C(_04053_));
 sg13g2_nand3_1 _17637_ (.B(_04052_),
    .C(_04053_),
    .A(_04050_),
    .Y(_04057_));
 sg13g2_nor3_1 _17638_ (.A(_04049_),
    .B(_04054_),
    .C(_04056_),
    .Y(_04058_));
 sg13g2_nand3_1 _17639_ (.B(_04055_),
    .C(_04057_),
    .A(_04048_),
    .Y(_04059_));
 sg13g2_a21oi_1 _17640_ (.A1(_04055_),
    .A2(_04057_),
    .Y(_04060_),
    .B1(_04048_));
 sg13g2_o21ai_1 _17641_ (.B1(_04049_),
    .Y(_04061_),
    .A1(_04054_),
    .A2(_04056_));
 sg13g2_nand3_1 _17642_ (.B(_03990_),
    .C(_03991_),
    .A(_03989_),
    .Y(_04062_));
 sg13g2_a21oi_1 _17643_ (.A1(_03990_),
    .A2(_03991_),
    .Y(_04063_),
    .B1(_03989_));
 sg13g2_a21oi_1 _17644_ (.A1(_03988_),
    .A2(_04062_),
    .Y(_04064_),
    .B1(_04063_));
 sg13g2_nor3_1 _17645_ (.A(_04058_),
    .B(_04060_),
    .C(_04064_),
    .Y(_04065_));
 sg13g2_o21ai_1 _17646_ (.B1(_04064_),
    .Y(_04066_),
    .A1(_04058_),
    .A2(_04060_));
 sg13g2_nand2b_1 _17647_ (.Y(_04067_),
    .B(_04066_),
    .A_N(_04065_));
 sg13g2_xnor2_1 _17648_ (.Y(_04068_),
    .A(net7069),
    .B(net7201));
 sg13g2_xnor2_1 _17649_ (.Y(_04069_),
    .A(_03968_),
    .B(_04068_));
 sg13g2_nand3_1 _17650_ (.B(_03953_),
    .C(_04069_),
    .A(_03950_),
    .Y(_04070_));
 sg13g2_nand2b_1 _17651_ (.Y(_04071_),
    .B(_03994_),
    .A_N(_03997_));
 sg13g2_xor2_1 _17652_ (.B(_04071_),
    .A(_04067_),
    .X(_04072_));
 sg13g2_xnor2_1 _17653_ (.Y(_04073_),
    .A(_04070_),
    .B(_04072_));
 sg13g2_or2_1 _17654_ (.X(_04074_),
    .B(_04073_),
    .A(_04040_));
 sg13g2_xnor2_1 _17655_ (.Y(_04075_),
    .A(_04040_),
    .B(_04073_));
 sg13g2_nor2_1 _17656_ (.A(_04005_),
    .B(_04075_),
    .Y(_04076_));
 sg13g2_xor2_1 _17657_ (.B(_04075_),
    .A(_04005_),
    .X(_04077_));
 sg13g2_a22oi_1 _17658_ (.Y(_04078_),
    .B1(net7632),
    .B2(_02066_),
    .A2(net7635),
    .A1(_03159_));
 sg13g2_nor2_1 _17659_ (.A(net7244),
    .B(net7188),
    .Y(_04079_));
 sg13g2_a22oi_1 _17660_ (.Y(_04080_),
    .B1(_03819_),
    .B2(_01641_),
    .A2(_03817_),
    .A1(_01658_));
 sg13g2_nor3_1 _17661_ (.A(net7235),
    .B(net7191),
    .C(_04080_),
    .Y(_04081_));
 sg13g2_o21ai_1 _17662_ (.B1(_04080_),
    .Y(_04082_),
    .A1(net7235),
    .A2(net7191));
 sg13g2_nand2b_1 _17663_ (.Y(_04083_),
    .B(_04082_),
    .A_N(_04081_));
 sg13g2_xnor2_1 _17664_ (.Y(_04084_),
    .A(_04079_),
    .B(_04083_));
 sg13g2_a21oi_1 _17665_ (.A1(_04042_),
    .A2(_04044_),
    .Y(_04085_),
    .B1(_04045_));
 sg13g2_a21oi_1 _17666_ (.A1(_04010_),
    .A2(_04011_),
    .Y(_04086_),
    .B1(_04012_));
 sg13g2_a21o_1 _17667_ (.A2(_04011_),
    .A1(_04010_),
    .B1(_04012_),
    .X(_04087_));
 sg13g2_nor2_1 _17668_ (.A(_04010_),
    .B(_04011_),
    .Y(_04088_));
 sg13g2_or2_1 _17669_ (.X(_04089_),
    .B(_04011_),
    .A(_04010_));
 sg13g2_nand3_1 _17670_ (.B(_04087_),
    .C(_04089_),
    .A(_04085_),
    .Y(_04090_));
 sg13g2_a21o_1 _17671_ (.A2(_04089_),
    .A1(_04087_),
    .B1(_04085_),
    .X(_04091_));
 sg13g2_and3_1 _17672_ (.X(_04092_),
    .A(_04084_),
    .B(_04090_),
    .C(_04091_));
 sg13g2_a21oi_1 _17673_ (.A1(_04090_),
    .A2(_04091_),
    .Y(_04093_),
    .B1(_04084_));
 sg13g2_or2_1 _17674_ (.X(_04094_),
    .B(_04093_),
    .A(_04092_));
 sg13g2_and3_1 _17675_ (.X(_04095_),
    .A(_04051_),
    .B(_04052_),
    .C(_04053_));
 sg13g2_a21o_1 _17676_ (.A2(_04053_),
    .A1(_04052_),
    .B1(_04051_),
    .X(_04096_));
 sg13g2_a21oi_1 _17677_ (.A1(_04049_),
    .A2(_04096_),
    .Y(_04097_),
    .B1(_04095_));
 sg13g2_o21ai_1 _17678_ (.B1(_04097_),
    .Y(_04098_),
    .A1(_04092_),
    .A2(_04093_));
 sg13g2_xnor2_1 _17679_ (.Y(_04099_),
    .A(_04094_),
    .B(_04097_));
 sg13g2_a21oi_1 _17680_ (.A1(_04059_),
    .A2(_04061_),
    .Y(_04100_),
    .B1(_04064_));
 sg13g2_xnor2_1 _17681_ (.Y(_04101_),
    .A(_04039_),
    .B(_04100_));
 sg13g2_nand2b_1 _17682_ (.Y(_04102_),
    .B(_04099_),
    .A_N(_04100_));
 sg13g2_nor2b_1 _17683_ (.A(_04099_),
    .B_N(_04100_),
    .Y(_04103_));
 sg13g2_xor2_1 _17684_ (.B(_04101_),
    .A(_04099_),
    .X(_04104_));
 sg13g2_nor2_1 _17685_ (.A(_04015_),
    .B(_04016_),
    .Y(_04105_));
 sg13g2_a221oi_1 _17686_ (.B2(_04105_),
    .C1(_04026_),
    .B1(_04025_),
    .A1(net7247),
    .Y(_04106_),
    .A2(_04017_));
 sg13g2_nor2_1 _17687_ (.A(net7230),
    .B(net7195),
    .Y(_04107_));
 sg13g2_xnor2_1 _17688_ (.Y(_04108_),
    .A(net7230),
    .B(net7195));
 sg13g2_and2_1 _17689_ (.A(net7068),
    .B(_04108_),
    .X(_04109_));
 sg13g2_a22oi_1 _17690_ (.Y(_04110_),
    .B1(_04109_),
    .B2(_03953_),
    .A2(_04106_),
    .A1(_04014_));
 sg13g2_nor2_1 _17691_ (.A(net7225),
    .B(net7198),
    .Y(_04111_));
 sg13g2_nor2_1 _17692_ (.A(net7217),
    .B(net7209),
    .Y(_04112_));
 sg13g2_nor2_1 _17693_ (.A(net7213),
    .B(net7211),
    .Y(_04113_));
 sg13g2_xnor2_1 _17694_ (.Y(_04114_),
    .A(_04112_),
    .B(_04113_));
 sg13g2_xnor2_1 _17695_ (.Y(_04115_),
    .A(_04111_),
    .B(_04114_));
 sg13g2_o21ai_1 _17696_ (.B1(_04018_),
    .Y(_04116_),
    .A1(_04025_),
    .A2(_04105_));
 sg13g2_nand2_1 _17697_ (.Y(_04117_),
    .A(_03836_),
    .B(_04022_));
 sg13g2_nor2_1 _17698_ (.A(net7224),
    .B(_03952_),
    .Y(_04118_));
 sg13g2_nor2_1 _17699_ (.A(net7230),
    .B(net7201),
    .Y(_04119_));
 sg13g2_xor2_1 _17700_ (.B(_04119_),
    .A(_04118_),
    .X(_04120_));
 sg13g2_xnor2_1 _17701_ (.Y(_04121_),
    .A(_04117_),
    .B(_04120_));
 sg13g2_nor2_1 _17702_ (.A(_04116_),
    .B(_04121_),
    .Y(_04122_));
 sg13g2_xor2_1 _17703_ (.B(_04121_),
    .A(_04116_),
    .X(_04123_));
 sg13g2_xnor2_1 _17704_ (.Y(_04124_),
    .A(_04115_),
    .B(_04123_));
 sg13g2_nor2_1 _17705_ (.A(_04110_),
    .B(_04124_),
    .Y(_04125_));
 sg13g2_or2_1 _17706_ (.X(_04126_),
    .B(_04124_),
    .A(_04110_));
 sg13g2_xnor2_1 _17707_ (.Y(_04127_),
    .A(_04110_),
    .B(_04124_));
 sg13g2_and4_1 _17708_ (.A(_02015_),
    .B(_02018_),
    .C(_02028_),
    .D(net7441),
    .X(_04128_));
 sg13g2_a22oi_1 _17709_ (.Y(_04129_),
    .B1(_04128_),
    .B2(_02012_),
    .A2(net7639),
    .A1(_03121_));
 sg13g2_inv_1 _17710_ (.Y(_04130_),
    .A(net7185));
 sg13g2_nor2_1 _17711_ (.A(net7249),
    .B(net7187),
    .Y(_04131_));
 sg13g2_nor2b_1 _17712_ (.A(_04127_),
    .B_N(net7066),
    .Y(_04132_));
 sg13g2_xnor2_1 _17713_ (.Y(_04133_),
    .A(_04127_),
    .B(net7066));
 sg13g2_xnor2_1 _17714_ (.Y(_04134_),
    .A(_04104_),
    .B(_04133_));
 sg13g2_nor2b_1 _17715_ (.A(_04067_),
    .B_N(_04070_),
    .Y(_04135_));
 sg13g2_nand2b_1 _17716_ (.Y(_04136_),
    .B(_04067_),
    .A_N(_04070_));
 sg13g2_o21ai_1 _17717_ (.B1(_04136_),
    .Y(_04137_),
    .A1(_04071_),
    .A2(_04135_));
 sg13g2_nor2_1 _17718_ (.A(_04134_),
    .B(_04137_),
    .Y(_04138_));
 sg13g2_nand2_1 _17719_ (.Y(_04139_),
    .A(_04134_),
    .B(_04137_));
 sg13g2_nand2b_1 _17720_ (.Y(_04140_),
    .B(_04139_),
    .A_N(_04138_));
 sg13g2_xor2_1 _17721_ (.B(_04140_),
    .A(_04074_),
    .X(_04141_));
 sg13g2_a22oi_1 _17722_ (.Y(_04142_),
    .B1(net7633),
    .B2(_02141_),
    .A2(net7635),
    .A1(_03225_));
 sg13g2_nor2_1 _17723_ (.A(net7244),
    .B(_04142_),
    .Y(_04143_));
 sg13g2_a22oi_1 _17724_ (.Y(_04144_),
    .B1(net7324),
    .B2(_01642_),
    .A2(_03817_),
    .A1(_01659_));
 sg13g2_nor3_1 _17725_ (.A(net7236),
    .B(net7188),
    .C(_04144_),
    .Y(_04145_));
 sg13g2_o21ai_1 _17726_ (.B1(_04144_),
    .Y(_04146_),
    .A1(net7236),
    .A2(net7188));
 sg13g2_nand2b_1 _17727_ (.Y(_04147_),
    .B(_04146_),
    .A_N(_04145_));
 sg13g2_xnor2_1 _17728_ (.Y(_04148_),
    .A(_04143_),
    .B(_04147_));
 sg13g2_a21oi_1 _17729_ (.A1(_04079_),
    .A2(_04082_),
    .Y(_04149_),
    .B1(_04081_));
 sg13g2_a21oi_1 _17730_ (.A1(_04111_),
    .A2(_04112_),
    .Y(_04150_),
    .B1(_04113_));
 sg13g2_a21o_1 _17731_ (.A2(_04112_),
    .A1(_04111_),
    .B1(_04113_),
    .X(_04151_));
 sg13g2_nor2_1 _17732_ (.A(_04111_),
    .B(_04112_),
    .Y(_04152_));
 sg13g2_or2_1 _17733_ (.X(_04153_),
    .B(_04112_),
    .A(_04111_));
 sg13g2_nand3_1 _17734_ (.B(_04151_),
    .C(_04153_),
    .A(_04149_),
    .Y(_04154_));
 sg13g2_a21o_1 _17735_ (.A2(_04153_),
    .A1(_04151_),
    .B1(_04149_),
    .X(_04155_));
 sg13g2_nand3_1 _17736_ (.B(_04154_),
    .C(_04155_),
    .A(_04148_),
    .Y(_04156_));
 sg13g2_a21o_1 _17737_ (.A2(_04155_),
    .A1(_04154_),
    .B1(_04148_),
    .X(_04157_));
 sg13g2_o21ai_1 _17738_ (.B1(_04085_),
    .Y(_04158_),
    .A1(_04086_),
    .A2(_04088_));
 sg13g2_nor3_1 _17739_ (.A(_04085_),
    .B(_04086_),
    .C(_04088_),
    .Y(_04159_));
 sg13g2_o21ai_1 _17740_ (.B1(_04158_),
    .Y(_04160_),
    .A1(_04084_),
    .A2(_04159_));
 sg13g2_a21oi_1 _17741_ (.A1(_04156_),
    .A2(_04157_),
    .Y(_04161_),
    .B1(_04160_));
 sg13g2_a21o_1 _17742_ (.A2(_04157_),
    .A1(_04156_),
    .B1(_04160_),
    .X(_04162_));
 sg13g2_and3_1 _17743_ (.X(_04163_),
    .A(_04156_),
    .B(_04157_),
    .C(_04160_));
 sg13g2_nand3_1 _17744_ (.B(_04157_),
    .C(_04160_),
    .A(_04156_),
    .Y(_04164_));
 sg13g2_nand2_1 _17745_ (.Y(_04165_),
    .A(_04162_),
    .B(_04164_));
 sg13g2_nor3_1 _17746_ (.A(_04098_),
    .B(_04161_),
    .C(_04163_),
    .Y(_04166_));
 sg13g2_nand4_1 _17747_ (.B(_04097_),
    .C(_04162_),
    .A(_04094_),
    .Y(_04167_),
    .D(_04164_));
 sg13g2_a22oi_1 _17748_ (.Y(_04168_),
    .B1(_04162_),
    .B2(_04164_),
    .A2(_04097_),
    .A1(_04094_));
 sg13g2_o21ai_1 _17749_ (.B1(_04098_),
    .Y(_04169_),
    .A1(_04161_),
    .A2(_04163_));
 sg13g2_nor3_1 _17750_ (.A(_04126_),
    .B(_04166_),
    .C(_04168_),
    .Y(_04170_));
 sg13g2_nand3_1 _17751_ (.B(_04167_),
    .C(_04169_),
    .A(_04125_),
    .Y(_04171_));
 sg13g2_a21oi_1 _17752_ (.A1(_04167_),
    .A2(_04169_),
    .Y(_04172_),
    .B1(_04125_));
 sg13g2_o21ai_1 _17753_ (.B1(_04126_),
    .Y(_04173_),
    .A1(_04166_),
    .A2(_04168_));
 sg13g2_nand2_1 _17754_ (.Y(_04174_),
    .A(_04171_),
    .B(_04173_));
 sg13g2_nand2b_1 _17755_ (.Y(_04175_),
    .B(net7441),
    .A_N(_02088_));
 sg13g2_nor3_1 _17756_ (.A(_02091_),
    .B(_02101_),
    .C(_04175_),
    .Y(_04176_));
 sg13g2_and3_1 _17757_ (.X(_04177_),
    .A(_03174_),
    .B(_03179_),
    .C(net7639));
 sg13g2_a22oi_1 _17758_ (.Y(_04178_),
    .B1(_04177_),
    .B2(_03190_),
    .A2(_04176_),
    .A1(_02086_));
 sg13g2_nor2_1 _17759_ (.A(net7249),
    .B(_04178_),
    .Y(_04179_));
 sg13g2_nor2_1 _17760_ (.A(net7070),
    .B(net7187),
    .Y(_04180_));
 sg13g2_xnor2_1 _17761_ (.Y(_04181_),
    .A(_04179_),
    .B(_04180_));
 sg13g2_nor2_1 _17762_ (.A(net7211),
    .B(net7204),
    .Y(_04182_));
 sg13g2_nor2_1 _17763_ (.A(net7224),
    .B(net7201),
    .Y(_04183_));
 sg13g2_xnor2_1 _17764_ (.Y(_04184_),
    .A(_04182_),
    .B(_04183_));
 sg13g2_xnor2_1 _17765_ (.Y(_04185_),
    .A(_04107_),
    .B(_04184_));
 sg13g2_nand2_1 _17766_ (.Y(_04186_),
    .A(_04118_),
    .B(_04119_));
 sg13g2_nor2_1 _17767_ (.A(_04118_),
    .B(_04119_),
    .Y(_04187_));
 sg13g2_o21ai_1 _17768_ (.B1(_04186_),
    .Y(_04188_),
    .A1(_04117_),
    .A2(_04187_));
 sg13g2_nor2_1 _17769_ (.A(net7225),
    .B(net7194),
    .Y(_04189_));
 sg13g2_nor2_1 _17770_ (.A(net7217),
    .B(net7199),
    .Y(_04190_));
 sg13g2_nor2_1 _17771_ (.A(net7214),
    .B(net7209),
    .Y(_04191_));
 sg13g2_xnor2_1 _17772_ (.Y(_04192_),
    .A(_04189_),
    .B(_04191_));
 sg13g2_xnor2_1 _17773_ (.Y(_04193_),
    .A(_04190_),
    .B(_04192_));
 sg13g2_nor2_1 _17774_ (.A(_04188_),
    .B(_04193_),
    .Y(_04194_));
 sg13g2_xnor2_1 _17775_ (.Y(_04195_),
    .A(_04188_),
    .B(_04193_));
 sg13g2_xnor2_1 _17776_ (.Y(_04196_),
    .A(_04185_),
    .B(_04195_));
 sg13g2_a21oi_1 _17777_ (.A1(_04116_),
    .A2(_04121_),
    .Y(_04197_),
    .B1(_04115_));
 sg13g2_nor2_1 _17778_ (.A(_04122_),
    .B(_04197_),
    .Y(_04198_));
 sg13g2_xnor2_1 _17779_ (.Y(_04199_),
    .A(_04196_),
    .B(_04198_));
 sg13g2_or2_1 _17780_ (.X(_04200_),
    .B(_04199_),
    .A(_04181_));
 sg13g2_xnor2_1 _17781_ (.Y(_04201_),
    .A(_04181_),
    .B(_04199_));
 sg13g2_xor2_1 _17782_ (.B(_04199_),
    .A(_04181_),
    .X(_04202_));
 sg13g2_nor2_1 _17783_ (.A(_04132_),
    .B(_04202_),
    .Y(_04203_));
 sg13g2_xnor2_1 _17784_ (.Y(_04204_),
    .A(_04132_),
    .B(_04202_));
 sg13g2_xnor2_1 _17785_ (.Y(_04205_),
    .A(_04174_),
    .B(_04204_));
 sg13g2_nand2b_1 _17786_ (.Y(_04206_),
    .B(_04133_),
    .A_N(_04104_));
 sg13g2_o21ai_1 _17787_ (.B1(_04102_),
    .Y(_04207_),
    .A1(_04038_),
    .A2(_04103_));
 sg13g2_and2_1 _17788_ (.A(_04206_),
    .B(_04207_),
    .X(_04208_));
 sg13g2_or2_1 _17789_ (.X(_04209_),
    .B(_04207_),
    .A(_04206_));
 sg13g2_nand2b_1 _17790_ (.Y(_04210_),
    .B(_04209_),
    .A_N(_04208_));
 sg13g2_xor2_1 _17791_ (.B(_04210_),
    .A(_04205_),
    .X(_04211_));
 sg13g2_o21ai_1 _17792_ (.B1(_04149_),
    .Y(_04212_),
    .A1(_04150_),
    .A2(_04152_));
 sg13g2_nor3_1 _17793_ (.A(_04149_),
    .B(_04150_),
    .C(_04152_),
    .Y(_04213_));
 sg13g2_o21ai_1 _17794_ (.B1(_04212_),
    .Y(_04214_),
    .A1(_04148_),
    .A2(_04213_));
 sg13g2_a22oi_1 _17795_ (.Y(_04215_),
    .B1(_03823_),
    .B2(_02205_),
    .A2(_03822_),
    .A1(_03293_));
 sg13g2_nor2_1 _17796_ (.A(net7244),
    .B(net7173),
    .Y(_04216_));
 sg13g2_a22oi_1 _17797_ (.Y(_04217_),
    .B1(net7324),
    .B2(_01643_),
    .A2(_03817_),
    .A1(_01661_));
 sg13g2_nor3_1 _17798_ (.A(net7236),
    .B(_04142_),
    .C(_04217_),
    .Y(_04218_));
 sg13g2_o21ai_1 _17799_ (.B1(_04217_),
    .Y(_04219_),
    .A1(net7236),
    .A2(_04142_));
 sg13g2_nand2b_1 _17800_ (.Y(_04220_),
    .B(_04219_),
    .A_N(_04218_));
 sg13g2_xnor2_1 _17801_ (.Y(_04221_),
    .A(_04216_),
    .B(_04220_));
 sg13g2_a21o_1 _17802_ (.A2(_04146_),
    .A1(_04143_),
    .B1(_04145_),
    .X(_04222_));
 sg13g2_nand2_1 _17803_ (.Y(_04223_),
    .A(_04190_),
    .B(_04191_));
 sg13g2_o21ai_1 _17804_ (.B1(_04189_),
    .Y(_04224_),
    .A1(_04190_),
    .A2(_04191_));
 sg13g2_nand2_1 _17805_ (.Y(_04225_),
    .A(_04223_),
    .B(_04224_));
 sg13g2_a21o_1 _17806_ (.A2(_04224_),
    .A1(_04223_),
    .B1(_04222_),
    .X(_04226_));
 sg13g2_nand3_1 _17807_ (.B(_04223_),
    .C(_04224_),
    .A(_04222_),
    .Y(_04227_));
 sg13g2_nand3_1 _17808_ (.B(_04226_),
    .C(_04227_),
    .A(_04221_),
    .Y(_04228_));
 sg13g2_a21o_1 _17809_ (.A2(_04227_),
    .A1(_04226_),
    .B1(_04221_),
    .X(_04229_));
 sg13g2_nand3_1 _17810_ (.B(_04228_),
    .C(_04229_),
    .A(_04214_),
    .Y(_04230_));
 sg13g2_a21o_1 _17811_ (.A2(_04229_),
    .A1(_04228_),
    .B1(_04214_),
    .X(_04231_));
 sg13g2_and4_1 _17812_ (.A(_04196_),
    .B(_04198_),
    .C(_04230_),
    .D(_04231_),
    .X(_04232_));
 sg13g2_nand4_1 _17813_ (.B(_04198_),
    .C(_04230_),
    .A(_04196_),
    .Y(_04233_),
    .D(_04231_));
 sg13g2_a22oi_1 _17814_ (.Y(_04234_),
    .B1(_04230_),
    .B2(_04231_),
    .A2(_04198_),
    .A1(_04196_));
 sg13g2_nand3b_1 _17815_ (.B(_04161_),
    .C(_04233_),
    .Y(_04235_),
    .A_N(_04234_));
 sg13g2_o21ai_1 _17816_ (.B1(_04162_),
    .Y(_04236_),
    .A1(_04232_),
    .A2(_04234_));
 sg13g2_nand2_1 _17817_ (.Y(_04237_),
    .A(_04235_),
    .B(_04236_));
 sg13g2_a21oi_1 _17818_ (.A1(_03833_),
    .A2(_03834_),
    .Y(_04238_),
    .B1(_04178_));
 sg13g2_or2_1 _17819_ (.X(_04239_),
    .B(_04178_),
    .A(_03835_));
 sg13g2_nor2_1 _17820_ (.A(net7232),
    .B(net7187),
    .Y(_04240_));
 sg13g2_and4_1 _17821_ (.A(_02159_),
    .B(_02161_),
    .C(_02170_),
    .D(net7441),
    .X(_04241_));
 sg13g2_and3_1 _17822_ (.X(_04242_),
    .A(_03239_),
    .B(_03244_),
    .C(net7639));
 sg13g2_a22oi_1 _17823_ (.Y(_04243_),
    .B1(_04242_),
    .B2(_03255_),
    .A2(_04241_),
    .A1(_02157_));
 sg13g2_nand3_1 _17824_ (.B(_04239_),
    .C(net7167),
    .A(net7187),
    .Y(_04244_));
 sg13g2_a21oi_1 _17825_ (.A1(net7187),
    .A2(_04238_),
    .Y(_04245_),
    .B1(_04240_));
 sg13g2_or3_1 _17826_ (.A(net7249),
    .B(net7167),
    .C(_04245_),
    .X(_04246_));
 sg13g2_nand3_1 _17827_ (.B(net7067),
    .C(net7167),
    .A(net7071),
    .Y(_04247_));
 sg13g2_o21ai_1 _17828_ (.B1(_04247_),
    .Y(_04248_),
    .A1(net7071),
    .A2(_04238_));
 sg13g2_inv_1 _17829_ (.Y(_04249_),
    .A(_04250_));
 sg13g2_nand2_1 _17830_ (.Y(_04250_),
    .A(_04238_),
    .B(_04240_));
 sg13g2_o21ai_1 _17831_ (.B1(_04250_),
    .Y(_04251_),
    .A1(net7067),
    .A2(_04238_));
 sg13g2_a22oi_1 _17832_ (.Y(_04252_),
    .B1(_04251_),
    .B2(net7249),
    .A2(_04248_),
    .A1(net7232));
 sg13g2_nand3_1 _17833_ (.B(_04246_),
    .C(_04252_),
    .A(_04244_),
    .Y(_04253_));
 sg13g2_a21oi_1 _17834_ (.A1(_04188_),
    .A2(_04193_),
    .Y(_04254_),
    .B1(_04185_));
 sg13g2_nor2_1 _17835_ (.A(_04194_),
    .B(_04254_),
    .Y(_04255_));
 sg13g2_nor2_1 _17836_ (.A(net7225),
    .B(net7188),
    .Y(_04256_));
 sg13g2_nor2_1 _17837_ (.A(net7218),
    .B(net7194),
    .Y(_04257_));
 sg13g2_nor2_1 _17838_ (.A(net7214),
    .B(net7199),
    .Y(_04258_));
 sg13g2_xnor2_1 _17839_ (.Y(_04259_),
    .A(_04257_),
    .B(_04258_));
 sg13g2_xnor2_1 _17840_ (.Y(_04260_),
    .A(_04256_),
    .B(_04259_));
 sg13g2_nor2_1 _17841_ (.A(_04182_),
    .B(_04183_),
    .Y(_04261_));
 sg13g2_a21oi_1 _17842_ (.A1(_04182_),
    .A2(_04183_),
    .Y(_04262_),
    .B1(_04107_));
 sg13g2_nor2_1 _17843_ (.A(_04261_),
    .B(_04262_),
    .Y(_04263_));
 sg13g2_nor2_1 _17844_ (.A(net7224),
    .B(net7195),
    .Y(_04264_));
 sg13g2_nor2_1 _17845_ (.A(net7209),
    .B(net7204),
    .Y(_04265_));
 sg13g2_nor2_1 _17846_ (.A(net7211),
    .B(net7201),
    .Y(_04266_));
 sg13g2_xnor2_1 _17847_ (.Y(_04267_),
    .A(_04264_),
    .B(_04266_));
 sg13g2_xnor2_1 _17848_ (.Y(_04268_),
    .A(_04265_),
    .B(_04267_));
 sg13g2_nand2_1 _17849_ (.Y(_04269_),
    .A(_04263_),
    .B(_04268_));
 sg13g2_xor2_1 _17850_ (.B(_04268_),
    .A(_04263_),
    .X(_04270_));
 sg13g2_xnor2_1 _17851_ (.Y(_04271_),
    .A(_04260_),
    .B(_04270_));
 sg13g2_xnor2_1 _17852_ (.Y(_04272_),
    .A(_04255_),
    .B(_04271_));
 sg13g2_nor2b_1 _17853_ (.A(_04253_),
    .B_N(_04272_),
    .Y(_04273_));
 sg13g2_inv_1 _17854_ (.Y(_04274_),
    .A(_04273_));
 sg13g2_xnor2_1 _17855_ (.Y(_04275_),
    .A(_04253_),
    .B(_04272_));
 sg13g2_xnor2_1 _17856_ (.Y(_04276_),
    .A(_04200_),
    .B(_04275_));
 sg13g2_xor2_1 _17857_ (.B(_04276_),
    .A(_04237_),
    .X(_04277_));
 sg13g2_a22oi_1 _17858_ (.Y(_04278_),
    .B1(_04202_),
    .B2(_04132_),
    .A2(_04173_),
    .A1(_04171_));
 sg13g2_o21ai_1 _17859_ (.B1(_04201_),
    .Y(_04279_),
    .A1(_04170_),
    .A2(_04172_));
 sg13g2_nor3_1 _17860_ (.A(_04170_),
    .B(_04172_),
    .C(_04201_),
    .Y(_04280_));
 sg13g2_o21ai_1 _17861_ (.B1(_04098_),
    .Y(_04281_),
    .A1(_04126_),
    .A2(_04165_));
 sg13g2_nand2_1 _17862_ (.Y(_04282_),
    .A(_04126_),
    .B(_04165_));
 sg13g2_nand2_1 _17863_ (.Y(_04283_),
    .A(_04281_),
    .B(_04282_));
 sg13g2_or3_1 _17864_ (.A(_04203_),
    .B(_04278_),
    .C(_04283_),
    .X(_04284_));
 sg13g2_a221oi_1 _17865_ (.B2(_04282_),
    .C1(_04280_),
    .B1(_04281_),
    .A1(_04132_),
    .Y(_04285_),
    .A2(_04279_));
 sg13g2_o21ai_1 _17866_ (.B1(_04283_),
    .Y(_04286_),
    .A1(_04203_),
    .A2(_04278_));
 sg13g2_nand2_1 _17867_ (.Y(_04287_),
    .A(_04284_),
    .B(_04286_));
 sg13g2_xor2_1 _17868_ (.B(_04287_),
    .A(_04277_),
    .X(_04288_));
 sg13g2_nor2_1 _17869_ (.A(_03835_),
    .B(net7168),
    .Y(_04289_));
 sg13g2_nor2_1 _17870_ (.A(net7232),
    .B(_04178_),
    .Y(_04290_));
 sg13g2_nor2_1 _17871_ (.A(net7224),
    .B(net7184),
    .Y(_04291_));
 sg13g2_xnor2_1 _17872_ (.Y(_04292_),
    .A(_04290_),
    .B(_04291_));
 sg13g2_inv_1 _17873_ (.Y(_04293_),
    .A(_04294_));
 sg13g2_xnor2_1 _17874_ (.Y(_04294_),
    .A(_04289_),
    .B(_04292_));
 sg13g2_and4_1 _17875_ (.A(_02237_),
    .B(_02240_),
    .C(_02250_),
    .D(net7441),
    .X(_04295_));
 sg13g2_and3_1 _17876_ (.X(_04296_),
    .A(_03310_),
    .B(_03315_),
    .C(_03815_));
 sg13g2_a22oi_1 _17877_ (.Y(_04297_),
    .B1(_04296_),
    .B2(_03326_),
    .A2(_04295_),
    .A1(_02234_));
 sg13g2_nor2_1 _17878_ (.A(_04238_),
    .B(_04240_),
    .Y(_04298_));
 sg13g2_nor2_1 _17879_ (.A(net7168),
    .B(_04298_),
    .Y(_04299_));
 sg13g2_nor2_1 _17880_ (.A(_04239_),
    .B(net7168),
    .Y(_04300_));
 sg13g2_nand2_1 _17881_ (.Y(_04301_),
    .A(_04239_),
    .B(net7168));
 sg13g2_o21ai_1 _17882_ (.B1(_04301_),
    .Y(_04302_),
    .A1(_04240_),
    .A2(_04300_));
 sg13g2_mux2_1 _17883_ (.A0(_04302_),
    .A1(_04299_),
    .S(net7162),
    .X(_04303_));
 sg13g2_or2_1 _17884_ (.X(_04304_),
    .B(_04297_),
    .A(_03825_));
 sg13g2_a22oi_1 _17885_ (.Y(_04305_),
    .B1(_04304_),
    .B2(_04249_),
    .A2(_04303_),
    .A1(net7071));
 sg13g2_xnor2_1 _17886_ (.Y(_04306_),
    .A(net6947),
    .B(_04305_));
 sg13g2_nor2_1 _17887_ (.A(net7225),
    .B(net7183),
    .Y(_04307_));
 sg13g2_nor2_1 _17888_ (.A(net7218),
    .B(net7188),
    .Y(_04308_));
 sg13g2_nor2_1 _17889_ (.A(net7214),
    .B(net7194),
    .Y(_04309_));
 sg13g2_xnor2_1 _17890_ (.Y(_04310_),
    .A(_04308_),
    .B(_04309_));
 sg13g2_xnor2_1 _17891_ (.Y(_04311_),
    .A(_04307_),
    .B(_04310_));
 sg13g2_nor2_1 _17892_ (.A(_04265_),
    .B(_04266_),
    .Y(_04312_));
 sg13g2_a21oi_1 _17893_ (.A1(_04265_),
    .A2(_04266_),
    .Y(_04313_),
    .B1(_04264_));
 sg13g2_nor2_1 _17894_ (.A(_04312_),
    .B(_04313_),
    .Y(_04314_));
 sg13g2_nor2_1 _17895_ (.A(_03908_),
    .B(net7195),
    .Y(_04315_));
 sg13g2_nor2_1 _17896_ (.A(net7204),
    .B(net7199),
    .Y(_04316_));
 sg13g2_nor2_1 _17897_ (.A(_03931_),
    .B(net7201),
    .Y(_04317_));
 sg13g2_xnor2_1 _17898_ (.Y(_04318_),
    .A(_04315_),
    .B(_04317_));
 sg13g2_xnor2_1 _17899_ (.Y(_04319_),
    .A(_04316_),
    .B(_04318_));
 sg13g2_nor2_1 _17900_ (.A(_04314_),
    .B(_04319_),
    .Y(_04320_));
 sg13g2_xor2_1 _17901_ (.B(_04319_),
    .A(_04314_),
    .X(_04321_));
 sg13g2_xnor2_1 _17902_ (.Y(_04322_),
    .A(_04311_),
    .B(_04321_));
 sg13g2_o21ai_1 _17903_ (.B1(_04260_),
    .Y(_04323_),
    .A1(_04263_),
    .A2(_04268_));
 sg13g2_nor2_1 _17904_ (.A(_03846_),
    .B(net7168),
    .Y(_04324_));
 sg13g2_xnor2_1 _17905_ (.Y(_04325_),
    .A(net7232),
    .B(net7167));
 sg13g2_nand3_1 _17906_ (.B(_04238_),
    .C(_04325_),
    .A(_04131_),
    .Y(_04326_));
 sg13g2_a21oi_1 _17907_ (.A1(_04269_),
    .A2(_04323_),
    .Y(_04327_),
    .B1(_04326_));
 sg13g2_nand3_1 _17908_ (.B(_04323_),
    .C(_04326_),
    .A(_04269_),
    .Y(_04328_));
 sg13g2_nor2b_1 _17909_ (.A(_04327_),
    .B_N(_04328_),
    .Y(_04329_));
 sg13g2_xnor2_1 _17910_ (.Y(_04330_),
    .A(_04322_),
    .B(_04329_));
 sg13g2_xnor2_1 _17911_ (.Y(_04331_),
    .A(_04306_),
    .B(_04330_));
 sg13g2_nand2b_1 _17912_ (.Y(_04332_),
    .B(_04255_),
    .A_N(_04271_));
 sg13g2_nand2_1 _17913_ (.Y(_04333_),
    .A(_04222_),
    .B(_04225_));
 sg13g2_o21ai_1 _17914_ (.B1(_04221_),
    .Y(_04334_),
    .A1(_04222_),
    .A2(_04225_));
 sg13g2_nand2_1 _17915_ (.Y(_04335_),
    .A(_04333_),
    .B(_04334_));
 sg13g2_a22oi_1 _17916_ (.Y(_04336_),
    .B1(net7633),
    .B2(_02282_),
    .A2(net7636),
    .A1(_03366_));
 sg13g2_nor2_1 _17917_ (.A(net7244),
    .B(net7161),
    .Y(_04337_));
 sg13g2_a22oi_1 _17918_ (.Y(_04338_),
    .B1(net7324),
    .B2(_01644_),
    .A2(net7326),
    .A1(_01662_));
 sg13g2_nor3_1 _17919_ (.A(net7236),
    .B(net7173),
    .C(_04338_),
    .Y(_04339_));
 sg13g2_o21ai_1 _17920_ (.B1(_04338_),
    .Y(_04340_),
    .A1(net7236),
    .A2(net7173));
 sg13g2_nor2b_1 _17921_ (.A(_04339_),
    .B_N(_04340_),
    .Y(_04341_));
 sg13g2_xnor2_1 _17922_ (.Y(_04342_),
    .A(_04337_),
    .B(_04341_));
 sg13g2_and2_1 _17923_ (.A(_04216_),
    .B(_04219_),
    .X(_04343_));
 sg13g2_nor2_1 _17924_ (.A(_04218_),
    .B(_04343_),
    .Y(_04344_));
 sg13g2_a21oi_1 _17925_ (.A1(_04256_),
    .A2(_04258_),
    .Y(_04345_),
    .B1(_04257_));
 sg13g2_nor2_1 _17926_ (.A(_04256_),
    .B(_04258_),
    .Y(_04346_));
 sg13g2_nor2_1 _17927_ (.A(_04345_),
    .B(_04346_),
    .Y(_04347_));
 sg13g2_xor2_1 _17928_ (.B(_04347_),
    .A(_04344_),
    .X(_04348_));
 sg13g2_xnor2_1 _17929_ (.Y(_04349_),
    .A(_04342_),
    .B(_04348_));
 sg13g2_nand2b_1 _17930_ (.Y(_04350_),
    .B(_04335_),
    .A_N(_04349_));
 sg13g2_xor2_1 _17931_ (.B(_04349_),
    .A(_04335_),
    .X(_04351_));
 sg13g2_xnor2_1 _17932_ (.Y(_04352_),
    .A(_04332_),
    .B(_04351_));
 sg13g2_xnor2_1 _17933_ (.Y(_04353_),
    .A(_04231_),
    .B(_04352_));
 sg13g2_nor2_1 _17934_ (.A(_04274_),
    .B(_04331_),
    .Y(_04354_));
 sg13g2_xnor2_1 _17935_ (.Y(_04355_),
    .A(_04274_),
    .B(_04331_));
 sg13g2_xnor2_1 _17936_ (.Y(_04356_),
    .A(_04353_),
    .B(_04355_));
 sg13g2_a21oi_1 _17937_ (.A1(_04235_),
    .A2(_04236_),
    .Y(_04357_),
    .B1(_04275_));
 sg13g2_nand3_1 _17938_ (.B(_04236_),
    .C(_04275_),
    .A(_04235_),
    .Y(_04358_));
 sg13g2_a21oi_1 _17939_ (.A1(_04200_),
    .A2(_04358_),
    .Y(_04359_),
    .B1(_04357_));
 sg13g2_a21oi_1 _17940_ (.A1(_04162_),
    .A2(_04233_),
    .Y(_04360_),
    .B1(_04234_));
 sg13g2_nand2_1 _17941_ (.Y(_04361_),
    .A(_04359_),
    .B(_04360_));
 sg13g2_nor2_1 _17942_ (.A(_04359_),
    .B(_04360_),
    .Y(_04362_));
 sg13g2_xor2_1 _17943_ (.B(_04360_),
    .A(_04359_),
    .X(_04363_));
 sg13g2_xnor2_1 _17944_ (.Y(_04364_),
    .A(_04356_),
    .B(_04363_));
 sg13g2_nor2b_1 _17945_ (.A(_04322_),
    .B_N(_04328_),
    .Y(_04365_));
 sg13g2_nor2_1 _17946_ (.A(_04327_),
    .B(_04365_),
    .Y(_04366_));
 sg13g2_a22oi_1 _17947_ (.Y(_04367_),
    .B1(net7633),
    .B2(_02362_),
    .A2(net7636),
    .A1(_03436_));
 sg13g2_nor2_1 _17948_ (.A(net7244),
    .B(net7156),
    .Y(_04368_));
 sg13g2_a22oi_1 _17949_ (.Y(_04369_),
    .B1(net7319),
    .B2(_01645_),
    .A2(net7326),
    .A1(_01663_));
 sg13g2_nor3_1 _17950_ (.A(net7236),
    .B(net7161),
    .C(_04369_),
    .Y(_04370_));
 sg13g2_o21ai_1 _17951_ (.B1(_04369_),
    .Y(_04371_),
    .A1(net7236),
    .A2(net7161));
 sg13g2_nand2b_1 _17952_ (.Y(_04372_),
    .B(_04371_),
    .A_N(_04370_));
 sg13g2_xnor2_1 _17953_ (.Y(_04373_),
    .A(_04368_),
    .B(_04372_));
 sg13g2_a21oi_1 _17954_ (.A1(_04337_),
    .A2(_04340_),
    .Y(_04374_),
    .B1(_04339_));
 sg13g2_a21oi_1 _17955_ (.A1(_04307_),
    .A2(_04308_),
    .Y(_04375_),
    .B1(_04309_));
 sg13g2_nor2_1 _17956_ (.A(_04307_),
    .B(_04308_),
    .Y(_04376_));
 sg13g2_nor2_1 _17957_ (.A(_04375_),
    .B(_04376_),
    .Y(_04377_));
 sg13g2_xnor2_1 _17958_ (.Y(_04378_),
    .A(_04374_),
    .B(_04377_));
 sg13g2_xnor2_1 _17959_ (.Y(_04379_),
    .A(_04373_),
    .B(_04378_));
 sg13g2_nor3_1 _17960_ (.A(_04218_),
    .B(_04343_),
    .C(_04347_),
    .Y(_04380_));
 sg13g2_nand2b_1 _17961_ (.Y(_04381_),
    .B(_04347_),
    .A_N(_04344_));
 sg13g2_a21o_1 _17962_ (.A2(_04381_),
    .A1(_04342_),
    .B1(_04380_),
    .X(_04382_));
 sg13g2_or2_1 _17963_ (.X(_04383_),
    .B(_04382_),
    .A(_04379_));
 sg13g2_xnor2_1 _17964_ (.Y(_04384_),
    .A(_04379_),
    .B(_04382_));
 sg13g2_nand2_1 _17965_ (.Y(_04385_),
    .A(_04350_),
    .B(_04384_));
 sg13g2_xnor2_1 _17966_ (.Y(_04386_),
    .A(_04350_),
    .B(_04384_));
 sg13g2_xnor2_1 _17967_ (.Y(_04387_),
    .A(_04366_),
    .B(_04386_));
 sg13g2_nand2_1 _17968_ (.Y(_04388_),
    .A(_04306_),
    .B(_04330_));
 sg13g2_nor2_1 _17969_ (.A(net7204),
    .B(net7194),
    .Y(_04389_));
 sg13g2_nor2_1 _17970_ (.A(net7201),
    .B(net7199),
    .Y(_04390_));
 sg13g2_nor2_1 _17971_ (.A(_03931_),
    .B(net7195),
    .Y(_04391_));
 sg13g2_xnor2_1 _17972_ (.Y(_04392_),
    .A(_04390_),
    .B(_04391_));
 sg13g2_xnor2_1 _17973_ (.Y(_04393_),
    .A(_04389_),
    .B(_04392_));
 sg13g2_nor2_1 _17974_ (.A(_04316_),
    .B(_04317_),
    .Y(_04394_));
 sg13g2_a21oi_1 _17975_ (.A1(_04316_),
    .A2(_04317_),
    .Y(_04395_),
    .B1(_04315_));
 sg13g2_nor2_1 _17976_ (.A(_04394_),
    .B(_04395_),
    .Y(_04396_));
 sg13g2_nor2_1 _17977_ (.A(net7225),
    .B(net7174),
    .Y(_04397_));
 sg13g2_nor2_1 _17978_ (.A(net7218),
    .B(_04142_),
    .Y(_04398_));
 sg13g2_nor2_1 _17979_ (.A(net7214),
    .B(net7190),
    .Y(_04399_));
 sg13g2_xor2_1 _17980_ (.B(_04399_),
    .A(_04398_),
    .X(_04400_));
 sg13g2_xnor2_1 _17981_ (.Y(_04401_),
    .A(_04397_),
    .B(_04400_));
 sg13g2_nor2b_1 _17982_ (.A(_04401_),
    .B_N(_04396_),
    .Y(_04402_));
 sg13g2_nand2b_1 _17983_ (.Y(_04403_),
    .B(_04401_),
    .A_N(_04396_));
 sg13g2_xor2_1 _17984_ (.B(_04401_),
    .A(_04396_),
    .X(_04404_));
 sg13g2_xnor2_1 _17985_ (.Y(_04405_),
    .A(_04393_),
    .B(_04404_));
 sg13g2_a21oi_1 _17986_ (.A1(_04314_),
    .A2(_04319_),
    .Y(_04406_),
    .B1(_04311_));
 sg13g2_nor2_1 _17987_ (.A(_04320_),
    .B(_04406_),
    .Y(_04407_));
 sg13g2_nand2_1 _17988_ (.Y(_04408_),
    .A(net7071),
    .B(_04299_));
 sg13g2_a21oi_1 _17989_ (.A1(_04250_),
    .A2(_04408_),
    .Y(_04409_),
    .B1(_04293_));
 sg13g2_xnor2_1 _17990_ (.Y(_04410_),
    .A(_04407_),
    .B(_04409_));
 sg13g2_xnor2_1 _17991_ (.Y(_04411_),
    .A(_04405_),
    .B(_04410_));
 sg13g2_xnor2_1 _17992_ (.Y(_04412_),
    .A(net6947),
    .B(_04302_));
 sg13g2_nand2b_1 _17993_ (.Y(_04413_),
    .B(_04412_),
    .A_N(_04304_));
 sg13g2_a22oi_1 _17994_ (.Y(_04414_),
    .B1(net7440),
    .B2(_02324_),
    .A2(net7638),
    .A1(_03403_));
 sg13g2_nor2_1 _17995_ (.A(net7250),
    .B(net7153),
    .Y(_04415_));
 sg13g2_nor2_1 _17996_ (.A(_03835_),
    .B(net7162),
    .Y(_04416_));
 sg13g2_xnor2_1 _17997_ (.Y(_04417_),
    .A(_04415_),
    .B(_04416_));
 sg13g2_nand2_1 _17998_ (.Y(_04418_),
    .A(_04290_),
    .B(_04291_));
 sg13g2_o21ai_1 _17999_ (.B1(_04289_),
    .Y(_04419_),
    .A1(_04290_),
    .A2(_04291_));
 sg13g2_nand2_1 _18000_ (.Y(_04420_),
    .A(_04418_),
    .B(_04419_));
 sg13g2_nor2_1 _18001_ (.A(net7224),
    .B(_04178_),
    .Y(_04421_));
 sg13g2_nor2_1 _18002_ (.A(_03908_),
    .B(net7184),
    .Y(_04422_));
 sg13g2_xnor2_1 _18003_ (.Y(_04423_),
    .A(_04421_),
    .B(_04422_));
 sg13g2_xnor2_1 _18004_ (.Y(_04424_),
    .A(_04324_),
    .B(_04423_));
 sg13g2_nand2_1 _18005_ (.Y(_04425_),
    .A(_04420_),
    .B(_04424_));
 sg13g2_xor2_1 _18006_ (.B(_04424_),
    .A(_04420_),
    .X(_04426_));
 sg13g2_nor2b_1 _18007_ (.A(_04417_),
    .B_N(_04426_),
    .Y(_04427_));
 sg13g2_xor2_1 _18008_ (.B(_04426_),
    .A(_04417_),
    .X(_04428_));
 sg13g2_nand2_1 _18009_ (.Y(_04429_),
    .A(_04413_),
    .B(_04428_));
 sg13g2_nor2_1 _18010_ (.A(_04413_),
    .B(_04428_),
    .Y(_04430_));
 sg13g2_xnor2_1 _18011_ (.Y(_04431_),
    .A(_04413_),
    .B(_04428_));
 sg13g2_xor2_1 _18012_ (.B(_04431_),
    .A(_04411_),
    .X(_04432_));
 sg13g2_nor2_1 _18013_ (.A(_04388_),
    .B(_04432_),
    .Y(_04433_));
 sg13g2_xnor2_1 _18014_ (.Y(_04434_),
    .A(_04388_),
    .B(_04432_));
 sg13g2_xnor2_1 _18015_ (.Y(_04435_),
    .A(_04387_),
    .B(_04434_));
 sg13g2_a21o_1 _18016_ (.A2(_04351_),
    .A1(_04231_),
    .B1(_04332_),
    .X(_04436_));
 sg13g2_o21ai_1 _18017_ (.B1(_04436_),
    .Y(_04437_),
    .A1(_04231_),
    .A2(_04351_));
 sg13g2_a21oi_1 _18018_ (.A1(_04274_),
    .A2(_04331_),
    .Y(_04438_),
    .B1(_04353_));
 sg13g2_o21ai_1 _18019_ (.B1(_04437_),
    .Y(_04439_),
    .A1(_04354_),
    .A2(_04438_));
 sg13g2_nor3_1 _18020_ (.A(_04354_),
    .B(_04437_),
    .C(_04438_),
    .Y(_04440_));
 sg13g2_or3_1 _18021_ (.A(_04354_),
    .B(_04437_),
    .C(_04438_),
    .X(_04441_));
 sg13g2_nand2_1 _18022_ (.Y(_04442_),
    .A(_04439_),
    .B(_04441_));
 sg13g2_xor2_1 _18023_ (.B(_04442_),
    .A(_04435_),
    .X(_04443_));
 sg13g2_a21o_1 _18024_ (.A2(_04409_),
    .A1(_04407_),
    .B1(_04405_),
    .X(_04444_));
 sg13g2_o21ai_1 _18025_ (.B1(_04444_),
    .Y(_04445_),
    .A1(_04407_),
    .A2(_04409_));
 sg13g2_a22oi_1 _18026_ (.Y(_04446_),
    .B1(net7633),
    .B2(_02438_),
    .A2(net7636),
    .A1(_03504_));
 sg13g2_nor2_1 _18027_ (.A(net7243),
    .B(net7149),
    .Y(_04447_));
 sg13g2_a22oi_1 _18028_ (.Y(_04448_),
    .B1(net7324),
    .B2(_01646_),
    .A2(net7326),
    .A1(_01664_));
 sg13g2_nor3_1 _18029_ (.A(net7238),
    .B(net7156),
    .C(_04448_),
    .Y(_04449_));
 sg13g2_o21ai_1 _18030_ (.B1(_04448_),
    .Y(_04450_),
    .A1(net7238),
    .A2(net7156));
 sg13g2_nand2b_1 _18031_ (.Y(_04451_),
    .B(_04450_),
    .A_N(_04449_));
 sg13g2_xnor2_1 _18032_ (.Y(_04452_),
    .A(_04447_),
    .B(_04451_));
 sg13g2_a21oi_1 _18033_ (.A1(_04368_),
    .A2(_04371_),
    .Y(_04453_),
    .B1(_04370_));
 sg13g2_a21oi_1 _18034_ (.A1(_04397_),
    .A2(_04398_),
    .Y(_04454_),
    .B1(_04399_));
 sg13g2_nor2_1 _18035_ (.A(_04397_),
    .B(_04398_),
    .Y(_04455_));
 sg13g2_nor2_1 _18036_ (.A(_04454_),
    .B(_04455_),
    .Y(_04456_));
 sg13g2_xnor2_1 _18037_ (.Y(_04457_),
    .A(_04453_),
    .B(_04456_));
 sg13g2_xnor2_1 _18038_ (.Y(_04458_),
    .A(_04452_),
    .B(_04457_));
 sg13g2_o21ai_1 _18039_ (.B1(_04374_),
    .Y(_04459_),
    .A1(_04375_),
    .A2(_04376_));
 sg13g2_nor3_1 _18040_ (.A(_04374_),
    .B(_04375_),
    .C(_04376_),
    .Y(_04460_));
 sg13g2_o21ai_1 _18041_ (.B1(_04459_),
    .Y(_04461_),
    .A1(_04373_),
    .A2(_04460_));
 sg13g2_nor2_1 _18042_ (.A(_04458_),
    .B(_04461_),
    .Y(_04462_));
 sg13g2_xnor2_1 _18043_ (.Y(_04463_),
    .A(_04458_),
    .B(_04461_));
 sg13g2_nand2_1 _18044_ (.Y(_04464_),
    .A(_04383_),
    .B(_04463_));
 sg13g2_xnor2_1 _18045_ (.Y(_04465_),
    .A(_04383_),
    .B(_04463_));
 sg13g2_xnor2_1 _18046_ (.Y(_04466_),
    .A(_04445_),
    .B(_04465_));
 sg13g2_a21oi_1 _18047_ (.A1(_04411_),
    .A2(_04429_),
    .Y(_04467_),
    .B1(_04430_));
 sg13g2_nor2_1 _18048_ (.A(net7204),
    .B(net7190),
    .Y(_04468_));
 sg13g2_nor2_1 _18049_ (.A(net7201),
    .B(net7192),
    .Y(_04469_));
 sg13g2_nor2_1 _18050_ (.A(net7199),
    .B(net7195),
    .Y(_04470_));
 sg13g2_xnor2_1 _18051_ (.Y(_04471_),
    .A(_04469_),
    .B(_04470_));
 sg13g2_xnor2_1 _18052_ (.Y(_04472_),
    .A(_04468_),
    .B(_04471_));
 sg13g2_nor2_1 _18053_ (.A(_04389_),
    .B(_04390_),
    .Y(_04473_));
 sg13g2_a21oi_1 _18054_ (.A1(_04389_),
    .A2(_04390_),
    .Y(_04474_),
    .B1(_04391_));
 sg13g2_nor2_1 _18055_ (.A(_04473_),
    .B(_04474_),
    .Y(_04475_));
 sg13g2_nor2_1 _18056_ (.A(net7225),
    .B(net7161),
    .Y(_04476_));
 sg13g2_nor2_1 _18057_ (.A(net7217),
    .B(_04215_),
    .Y(_04477_));
 sg13g2_nor2_1 _18058_ (.A(net7214),
    .B(net7183),
    .Y(_04478_));
 sg13g2_xor2_1 _18059_ (.B(_04478_),
    .A(_04476_),
    .X(_04479_));
 sg13g2_xnor2_1 _18060_ (.Y(_04480_),
    .A(_04477_),
    .B(_04479_));
 sg13g2_nor2b_1 _18061_ (.A(_04480_),
    .B_N(_04475_),
    .Y(_04481_));
 sg13g2_nand2b_1 _18062_ (.Y(_04482_),
    .B(_04480_),
    .A_N(_04475_));
 sg13g2_nor2b_1 _18063_ (.A(_04481_),
    .B_N(_04482_),
    .Y(_04483_));
 sg13g2_xor2_1 _18064_ (.B(_04483_),
    .A(_04472_),
    .X(_04484_));
 sg13g2_a21oi_1 _18065_ (.A1(_04393_),
    .A2(_04403_),
    .Y(_04485_),
    .B1(_04402_));
 sg13g2_nand2_1 _18066_ (.Y(_04486_),
    .A(_04425_),
    .B(_04485_));
 sg13g2_nor2_1 _18067_ (.A(_04425_),
    .B(_04485_),
    .Y(_04487_));
 sg13g2_xnor2_1 _18068_ (.Y(_04488_),
    .A(_04425_),
    .B(_04485_));
 sg13g2_xnor2_1 _18069_ (.Y(_04489_),
    .A(_04484_),
    .B(_04488_));
 sg13g2_or2_1 _18070_ (.X(_04490_),
    .B(net7168),
    .A(net7223));
 sg13g2_or2_1 _18071_ (.X(_04491_),
    .B(net7184),
    .A(_03931_));
 sg13g2_or2_1 _18072_ (.X(_04492_),
    .B(_04178_),
    .A(_03908_));
 sg13g2_xor2_1 _18073_ (.B(_04492_),
    .A(_04491_),
    .X(_04493_));
 sg13g2_xnor2_1 _18074_ (.Y(_04494_),
    .A(_04490_),
    .B(_04493_));
 sg13g2_a21oi_1 _18075_ (.A1(_04324_),
    .A2(_04421_),
    .Y(_04495_),
    .B1(_04422_));
 sg13g2_nor2_1 _18076_ (.A(_04324_),
    .B(_04421_),
    .Y(_04496_));
 sg13g2_a21oi_1 _18077_ (.A1(_03833_),
    .A2(_03834_),
    .Y(_04497_),
    .B1(_04414_));
 sg13g2_nand2b_1 _18078_ (.Y(_04498_),
    .B(_04497_),
    .A_N(_04304_));
 sg13g2_nor3_1 _18079_ (.A(_04495_),
    .B(_04496_),
    .C(_04498_),
    .Y(_04499_));
 sg13g2_o21ai_1 _18080_ (.B1(_04498_),
    .Y(_04500_),
    .A1(_04495_),
    .A2(_04496_));
 sg13g2_nand2b_1 _18081_ (.Y(_04501_),
    .B(_04500_),
    .A_N(_04499_));
 sg13g2_xnor2_1 _18082_ (.Y(_04502_),
    .A(_04494_),
    .B(_04501_));
 sg13g2_a22oi_1 _18083_ (.Y(_04503_),
    .B1(net7440),
    .B2(_02399_),
    .A2(net7638),
    .A1(net7330));
 sg13g2_nor2_1 _18084_ (.A(net7250),
    .B(net7144),
    .Y(_04504_));
 sg13g2_nor2_1 _18085_ (.A(net7233),
    .B(net7162),
    .Y(_04505_));
 sg13g2_xnor2_1 _18086_ (.Y(_04506_),
    .A(_04504_),
    .B(_04505_));
 sg13g2_xnor2_1 _18087_ (.Y(_04507_),
    .A(_04497_),
    .B(_04506_));
 sg13g2_nand2_1 _18088_ (.Y(_04508_),
    .A(_04502_),
    .B(_04507_));
 sg13g2_xor2_1 _18089_ (.B(_04507_),
    .A(_04502_),
    .X(_04509_));
 sg13g2_and2_1 _18090_ (.A(_04427_),
    .B(_04509_),
    .X(_04510_));
 sg13g2_or2_1 _18091_ (.X(_04511_),
    .B(_04509_),
    .A(_04427_));
 sg13g2_xor2_1 _18092_ (.B(_04509_),
    .A(_04427_),
    .X(_04512_));
 sg13g2_xnor2_1 _18093_ (.Y(_04513_),
    .A(_04489_),
    .B(_04512_));
 sg13g2_nor2_1 _18094_ (.A(_04467_),
    .B(_04513_),
    .Y(_04514_));
 sg13g2_xor2_1 _18095_ (.B(_04513_),
    .A(_04467_),
    .X(_04515_));
 sg13g2_xor2_1 _18096_ (.B(_04515_),
    .A(_04466_),
    .X(_04516_));
 sg13g2_o21ai_1 _18097_ (.B1(_04366_),
    .Y(_04517_),
    .A1(_04350_),
    .A2(_04384_));
 sg13g2_and2_1 _18098_ (.A(_04385_),
    .B(_04517_),
    .X(_04518_));
 sg13g2_a21oi_1 _18099_ (.A1(_04388_),
    .A2(_04432_),
    .Y(_04519_),
    .B1(_04387_));
 sg13g2_o21ai_1 _18100_ (.B1(_04518_),
    .Y(_04520_),
    .A1(_04433_),
    .A2(_04519_));
 sg13g2_nor3_1 _18101_ (.A(_04433_),
    .B(_04518_),
    .C(_04519_),
    .Y(_04521_));
 sg13g2_or3_1 _18102_ (.A(_04433_),
    .B(_04518_),
    .C(_04519_),
    .X(_04522_));
 sg13g2_and2_1 _18103_ (.A(_04520_),
    .B(_04522_),
    .X(_04523_));
 sg13g2_xnor2_1 _18104_ (.Y(_04524_),
    .A(_04516_),
    .B(_04523_));
 sg13g2_o21ai_1 _18105_ (.B1(_04511_),
    .Y(_04525_),
    .A1(_04489_),
    .A2(_04510_));
 sg13g2_nor2_1 _18106_ (.A(net7207),
    .B(net7181),
    .Y(_04526_));
 sg13g2_nor2_1 _18107_ (.A(net7203),
    .B(net7190),
    .Y(_04527_));
 sg13g2_nor2_1 _18108_ (.A(net7197),
    .B(net7192),
    .Y(_04528_));
 sg13g2_xnor2_1 _18109_ (.Y(_04529_),
    .A(_04527_),
    .B(_04528_));
 sg13g2_xnor2_1 _18110_ (.Y(_04530_),
    .A(_04526_),
    .B(_04529_));
 sg13g2_a21oi_1 _18111_ (.A1(_04468_),
    .A2(_04470_),
    .Y(_04531_),
    .B1(_04469_));
 sg13g2_nor2_1 _18112_ (.A(_04468_),
    .B(_04470_),
    .Y(_04532_));
 sg13g2_nor2_1 _18113_ (.A(_04531_),
    .B(_04532_),
    .Y(_04533_));
 sg13g2_nor2_1 _18114_ (.A(net7228),
    .B(net7156),
    .Y(_04534_));
 sg13g2_nor2_1 _18115_ (.A(net7217),
    .B(net7159),
    .Y(_04535_));
 sg13g2_nor2_1 _18116_ (.A(net7215),
    .B(_04215_),
    .Y(_04536_));
 sg13g2_xnor2_1 _18117_ (.Y(_04537_),
    .A(_04535_),
    .B(_04536_));
 sg13g2_xnor2_1 _18118_ (.Y(_04538_),
    .A(_04534_),
    .B(_04537_));
 sg13g2_nand2_1 _18119_ (.Y(_04539_),
    .A(_04533_),
    .B(_04538_));
 sg13g2_xnor2_1 _18120_ (.Y(_04540_),
    .A(_04533_),
    .B(_04538_));
 sg13g2_xnor2_1 _18121_ (.Y(_04541_),
    .A(_04530_),
    .B(_04540_));
 sg13g2_a21oi_1 _18122_ (.A1(_04472_),
    .A2(_04482_),
    .Y(_04542_),
    .B1(_04481_));
 sg13g2_a21oi_1 _18123_ (.A1(_04494_),
    .A2(_04500_),
    .Y(_04543_),
    .B1(_04499_));
 sg13g2_xnor2_1 _18124_ (.Y(_04544_),
    .A(_04542_),
    .B(_04543_));
 sg13g2_xnor2_1 _18125_ (.Y(_04545_),
    .A(_04541_),
    .B(_04544_));
 sg13g2_or2_1 _18126_ (.X(_04546_),
    .B(_04492_),
    .A(_04491_));
 sg13g2_a21o_1 _18127_ (.A2(_04492_),
    .A1(_04491_),
    .B1(_04490_),
    .X(_04547_));
 sg13g2_nand2_1 _18128_ (.Y(_04548_),
    .A(_04546_),
    .B(_04547_));
 sg13g2_nand2_1 _18129_ (.Y(_04549_),
    .A(_04497_),
    .B(_04505_));
 sg13g2_o21ai_1 _18130_ (.B1(_04504_),
    .Y(_04550_),
    .A1(_04497_),
    .A2(_04505_));
 sg13g2_nand2_1 _18131_ (.Y(_04551_),
    .A(_04549_),
    .B(_04550_));
 sg13g2_nor2_1 _18132_ (.A(_03908_),
    .B(net7168),
    .Y(_04552_));
 sg13g2_or2_1 _18133_ (.X(_04553_),
    .B(net7184),
    .A(_03981_));
 sg13g2_or2_1 _18134_ (.X(_04554_),
    .B(_04178_),
    .A(_03931_));
 sg13g2_xnor2_1 _18135_ (.Y(_04555_),
    .A(_04553_),
    .B(_04554_));
 sg13g2_xnor2_1 _18136_ (.Y(_04556_),
    .A(_04552_),
    .B(_04555_));
 sg13g2_xnor2_1 _18137_ (.Y(_04557_),
    .A(_04548_),
    .B(net6946));
 sg13g2_xnor2_1 _18138_ (.Y(_04558_),
    .A(_04551_),
    .B(_04557_));
 sg13g2_and3_1 _18139_ (.X(_04559_),
    .A(_03520_),
    .B(_03525_),
    .C(_03815_));
 sg13g2_a22oi_1 _18140_ (.Y(_04560_),
    .B1(_04559_),
    .B2(_03536_),
    .A2(net7440),
    .A1(_02475_));
 sg13g2_nor2_1 _18141_ (.A(net7249),
    .B(net7143),
    .Y(_04561_));
 sg13g2_or2_1 _18142_ (.X(_04562_),
    .B(net7153),
    .A(net7233));
 sg13g2_nor2_1 _18143_ (.A(_03835_),
    .B(net7144),
    .Y(_04563_));
 sg13g2_or2_1 _18144_ (.X(_04564_),
    .B(net7162),
    .A(net7223));
 sg13g2_xnor2_1 _18145_ (.Y(_04565_),
    .A(_04562_),
    .B(_04564_));
 sg13g2_xnor2_1 _18146_ (.Y(_04566_),
    .A(_04563_),
    .B(_04565_));
 sg13g2_xor2_1 _18147_ (.B(_04566_),
    .A(_04561_),
    .X(_04567_));
 sg13g2_nand2_1 _18148_ (.Y(_04568_),
    .A(_04558_),
    .B(_04567_));
 sg13g2_xnor2_1 _18149_ (.Y(_04569_),
    .A(_04558_),
    .B(_04567_));
 sg13g2_xor2_1 _18150_ (.B(_04569_),
    .A(_04508_),
    .X(_04570_));
 sg13g2_xnor2_1 _18151_ (.Y(_04571_),
    .A(_04545_),
    .B(_04570_));
 sg13g2_a21oi_1 _18152_ (.A1(_04484_),
    .A2(_04486_),
    .Y(_04572_),
    .B1(_04487_));
 sg13g2_o21ai_1 _18153_ (.B1(_04453_),
    .Y(_04573_),
    .A1(_04454_),
    .A2(_04455_));
 sg13g2_nor3_1 _18154_ (.A(_04453_),
    .B(_04454_),
    .C(_04455_),
    .Y(_04574_));
 sg13g2_o21ai_1 _18155_ (.B1(_04573_),
    .Y(_04575_),
    .A1(_04452_),
    .A2(_04574_));
 sg13g2_a22oi_1 _18156_ (.Y(_04576_),
    .B1(net7633),
    .B2(_02502_),
    .A2(net7636),
    .A1(_03575_));
 sg13g2_nor2_1 _18157_ (.A(net7243),
    .B(_04576_),
    .Y(_04577_));
 sg13g2_a22oi_1 _18158_ (.Y(_04578_),
    .B1(net7324),
    .B2(_01647_),
    .A2(net7326),
    .A1(_01665_));
 sg13g2_nor3_1 _18159_ (.A(net7238),
    .B(net7149),
    .C(_04578_),
    .Y(_04579_));
 sg13g2_o21ai_1 _18160_ (.B1(_04578_),
    .Y(_04580_),
    .A1(net7238),
    .A2(net7149));
 sg13g2_nor2b_1 _18161_ (.A(_04579_),
    .B_N(_04580_),
    .Y(_04581_));
 sg13g2_xnor2_1 _18162_ (.Y(_04582_),
    .A(_04577_),
    .B(_04581_));
 sg13g2_and2_1 _18163_ (.A(_04447_),
    .B(_04450_),
    .X(_04583_));
 sg13g2_nor2_1 _18164_ (.A(_04449_),
    .B(_04583_),
    .Y(_04584_));
 sg13g2_nor2_1 _18165_ (.A(_04477_),
    .B(_04478_),
    .Y(_04585_));
 sg13g2_a21oi_1 _18166_ (.A1(_04477_),
    .A2(_04478_),
    .Y(_04586_),
    .B1(_04476_));
 sg13g2_nor2_1 _18167_ (.A(_04585_),
    .B(_04586_),
    .Y(_04587_));
 sg13g2_xor2_1 _18168_ (.B(_04587_),
    .A(_04584_),
    .X(_04588_));
 sg13g2_xnor2_1 _18169_ (.Y(_04589_),
    .A(_04582_),
    .B(_04588_));
 sg13g2_nor2_1 _18170_ (.A(_04575_),
    .B(_04589_),
    .Y(_04590_));
 sg13g2_xnor2_1 _18171_ (.Y(_04591_),
    .A(_04575_),
    .B(_04589_));
 sg13g2_nand2b_1 _18172_ (.Y(_04592_),
    .B(_04462_),
    .A_N(_04591_));
 sg13g2_nor2b_1 _18173_ (.A(_04462_),
    .B_N(_04591_),
    .Y(_04593_));
 sg13g2_xnor2_1 _18174_ (.Y(_04594_),
    .A(_04462_),
    .B(_04591_));
 sg13g2_xor2_1 _18175_ (.B(_04594_),
    .A(_04572_),
    .X(_04595_));
 sg13g2_xnor2_1 _18176_ (.Y(_04596_),
    .A(_04525_),
    .B(_04595_));
 sg13g2_xnor2_1 _18177_ (.Y(_04597_),
    .A(_04571_),
    .B(_04596_));
 sg13g2_a21oi_1 _18178_ (.A1(_04467_),
    .A2(_04513_),
    .Y(_04598_),
    .B1(_04466_));
 sg13g2_o21ai_1 _18179_ (.B1(_04445_),
    .Y(_04599_),
    .A1(_04383_),
    .A2(_04463_));
 sg13g2_and2_1 _18180_ (.A(_04464_),
    .B(_04599_),
    .X(_04600_));
 sg13g2_nor3_1 _18181_ (.A(_04514_),
    .B(_04598_),
    .C(_04600_),
    .Y(_04601_));
 sg13g2_o21ai_1 _18182_ (.B1(_04600_),
    .Y(_04602_),
    .A1(_04514_),
    .A2(_04598_));
 sg13g2_nor2b_1 _18183_ (.A(_04601_),
    .B_N(_04602_),
    .Y(_04603_));
 sg13g2_xnor2_1 _18184_ (.Y(_04604_),
    .A(_04597_),
    .B(_04603_));
 sg13g2_nand2_1 _18185_ (.Y(_04605_),
    .A(_04508_),
    .B(_04569_));
 sg13g2_nor2_1 _18186_ (.A(_04508_),
    .B(_04569_),
    .Y(_04606_));
 sg13g2_a21oi_1 _18187_ (.A1(_04545_),
    .A2(_04605_),
    .Y(_04607_),
    .B1(_04606_));
 sg13g2_nor2_1 _18188_ (.A(net7207),
    .B(net7175),
    .Y(_04608_));
 sg13g2_nor2_1 _18189_ (.A(net7203),
    .B(net7181),
    .Y(_04609_));
 sg13g2_nor2_1 _18190_ (.A(net7197),
    .B(net7190),
    .Y(_04610_));
 sg13g2_xor2_1 _18191_ (.B(_04610_),
    .A(_04609_),
    .X(_04611_));
 sg13g2_xnor2_1 _18192_ (.Y(_04612_),
    .A(_04608_),
    .B(_04611_));
 sg13g2_a21o_1 _18193_ (.A2(_04528_),
    .A1(_04526_),
    .B1(_04527_),
    .X(_04613_));
 sg13g2_o21ai_1 _18194_ (.B1(_04613_),
    .Y(_04614_),
    .A1(_04526_),
    .A2(_04528_));
 sg13g2_nor2_1 _18195_ (.A(net7228),
    .B(net7149),
    .Y(_04615_));
 sg13g2_nor2_1 _18196_ (.A(net7219),
    .B(net7156),
    .Y(_04616_));
 sg13g2_nor2_1 _18197_ (.A(net7215),
    .B(net7159),
    .Y(_04617_));
 sg13g2_xor2_1 _18198_ (.B(_04617_),
    .A(_04615_),
    .X(_04618_));
 sg13g2_xnor2_1 _18199_ (.Y(_04619_),
    .A(_04616_),
    .B(_04618_));
 sg13g2_nand2_1 _18200_ (.Y(_04620_),
    .A(_04614_),
    .B(_04619_));
 sg13g2_xor2_1 _18201_ (.B(_04619_),
    .A(_04614_),
    .X(_04621_));
 sg13g2_xor2_1 _18202_ (.B(_04621_),
    .A(_04612_),
    .X(_04622_));
 sg13g2_xnor2_1 _18203_ (.Y(_04623_),
    .A(_04612_),
    .B(_04621_));
 sg13g2_o21ai_1 _18204_ (.B1(_04530_),
    .Y(_04624_),
    .A1(_04533_),
    .A2(_04538_));
 sg13g2_a22oi_1 _18205_ (.Y(_04625_),
    .B1(_04549_),
    .B2(_04550_),
    .A2(_04547_),
    .A1(_04546_));
 sg13g2_nand4_1 _18206_ (.B(_04547_),
    .C(_04549_),
    .A(_04546_),
    .Y(_04626_),
    .D(_04550_));
 sg13g2_o21ai_1 _18207_ (.B1(_04626_),
    .Y(_04627_),
    .A1(_04556_),
    .A2(_04625_));
 sg13g2_nand3_1 _18208_ (.B(_04624_),
    .C(_04627_),
    .A(_04539_),
    .Y(_04628_));
 sg13g2_a21oi_1 _18209_ (.A1(_04539_),
    .A2(_04624_),
    .Y(_04629_),
    .B1(net6898));
 sg13g2_a21o_1 _18210_ (.A2(_04624_),
    .A1(_04539_),
    .B1(net6898),
    .X(_04630_));
 sg13g2_and3_1 _18211_ (.X(_04631_),
    .A(_04622_),
    .B(_04628_),
    .C(_04630_));
 sg13g2_a21oi_1 _18212_ (.A1(_04628_),
    .A2(_04630_),
    .Y(_04632_),
    .B1(_04622_));
 sg13g2_nor2_1 _18213_ (.A(_04631_),
    .B(_04632_),
    .Y(_04633_));
 sg13g2_nor2_1 _18214_ (.A(net7210),
    .B(net7168),
    .Y(_04634_));
 sg13g2_nor2_1 _18215_ (.A(_03981_),
    .B(net7177),
    .Y(_04635_));
 sg13g2_nor2_1 _18216_ (.A(net7193),
    .B(net7184),
    .Y(_04636_));
 sg13g2_xor2_1 _18217_ (.B(_04636_),
    .A(_04635_),
    .X(_04637_));
 sg13g2_xnor2_1 _18218_ (.Y(_04638_),
    .A(_04634_),
    .B(_04637_));
 sg13g2_nor2_1 _18219_ (.A(_04562_),
    .B(_04564_),
    .Y(_04639_));
 sg13g2_nand2_1 _18220_ (.Y(_04640_),
    .A(_04562_),
    .B(_04564_));
 sg13g2_a21oi_1 _18221_ (.A1(_04563_),
    .A2(_04640_),
    .Y(_04641_),
    .B1(_04639_));
 sg13g2_nor2_1 _18222_ (.A(_04553_),
    .B(_04554_),
    .Y(_04642_));
 sg13g2_nand2_1 _18223_ (.Y(_04643_),
    .A(_04553_),
    .B(_04554_));
 sg13g2_a21oi_1 _18224_ (.A1(_04552_),
    .A2(_04643_),
    .Y(_04644_),
    .B1(_04642_));
 sg13g2_xor2_1 _18225_ (.B(_04644_),
    .A(_04641_),
    .X(_04645_));
 sg13g2_xnor2_1 _18226_ (.Y(_04646_),
    .A(_04638_),
    .B(_04645_));
 sg13g2_and4_1 _18227_ (.A(_02519_),
    .B(_02521_),
    .C(_02523_),
    .D(net7440),
    .X(_04647_));
 sg13g2_and3_1 _18228_ (.X(_04648_),
    .A(_03601_),
    .B(_03606_),
    .C(_03815_));
 sg13g2_a22oi_1 _18229_ (.Y(_04649_),
    .B1(_04648_),
    .B2(_03592_),
    .A2(_04647_),
    .A1(_02533_));
 sg13g2_inv_1 _18230_ (.Y(_04650_),
    .A(net7134));
 sg13g2_nor2_1 _18231_ (.A(net7250),
    .B(net7135),
    .Y(_04651_));
 sg13g2_nor2_1 _18232_ (.A(_03835_),
    .B(net7140),
    .Y(_04652_));
 sg13g2_xnor2_1 _18233_ (.Y(_04653_),
    .A(_04651_),
    .B(_04652_));
 sg13g2_or2_1 _18234_ (.X(_04654_),
    .B(net7144),
    .A(net7233));
 sg13g2_or2_1 _18235_ (.X(_04655_),
    .B(net7162),
    .A(net7212));
 sg13g2_or2_1 _18236_ (.X(_04656_),
    .B(net7153),
    .A(net7223));
 sg13g2_xnor2_1 _18237_ (.Y(_04657_),
    .A(_04654_),
    .B(_04656_));
 sg13g2_xor2_1 _18238_ (.B(_04657_),
    .A(_04655_),
    .X(_04658_));
 sg13g2_nor2b_1 _18239_ (.A(_04653_),
    .B_N(_04658_),
    .Y(_04659_));
 sg13g2_xor2_1 _18240_ (.B(_04658_),
    .A(_04653_),
    .X(_04660_));
 sg13g2_nand2_1 _18241_ (.Y(_04661_),
    .A(_04561_),
    .B(_04566_));
 sg13g2_xnor2_1 _18242_ (.Y(_04662_),
    .A(_04660_),
    .B(_04661_));
 sg13g2_xnor2_1 _18243_ (.Y(_04663_),
    .A(_04646_),
    .B(_04662_));
 sg13g2_xor2_1 _18244_ (.B(_04663_),
    .A(_04568_),
    .X(_04664_));
 sg13g2_xnor2_1 _18245_ (.Y(_04665_),
    .A(_04633_),
    .B(_04664_));
 sg13g2_nand2_1 _18246_ (.Y(_04666_),
    .A(_04542_),
    .B(_04543_));
 sg13g2_nor2_1 _18247_ (.A(_04542_),
    .B(_04543_),
    .Y(_04667_));
 sg13g2_o21ai_1 _18248_ (.B1(_04666_),
    .Y(_04668_),
    .A1(_04541_),
    .A2(_04667_));
 sg13g2_nor3_1 _18249_ (.A(_04449_),
    .B(_04583_),
    .C(_04587_),
    .Y(_04669_));
 sg13g2_nand2b_1 _18250_ (.Y(_04670_),
    .B(_04587_),
    .A_N(_04584_));
 sg13g2_a21oi_1 _18251_ (.A1(_04582_),
    .A2(_04670_),
    .Y(_04671_),
    .B1(_04669_));
 sg13g2_mux2_1 _18252_ (.A0(_03625_),
    .A1(_03627_),
    .S(net7807),
    .X(_04672_));
 sg13g2_mux4_1 _18253_ (.S0(net7483),
    .A0(_03614_),
    .A1(_03615_),
    .A2(_03618_),
    .A3(_03617_),
    .S1(net7807),
    .X(_04673_));
 sg13g2_a221oi_1 _18254_ (.B2(_03822_),
    .C1(net7805),
    .B1(_04672_),
    .A1(_02548_),
    .Y(_04674_),
    .A2(net7634));
 sg13g2_a22oi_1 _18255_ (.Y(_04675_),
    .B1(_04673_),
    .B2(_03822_),
    .A2(net7634),
    .A1(_02540_));
 sg13g2_nand2_1 _18256_ (.Y(_04676_),
    .A(net7805),
    .B(_04675_));
 sg13g2_nor2b_1 _18257_ (.A(_04674_),
    .B_N(_04676_),
    .Y(_04677_));
 sg13g2_nand2b_1 _18258_ (.Y(_04678_),
    .B(_04676_),
    .A_N(_04674_));
 sg13g2_nor2_1 _18259_ (.A(net7243),
    .B(_04678_),
    .Y(_04679_));
 sg13g2_and2_1 _18260_ (.A(_01666_),
    .B(net7326),
    .X(_04680_));
 sg13g2_a21o_1 _18261_ (.A2(net7324),
    .A1(_01648_),
    .B1(_04680_),
    .X(_04681_));
 sg13g2_nor2_1 _18262_ (.A(net7237),
    .B(_04576_),
    .Y(_04682_));
 sg13g2_xnor2_1 _18263_ (.Y(_04683_),
    .A(_04681_),
    .B(_04682_));
 sg13g2_xnor2_1 _18264_ (.Y(_04684_),
    .A(_04679_),
    .B(_04683_));
 sg13g2_a21oi_1 _18265_ (.A1(_04577_),
    .A2(_04580_),
    .Y(_04685_),
    .B1(_04579_));
 sg13g2_a21oi_1 _18266_ (.A1(_04534_),
    .A2(_04536_),
    .Y(_04686_),
    .B1(_04535_));
 sg13g2_nor2_1 _18267_ (.A(_04534_),
    .B(_04536_),
    .Y(_04687_));
 sg13g2_nor2_1 _18268_ (.A(_04686_),
    .B(_04687_),
    .Y(_04688_));
 sg13g2_xnor2_1 _18269_ (.Y(_04689_),
    .A(_04685_),
    .B(_04688_));
 sg13g2_xnor2_1 _18270_ (.Y(_04690_),
    .A(_04684_),
    .B(_04689_));
 sg13g2_nand2b_1 _18271_ (.Y(_04691_),
    .B(_04671_),
    .A_N(_04690_));
 sg13g2_xnor2_1 _18272_ (.Y(_04692_),
    .A(_04671_),
    .B(_04690_));
 sg13g2_nand2_1 _18273_ (.Y(_04693_),
    .A(_04590_),
    .B(_04692_));
 sg13g2_nor2_1 _18274_ (.A(_04590_),
    .B(_04692_),
    .Y(_04694_));
 sg13g2_xnor2_1 _18275_ (.Y(_04695_),
    .A(_04590_),
    .B(_04692_));
 sg13g2_xnor2_1 _18276_ (.Y(_04696_),
    .A(_04668_),
    .B(_04695_));
 sg13g2_nand2_1 _18277_ (.Y(_04697_),
    .A(_04665_),
    .B(_04696_));
 sg13g2_xnor2_1 _18278_ (.Y(_04698_),
    .A(_04607_),
    .B(_04696_));
 sg13g2_xnor2_1 _18279_ (.Y(_04699_),
    .A(_04665_),
    .B(_04698_));
 sg13g2_a21oi_1 _18280_ (.A1(_04572_),
    .A2(_04592_),
    .Y(_04700_),
    .B1(_04593_));
 sg13g2_nand2_1 _18281_ (.Y(_04701_),
    .A(_04571_),
    .B(_04595_));
 sg13g2_o21ai_1 _18282_ (.B1(_04525_),
    .Y(_04702_),
    .A1(_04571_),
    .A2(_04595_));
 sg13g2_nand2_1 _18283_ (.Y(_04703_),
    .A(_04701_),
    .B(_04702_));
 sg13g2_xnor2_1 _18284_ (.Y(_04704_),
    .A(_04700_),
    .B(_04703_));
 sg13g2_xnor2_1 _18285_ (.Y(_04705_),
    .A(_04699_),
    .B(_04704_));
 sg13g2_nor2_1 _18286_ (.A(net7207),
    .B(net7159),
    .Y(_04706_));
 sg13g2_nor2_1 _18287_ (.A(net7197),
    .B(net7181),
    .Y(_04707_));
 sg13g2_nor2_1 _18288_ (.A(net7203),
    .B(net7175),
    .Y(_04708_));
 sg13g2_xnor2_1 _18289_ (.Y(_04709_),
    .A(_04707_),
    .B(_04708_));
 sg13g2_xnor2_1 _18290_ (.Y(_04710_),
    .A(_04706_),
    .B(_04709_));
 sg13g2_a21oi_1 _18291_ (.A1(_04608_),
    .A2(_04610_),
    .Y(_04711_),
    .B1(_04609_));
 sg13g2_nor2_1 _18292_ (.A(_04608_),
    .B(_04610_),
    .Y(_04712_));
 sg13g2_nor2_1 _18293_ (.A(_04711_),
    .B(_04712_),
    .Y(_04713_));
 sg13g2_nor2_1 _18294_ (.A(net7228),
    .B(_04576_),
    .Y(_04714_));
 sg13g2_nor2_1 _18295_ (.A(net7215),
    .B(net7156),
    .Y(_04715_));
 sg13g2_nor2_1 _18296_ (.A(net7219),
    .B(net7148),
    .Y(_04716_));
 sg13g2_xnor2_1 _18297_ (.Y(_04717_),
    .A(_04715_),
    .B(_04716_));
 sg13g2_xnor2_1 _18298_ (.Y(_04718_),
    .A(_04714_),
    .B(_04717_));
 sg13g2_nand2_1 _18299_ (.Y(_04719_),
    .A(_04713_),
    .B(_04718_));
 sg13g2_xor2_1 _18300_ (.B(_04718_),
    .A(_04713_),
    .X(_04720_));
 sg13g2_xnor2_1 _18301_ (.Y(_04721_),
    .A(_04710_),
    .B(_04720_));
 sg13g2_o21ai_1 _18302_ (.B1(_04612_),
    .Y(_04722_),
    .A1(_04614_),
    .A2(_04619_));
 sg13g2_nand2_1 _18303_ (.Y(_04723_),
    .A(_04641_),
    .B(_04644_));
 sg13g2_o21ai_1 _18304_ (.B1(_04638_),
    .Y(_04724_),
    .A1(_04641_),
    .A2(_04644_));
 sg13g2_a22oi_1 _18305_ (.Y(_04725_),
    .B1(_04723_),
    .B2(_04724_),
    .A2(_04722_),
    .A1(_04620_));
 sg13g2_nand4_1 _18306_ (.B(_04722_),
    .C(_04723_),
    .A(_04620_),
    .Y(_04726_),
    .D(_04724_));
 sg13g2_nor2b_1 _18307_ (.A(_04725_),
    .B_N(_04726_),
    .Y(_04727_));
 sg13g2_xor2_1 _18308_ (.B(_04727_),
    .A(_04721_),
    .X(_04728_));
 sg13g2_nor2_1 _18309_ (.A(net7222),
    .B(net7144),
    .Y(_04729_));
 sg13g2_nor2_1 _18310_ (.A(net7210),
    .B(net7163),
    .Y(_04730_));
 sg13g2_nor2_1 _18311_ (.A(net7212),
    .B(net7152),
    .Y(_04731_));
 sg13g2_xnor2_1 _18312_ (.Y(_04732_),
    .A(_04729_),
    .B(_04731_));
 sg13g2_xnor2_1 _18313_ (.Y(_04733_),
    .A(_04730_),
    .B(_04732_));
 sg13g2_a21oi_1 _18314_ (.A1(_03833_),
    .A2(_03834_),
    .Y(_04734_),
    .B1(_04649_));
 sg13g2_nand4_1 _18315_ (.B(_08239_),
    .C(_03601_),
    .A(_08032_),
    .Y(_04735_),
    .D(_03606_));
 sg13g2_nor2b_1 _18316_ (.A(_04735_),
    .B_N(_03592_),
    .Y(_04736_));
 sg13g2_and2_1 _18317_ (.A(net7637),
    .B(_04736_),
    .X(_04737_));
 sg13g2_nand3b_1 _18318_ (.B(net7637),
    .C(_03592_),
    .Y(_04738_),
    .A_N(_04735_));
 sg13g2_nor2_1 _18319_ (.A(_03846_),
    .B(net7143),
    .Y(_04739_));
 sg13g2_nor3_1 _18320_ (.A(net7065),
    .B(_04738_),
    .C(_04739_),
    .Y(_04740_));
 sg13g2_and3_1 _18321_ (.X(_04741_),
    .A(net7230),
    .B(_04734_),
    .C(_04738_));
 sg13g2_and4_1 _18322_ (.A(_08032_),
    .B(_08249_),
    .C(_03592_),
    .D(_03607_),
    .X(_04742_));
 sg13g2_and2_1 _18323_ (.A(net7637),
    .B(_04742_),
    .X(_04743_));
 sg13g2_inv_1 _18324_ (.Y(_04744_),
    .A(_04743_));
 sg13g2_xnor2_1 _18325_ (.Y(_04745_),
    .A(net7065),
    .B(_04743_));
 sg13g2_o21ai_1 _18326_ (.B1(net7249),
    .Y(_04746_),
    .A1(_04740_),
    .A2(_04741_));
 sg13g2_and2_1 _18327_ (.A(_04739_),
    .B(_04745_),
    .X(_04747_));
 sg13g2_and2_1 _18328_ (.A(net7143),
    .B(net7065),
    .X(_04748_));
 sg13g2_a22oi_1 _18329_ (.Y(_04749_),
    .B1(_04748_),
    .B2(_04744_),
    .A2(_04745_),
    .A1(_04739_));
 sg13g2_o21ai_1 _18330_ (.B1(net7071),
    .Y(_04750_),
    .A1(_04739_),
    .A2(_04748_));
 sg13g2_nand3_1 _18331_ (.B(_04749_),
    .C(_04750_),
    .A(_04746_),
    .Y(_04751_));
 sg13g2_xnor2_1 _18332_ (.Y(_04752_),
    .A(_04733_),
    .B(_04751_));
 sg13g2_nor2_1 _18333_ (.A(_03981_),
    .B(net7169),
    .Y(_04753_));
 sg13g2_nor2_1 _18334_ (.A(net7190),
    .B(net7186),
    .Y(_04754_));
 sg13g2_nor2_1 _18335_ (.A(net7193),
    .B(net7177),
    .Y(_04755_));
 sg13g2_xor2_1 _18336_ (.B(_04755_),
    .A(_04754_),
    .X(_04756_));
 sg13g2_xnor2_1 _18337_ (.Y(_04757_),
    .A(_04753_),
    .B(_04756_));
 sg13g2_or4_1 _18338_ (.A(net7222),
    .B(net7212),
    .C(net7162),
    .D(net7153),
    .X(_04758_));
 sg13g2_nand2_1 _18339_ (.Y(_04759_),
    .A(_04655_),
    .B(_04656_));
 sg13g2_a21o_1 _18340_ (.A2(_04656_),
    .A1(_04655_),
    .B1(_04654_),
    .X(_04760_));
 sg13g2_nand2_1 _18341_ (.Y(_04761_),
    .A(_04654_),
    .B(_04758_));
 sg13g2_o21ai_1 _18342_ (.B1(_04634_),
    .Y(_04762_),
    .A1(_04635_),
    .A2(_04636_));
 sg13g2_nand2_1 _18343_ (.Y(_04763_),
    .A(_04635_),
    .B(_04636_));
 sg13g2_a21o_1 _18344_ (.A2(_04635_),
    .A1(_04634_),
    .B1(_04636_),
    .X(_04764_));
 sg13g2_or2_1 _18345_ (.X(_04765_),
    .B(_04635_),
    .A(_04634_));
 sg13g2_nand4_1 _18346_ (.B(_04761_),
    .C(_04762_),
    .A(_04759_),
    .Y(_04766_),
    .D(_04763_));
 sg13g2_nand4_1 _18347_ (.B(_04760_),
    .C(_04764_),
    .A(_04758_),
    .Y(_04767_),
    .D(_04765_));
 sg13g2_and3_1 _18348_ (.X(_04768_),
    .A(_04757_),
    .B(_04766_),
    .C(_04767_));
 sg13g2_a21oi_1 _18349_ (.A1(_04766_),
    .A2(_04767_),
    .Y(_04769_),
    .B1(_04757_));
 sg13g2_or2_1 _18350_ (.X(_04770_),
    .B(_04769_),
    .A(_04768_));
 sg13g2_o21ai_1 _18351_ (.B1(_04659_),
    .Y(_04771_),
    .A1(_04768_),
    .A2(_04769_));
 sg13g2_or3_1 _18352_ (.A(_04659_),
    .B(_04768_),
    .C(_04769_),
    .X(_04772_));
 sg13g2_nand3_1 _18353_ (.B(_04771_),
    .C(_04772_),
    .A(_04752_),
    .Y(_04773_));
 sg13g2_a21o_1 _18354_ (.A2(_04772_),
    .A1(_04771_),
    .B1(_04752_),
    .X(_04774_));
 sg13g2_nand2_1 _18355_ (.Y(_04775_),
    .A(_04773_),
    .B(_04774_));
 sg13g2_nor2_1 _18356_ (.A(_04660_),
    .B(_04661_),
    .Y(_04776_));
 sg13g2_nand2_1 _18357_ (.Y(_04777_),
    .A(_04660_),
    .B(_04661_));
 sg13g2_a21o_1 _18358_ (.A2(_04777_),
    .A1(_04646_),
    .B1(_04776_),
    .X(_04778_));
 sg13g2_nand3_1 _18359_ (.B(_04774_),
    .C(_04778_),
    .A(_04773_),
    .Y(_04779_));
 sg13g2_a21oi_1 _18360_ (.A1(_04773_),
    .A2(_04774_),
    .Y(_04780_),
    .B1(_04778_));
 sg13g2_xnor2_1 _18361_ (.Y(_04781_),
    .A(_04775_),
    .B(_04778_));
 sg13g2_xor2_1 _18362_ (.B(_04781_),
    .A(_04728_),
    .X(_04782_));
 sg13g2_nand2_1 _18363_ (.Y(_04783_),
    .A(_04679_),
    .B(_04681_));
 sg13g2_o21ai_1 _18364_ (.B1(_04682_),
    .Y(_04784_),
    .A1(_04679_),
    .A2(_04681_));
 sg13g2_and2_1 _18365_ (.A(_04783_),
    .B(_04784_),
    .X(_04785_));
 sg13g2_a21oi_1 _18366_ (.A1(_04616_),
    .A2(_04617_),
    .Y(_04786_),
    .B1(_04615_));
 sg13g2_nor2_1 _18367_ (.A(_04616_),
    .B(_04617_),
    .Y(_04787_));
 sg13g2_nor2_1 _18368_ (.A(_04786_),
    .B(_04787_),
    .Y(_04788_));
 sg13g2_nand2_1 _18369_ (.Y(_04789_),
    .A(_09324_),
    .B(_07783_));
 sg13g2_o21ai_1 _18370_ (.B1(_04789_),
    .Y(_04790_),
    .A1(net7683),
    .A2(_08028_));
 sg13g2_and2_1 _18371_ (.A(_08239_),
    .B(_04790_),
    .X(_04791_));
 sg13g2_inv_1 _18372_ (.Y(_04792_),
    .A(_04791_));
 sg13g2_nor3_1 _18373_ (.A(_03628_),
    .B(_03821_),
    .C(_04792_),
    .Y(_04793_));
 sg13g2_nand3_1 _18374_ (.B(_03822_),
    .C(_04791_),
    .A(_03629_),
    .Y(_04794_));
 sg13g2_nor2_1 _18375_ (.A(net7243),
    .B(_04794_),
    .Y(_04795_));
 sg13g2_nand3_1 _18376_ (.B(_03629_),
    .C(_04790_),
    .A(_08249_),
    .Y(_04796_));
 sg13g2_nor2_1 _18377_ (.A(_03821_),
    .B(_04796_),
    .Y(_04797_));
 sg13g2_nand2b_1 _18378_ (.Y(_04798_),
    .B(_03822_),
    .A_N(_04796_));
 sg13g2_nor2_1 _18379_ (.A(net7243),
    .B(_04798_),
    .Y(_04799_));
 sg13g2_nor2_1 _18380_ (.A(net7237),
    .B(_04678_),
    .Y(_04800_));
 sg13g2_mux2_1 _18381_ (.A0(_04800_),
    .A1(net7237),
    .S(_04799_),
    .X(_04801_));
 sg13g2_xnor2_1 _18382_ (.Y(_04802_),
    .A(_04738_),
    .B(_04801_));
 sg13g2_xor2_1 _18383_ (.B(_04788_),
    .A(_04785_),
    .X(_04803_));
 sg13g2_xnor2_1 _18384_ (.Y(_04804_),
    .A(_04802_),
    .B(_04803_));
 sg13g2_o21ai_1 _18385_ (.B1(_04685_),
    .Y(_04805_),
    .A1(_04686_),
    .A2(_04687_));
 sg13g2_nor3_1 _18386_ (.A(_04685_),
    .B(_04686_),
    .C(_04687_),
    .Y(_04806_));
 sg13g2_o21ai_1 _18387_ (.B1(_04805_),
    .Y(_04807_),
    .A1(_04684_),
    .A2(_04806_));
 sg13g2_a22oi_1 _18388_ (.Y(_04808_),
    .B1(net7325),
    .B2(_01650_),
    .A2(_00538_),
    .A1(_01667_));
 sg13g2_nor2_1 _18389_ (.A(_04807_),
    .B(_04808_),
    .Y(_04809_));
 sg13g2_nand2_1 _18390_ (.Y(_04810_),
    .A(_04807_),
    .B(_04808_));
 sg13g2_nand2b_1 _18391_ (.Y(_04811_),
    .B(_04810_),
    .A_N(_04809_));
 sg13g2_xnor2_1 _18392_ (.Y(_04812_),
    .A(_04804_),
    .B(_04811_));
 sg13g2_a21oi_1 _18393_ (.A1(_04623_),
    .A2(_04628_),
    .Y(_04813_),
    .B1(_04629_));
 sg13g2_nand2_1 _18394_ (.Y(_04814_),
    .A(_04691_),
    .B(net6831));
 sg13g2_nor2_1 _18395_ (.A(_04691_),
    .B(net6831),
    .Y(_04815_));
 sg13g2_xnor2_1 _18396_ (.Y(_04816_),
    .A(_04691_),
    .B(_04813_));
 sg13g2_xnor2_1 _18397_ (.Y(_04817_),
    .A(_04812_),
    .B(_04816_));
 sg13g2_o21ai_1 _18398_ (.B1(_04663_),
    .Y(_04818_),
    .A1(_04631_),
    .A2(_04632_));
 sg13g2_nor3_1 _18399_ (.A(_04631_),
    .B(_04632_),
    .C(_04663_),
    .Y(_04819_));
 sg13g2_o21ai_1 _18400_ (.B1(_04818_),
    .Y(_04820_),
    .A1(_04568_),
    .A2(_04819_));
 sg13g2_nand2_1 _18401_ (.Y(_04821_),
    .A(net6741),
    .B(_04820_));
 sg13g2_nor2_1 _18402_ (.A(net6741),
    .B(_04820_),
    .Y(_04822_));
 sg13g2_xnor2_1 _18403_ (.Y(_04823_),
    .A(_04817_),
    .B(_04820_));
 sg13g2_xnor2_1 _18404_ (.Y(_04824_),
    .A(_04782_),
    .B(_04823_));
 sg13g2_o21ai_1 _18405_ (.B1(_04607_),
    .Y(_04825_),
    .A1(_04665_),
    .A2(_04696_));
 sg13g2_o21ai_1 _18406_ (.B1(_04693_),
    .Y(_04826_),
    .A1(_04668_),
    .A2(_04694_));
 sg13g2_and3_1 _18407_ (.X(_04827_),
    .A(_04697_),
    .B(_04825_),
    .C(_04826_));
 sg13g2_nand3_1 _18408_ (.B(_04825_),
    .C(_04826_),
    .A(_04697_),
    .Y(_04828_));
 sg13g2_a21oi_1 _18409_ (.A1(_04697_),
    .A2(_04825_),
    .Y(_04829_),
    .B1(_04826_));
 sg13g2_nor2_1 _18410_ (.A(_04827_),
    .B(_04829_),
    .Y(_04830_));
 sg13g2_xnor2_1 _18411_ (.Y(_04831_),
    .A(_04824_),
    .B(_04830_));
 sg13g2_nor2_1 _18412_ (.A(_04752_),
    .B(_04770_),
    .Y(_04832_));
 sg13g2_nand2_1 _18413_ (.Y(_04833_),
    .A(_04752_),
    .B(_04770_));
 sg13g2_a21oi_1 _18414_ (.A1(_04659_),
    .A2(_04833_),
    .Y(_04834_),
    .B1(_04832_));
 sg13g2_or2_1 _18415_ (.X(_04835_),
    .B(net7143),
    .A(net7222));
 sg13g2_a21o_1 _18416_ (.A2(_04743_),
    .A1(net7070),
    .B1(net7231),
    .X(_04836_));
 sg13g2_nand3_1 _18417_ (.B(net7231),
    .C(net7063),
    .A(net7070),
    .Y(_04837_));
 sg13g2_a21oi_1 _18418_ (.A1(_04836_),
    .A2(_04837_),
    .Y(_04838_),
    .B1(net7135));
 sg13g2_xnor2_1 _18419_ (.Y(_04839_),
    .A(_04835_),
    .B(_04838_));
 sg13g2_or2_1 _18420_ (.X(_04840_),
    .B(net7147),
    .A(net7212));
 sg13g2_or2_1 _18421_ (.X(_04841_),
    .B(net7163),
    .A(net7200));
 sg13g2_or2_1 _18422_ (.X(_04842_),
    .B(net7152),
    .A(net7210));
 sg13g2_xor2_1 _18423_ (.B(_04842_),
    .A(_04840_),
    .X(_04843_));
 sg13g2_xnor2_1 _18424_ (.Y(_04844_),
    .A(_04841_),
    .B(_04843_));
 sg13g2_nand2_1 _18425_ (.Y(_04845_),
    .A(net7065),
    .B(_04739_));
 sg13g2_nor2_1 _18426_ (.A(net7065),
    .B(_04739_),
    .Y(_04846_));
 sg13g2_nand3_1 _18427_ (.B(net7248),
    .C(_04742_),
    .A(net7637),
    .Y(_04847_));
 sg13g2_a21oi_1 _18428_ (.A1(_04845_),
    .A2(_04847_),
    .Y(_04848_),
    .B1(_04846_));
 sg13g2_or2_1 _18429_ (.X(_04849_),
    .B(_04848_),
    .A(_04844_));
 sg13g2_and2_1 _18430_ (.A(_04844_),
    .B(_04848_),
    .X(_04850_));
 sg13g2_xnor2_1 _18431_ (.Y(_04851_),
    .A(_04844_),
    .B(_04848_));
 sg13g2_xnor2_1 _18432_ (.Y(_04852_),
    .A(_04839_),
    .B(_04851_));
 sg13g2_xor2_1 _18433_ (.B(_04851_),
    .A(_04839_),
    .X(_04853_));
 sg13g2_mux2_1 _18434_ (.A0(_04847_),
    .A1(_04743_),
    .S(net7065),
    .X(_04854_));
 sg13g2_o21ai_1 _18435_ (.B1(net7071),
    .Y(_04855_),
    .A1(net7065),
    .A2(_04739_));
 sg13g2_o21ai_1 _18436_ (.B1(_04855_),
    .Y(_04856_),
    .A1(_04739_),
    .A2(_04854_));
 sg13g2_o21ai_1 _18437_ (.B1(_04733_),
    .Y(_04857_),
    .A1(_04747_),
    .A2(_04856_));
 sg13g2_nand3_1 _18438_ (.B(_04561_),
    .C(net7065),
    .A(net7231),
    .Y(_04858_));
 sg13g2_or2_1 _18439_ (.X(_04859_),
    .B(net7169),
    .A(net7194));
 sg13g2_or2_1 _18440_ (.X(_04860_),
    .B(net7182),
    .A(net7186));
 sg13g2_or2_1 _18441_ (.X(_04861_),
    .B(net7177),
    .A(net7189));
 sg13g2_xor2_1 _18442_ (.B(_04861_),
    .A(_04859_),
    .X(_04862_));
 sg13g2_xnor2_1 _18443_ (.Y(_04863_),
    .A(_04860_),
    .B(_04862_));
 sg13g2_nand2_1 _18444_ (.Y(_04864_),
    .A(_04730_),
    .B(_04731_));
 sg13g2_or2_1 _18445_ (.X(_04865_),
    .B(_04731_),
    .A(_04730_));
 sg13g2_o21ai_1 _18446_ (.B1(_04729_),
    .Y(_04866_),
    .A1(_04730_),
    .A2(_04731_));
 sg13g2_a21o_1 _18447_ (.A2(_04731_),
    .A1(_04730_),
    .B1(_04729_),
    .X(_04867_));
 sg13g2_nand2_1 _18448_ (.Y(_04868_),
    .A(_04754_),
    .B(_04755_));
 sg13g2_or2_1 _18449_ (.X(_04869_),
    .B(_04755_),
    .A(_04754_));
 sg13g2_o21ai_1 _18450_ (.B1(_04753_),
    .Y(_04870_),
    .A1(_04754_),
    .A2(_04755_));
 sg13g2_a21o_1 _18451_ (.A2(_04755_),
    .A1(_04754_),
    .B1(_04753_),
    .X(_04871_));
 sg13g2_nand4_1 _18452_ (.B(_04867_),
    .C(_04868_),
    .A(_04865_),
    .Y(_04872_),
    .D(_04870_));
 sg13g2_nand4_1 _18453_ (.B(_04866_),
    .C(_04869_),
    .A(_04864_),
    .Y(_04873_),
    .D(_04871_));
 sg13g2_nand3_1 _18454_ (.B(_04872_),
    .C(_04873_),
    .A(_04863_),
    .Y(_04874_));
 sg13g2_a21o_1 _18455_ (.A2(_04873_),
    .A1(_04872_),
    .B1(_04863_),
    .X(_04875_));
 sg13g2_a22oi_1 _18456_ (.Y(_04876_),
    .B1(_04874_),
    .B2(_04875_),
    .A2(_04858_),
    .A1(_04857_));
 sg13g2_and4_1 _18457_ (.A(_04857_),
    .B(_04858_),
    .C(_04874_),
    .D(_04875_),
    .X(_04877_));
 sg13g2_nand4_1 _18458_ (.B(_04858_),
    .C(_04874_),
    .A(_04857_),
    .Y(_04878_),
    .D(_04875_));
 sg13g2_nand3b_1 _18459_ (.B(_04878_),
    .C(_04852_),
    .Y(_04879_),
    .A_N(_04876_));
 sg13g2_o21ai_1 _18460_ (.B1(_04853_),
    .Y(_04880_),
    .A1(_04876_),
    .A2(_04877_));
 sg13g2_nor2_1 _18461_ (.A(net7206),
    .B(net7156),
    .Y(_04881_));
 sg13g2_nor2_1 _18462_ (.A(net7202),
    .B(net7159),
    .Y(_04882_));
 sg13g2_nor2_1 _18463_ (.A(net7196),
    .B(net7175),
    .Y(_04883_));
 sg13g2_xnor2_1 _18464_ (.Y(_04884_),
    .A(_04882_),
    .B(_04883_));
 sg13g2_xnor2_1 _18465_ (.Y(_04885_),
    .A(_04881_),
    .B(_04884_));
 sg13g2_nor2_1 _18466_ (.A(_04707_),
    .B(_04708_),
    .Y(_04886_));
 sg13g2_a21oi_1 _18467_ (.A1(_04707_),
    .A2(_04708_),
    .Y(_04887_),
    .B1(_04706_));
 sg13g2_nor2_1 _18468_ (.A(_04886_),
    .B(_04887_),
    .Y(_04888_));
 sg13g2_nor2_1 _18469_ (.A(net7227),
    .B(net7132),
    .Y(_04889_));
 sg13g2_nor2_1 _18470_ (.A(net7215),
    .B(net7148),
    .Y(_04890_));
 sg13g2_nor2_1 _18471_ (.A(net7219),
    .B(net7139),
    .Y(_04891_));
 sg13g2_xnor2_1 _18472_ (.Y(_04892_),
    .A(_04890_),
    .B(_04891_));
 sg13g2_xnor2_1 _18473_ (.Y(_04893_),
    .A(_04889_),
    .B(_04892_));
 sg13g2_nand2_1 _18474_ (.Y(_04894_),
    .A(_04888_),
    .B(_04893_));
 sg13g2_xor2_1 _18475_ (.B(_04893_),
    .A(_04888_),
    .X(_04895_));
 sg13g2_xnor2_1 _18476_ (.Y(_04896_),
    .A(_04885_),
    .B(_04895_));
 sg13g2_xor2_1 _18477_ (.B(_04895_),
    .A(_04885_),
    .X(_04897_));
 sg13g2_o21ai_1 _18478_ (.B1(_04710_),
    .Y(_04898_),
    .A1(_04713_),
    .A2(_04718_));
 sg13g2_a22oi_1 _18479_ (.Y(_04899_),
    .B1(_04764_),
    .B2(_04765_),
    .A2(_04761_),
    .A1(_04759_));
 sg13g2_nand4_1 _18480_ (.B(_04761_),
    .C(_04764_),
    .A(_04759_),
    .Y(_04900_),
    .D(_04765_));
 sg13g2_a21o_1 _18481_ (.A2(_04900_),
    .A1(_04757_),
    .B1(_04899_),
    .X(_04901_));
 sg13g2_a21oi_1 _18482_ (.A1(_04719_),
    .A2(_04898_),
    .Y(_04902_),
    .B1(_04901_));
 sg13g2_and3_1 _18483_ (.X(_04903_),
    .A(_04719_),
    .B(_04898_),
    .C(_04901_));
 sg13g2_nand3_1 _18484_ (.B(_04898_),
    .C(_04901_),
    .A(_04719_),
    .Y(_04904_));
 sg13g2_o21ai_1 _18485_ (.B1(_04896_),
    .Y(_04905_),
    .A1(_04902_),
    .A2(_04903_));
 sg13g2_or3_1 _18486_ (.A(_04896_),
    .B(_04902_),
    .C(_04903_),
    .X(_04906_));
 sg13g2_and4_1 _18487_ (.A(_04879_),
    .B(_04880_),
    .C(_04905_),
    .D(_04906_),
    .X(_04907_));
 sg13g2_nand4_1 _18488_ (.B(_04880_),
    .C(_04905_),
    .A(_04879_),
    .Y(_04908_),
    .D(_04906_));
 sg13g2_a22oi_1 _18489_ (.Y(_04909_),
    .B1(_04905_),
    .B2(_04906_),
    .A2(_04880_),
    .A1(_04879_));
 sg13g2_nor2_1 _18490_ (.A(_04907_),
    .B(_04909_),
    .Y(_04910_));
 sg13g2_xnor2_1 _18491_ (.Y(_04911_),
    .A(_04834_),
    .B(_04910_));
 sg13g2_o21ai_1 _18492_ (.B1(_04779_),
    .Y(_04912_),
    .A1(_04728_),
    .A2(_04780_));
 sg13g2_a21oi_1 _18493_ (.A1(_04804_),
    .A2(_04810_),
    .Y(_04913_),
    .B1(_04809_));
 sg13g2_a22oi_1 _18494_ (.Y(_04914_),
    .B1(_03818_),
    .B2(_01651_),
    .A2(_00538_),
    .A1(_01668_));
 sg13g2_xnor2_1 _18495_ (.Y(_04915_),
    .A(net7246),
    .B(net7240));
 sg13g2_nor2_1 _18496_ (.A(net7120),
    .B(_04915_),
    .Y(_04916_));
 sg13g2_nand2b_1 _18497_ (.Y(_04917_),
    .B(net7061),
    .A_N(_04915_));
 sg13g2_nor2_2 _18498_ (.A(net7116),
    .B(_04915_),
    .Y(_04918_));
 sg13g2_nand2b_1 _18499_ (.Y(_04919_),
    .B(_04797_),
    .A_N(_04915_));
 sg13g2_xnor2_1 _18500_ (.Y(_04920_),
    .A(_04914_),
    .B(_04918_));
 sg13g2_nor2_1 _18501_ (.A(_04715_),
    .B(_04716_),
    .Y(_04921_));
 sg13g2_a21oi_1 _18502_ (.A1(_04715_),
    .A2(_04716_),
    .Y(_04922_),
    .B1(_04714_));
 sg13g2_nor2_1 _18503_ (.A(_04921_),
    .B(_04922_),
    .Y(_04923_));
 sg13g2_nand2_1 _18504_ (.Y(_04924_),
    .A(net7237),
    .B(_04738_));
 sg13g2_nor2_1 _18505_ (.A(net7237),
    .B(_04738_),
    .Y(_04925_));
 sg13g2_a22oi_1 _18506_ (.Y(_04926_),
    .B1(_04925_),
    .B2(_04677_),
    .A2(_04924_),
    .A1(_04795_));
 sg13g2_a22oi_1 _18507_ (.Y(_04927_),
    .B1(_04924_),
    .B2(_04799_),
    .A2(_04800_),
    .A1(_04743_));
 sg13g2_nor2b_1 _18508_ (.A(_04923_),
    .B_N(_04926_),
    .Y(_04928_));
 sg13g2_o21ai_1 _18509_ (.B1(_04926_),
    .Y(_04929_),
    .A1(_04921_),
    .A2(_04922_));
 sg13g2_nor3_1 _18510_ (.A(_04921_),
    .B(_04922_),
    .C(_04927_),
    .Y(_04930_));
 sg13g2_xnor2_1 _18511_ (.Y(_04931_),
    .A(_04923_),
    .B(_04926_));
 sg13g2_xnor2_1 _18512_ (.Y(_04932_),
    .A(_04920_),
    .B(_04931_));
 sg13g2_nand2b_1 _18513_ (.Y(_04933_),
    .B(_04785_),
    .A_N(_04802_));
 sg13g2_nor2b_1 _18514_ (.A(_04785_),
    .B_N(_04802_),
    .Y(_04934_));
 sg13g2_a21o_1 _18515_ (.A2(_04933_),
    .A1(_04788_),
    .B1(_04934_),
    .X(_04935_));
 sg13g2_nand2b_1 _18516_ (.Y(_04936_),
    .B(_04935_),
    .A_N(_04932_));
 sg13g2_xor2_1 _18517_ (.B(_04935_),
    .A(_04932_),
    .X(_04937_));
 sg13g2_o21ai_1 _18518_ (.B1(_04726_),
    .Y(_04938_),
    .A1(_04721_),
    .A2(_04725_));
 sg13g2_xnor2_1 _18519_ (.Y(_04939_),
    .A(_04913_),
    .B(_04938_));
 sg13g2_xnor2_1 _18520_ (.Y(_04940_),
    .A(_04937_),
    .B(_04939_));
 sg13g2_nand2_1 _18521_ (.Y(_04941_),
    .A(_04912_),
    .B(_04940_));
 sg13g2_xnor2_1 _18522_ (.Y(_04942_),
    .A(_04912_),
    .B(_04940_));
 sg13g2_xnor2_1 _18523_ (.Y(_04943_),
    .A(_04911_),
    .B(_04942_));
 sg13g2_a21oi_1 _18524_ (.A1(_04812_),
    .A2(_04814_),
    .Y(_04944_),
    .B1(_04815_));
 sg13g2_inv_1 _18525_ (.Y(_04945_),
    .A(_04944_));
 sg13g2_a21oi_1 _18526_ (.A1(_04782_),
    .A2(_04821_),
    .Y(_04946_),
    .B1(_04822_));
 sg13g2_nand2_1 _18527_ (.Y(_04947_),
    .A(_04945_),
    .B(_04946_));
 sg13g2_xnor2_1 _18528_ (.Y(_04948_),
    .A(_04945_),
    .B(_04946_));
 sg13g2_xnor2_1 _18529_ (.Y(_04949_),
    .A(_04943_),
    .B(_04948_));
 sg13g2_or2_1 _18530_ (.X(_04950_),
    .B(net7134),
    .A(net7231));
 sg13g2_a21oi_1 _18531_ (.A1(_04835_),
    .A2(_04950_),
    .Y(_04951_),
    .B1(_03836_));
 sg13g2_nor2_1 _18532_ (.A(_04650_),
    .B(_04835_),
    .Y(_04952_));
 sg13g2_o21ai_1 _18533_ (.B1(net7063),
    .Y(_04953_),
    .A1(_04951_),
    .A2(_04952_));
 sg13g2_o21ai_1 _18534_ (.B1(_04953_),
    .Y(_04954_),
    .A1(_04835_),
    .A2(_04950_));
 sg13g2_nor2_1 _18535_ (.A(net7212),
    .B(net7140),
    .Y(_04955_));
 sg13g2_nor2_1 _18536_ (.A(net7222),
    .B(net7135),
    .Y(_04956_));
 sg13g2_xor2_1 _18537_ (.B(_04956_),
    .A(_04955_),
    .X(_04957_));
 sg13g2_nand2_1 _18538_ (.Y(_04958_),
    .A(net7231),
    .B(_04743_));
 sg13g2_xnor2_1 _18539_ (.Y(_04959_),
    .A(_04957_),
    .B(_04958_));
 sg13g2_nor2_1 _18540_ (.A(net7210),
    .B(net7147),
    .Y(_04960_));
 sg13g2_nor2_1 _18541_ (.A(net7193),
    .B(net7163),
    .Y(_04961_));
 sg13g2_nor2_1 _18542_ (.A(net7200),
    .B(net7152),
    .Y(_04962_));
 sg13g2_xnor2_1 _18543_ (.Y(_04963_),
    .A(_04961_),
    .B(_04962_));
 sg13g2_xnor2_1 _18544_ (.Y(_04964_),
    .A(_04960_),
    .B(_04963_));
 sg13g2_xor2_1 _18545_ (.B(_04964_),
    .A(_04959_),
    .X(_04965_));
 sg13g2_xnor2_1 _18546_ (.Y(_04966_),
    .A(_04954_),
    .B(_04965_));
 sg13g2_nor2_1 _18547_ (.A(net7190),
    .B(net7169),
    .Y(_04967_));
 sg13g2_nor2_1 _18548_ (.A(net7182),
    .B(net7177),
    .Y(_04968_));
 sg13g2_nor2_1 _18549_ (.A(net7186),
    .B(net7175),
    .Y(_04969_));
 sg13g2_xnor2_1 _18550_ (.Y(_04970_),
    .A(_04968_),
    .B(_04969_));
 sg13g2_xnor2_1 _18551_ (.Y(_04971_),
    .A(_04967_),
    .B(_04970_));
 sg13g2_or2_1 _18552_ (.X(_04972_),
    .B(_04842_),
    .A(_04841_));
 sg13g2_a21o_1 _18553_ (.A2(_04842_),
    .A1(_04841_),
    .B1(_04840_),
    .X(_04973_));
 sg13g2_nand2_1 _18554_ (.Y(_04974_),
    .A(_04972_),
    .B(_04973_));
 sg13g2_or2_1 _18555_ (.X(_04975_),
    .B(_04861_),
    .A(_04860_));
 sg13g2_a21o_1 _18556_ (.A2(_04861_),
    .A1(_04860_),
    .B1(_04859_),
    .X(_04976_));
 sg13g2_nand2_1 _18557_ (.Y(_04977_),
    .A(_04975_),
    .B(_04976_));
 sg13g2_xor2_1 _18558_ (.B(_04977_),
    .A(_04974_),
    .X(_04978_));
 sg13g2_xnor2_1 _18559_ (.Y(_04979_),
    .A(_04971_),
    .B(_04978_));
 sg13g2_a21oi_1 _18560_ (.A1(_04839_),
    .A2(_04849_),
    .Y(_04980_),
    .B1(_04850_));
 sg13g2_nand2_1 _18561_ (.Y(_04981_),
    .A(_04979_),
    .B(_04980_));
 sg13g2_xor2_1 _18562_ (.B(_04980_),
    .A(_04979_),
    .X(_04982_));
 sg13g2_xnor2_1 _18563_ (.Y(_04983_),
    .A(_04966_),
    .B(_04982_));
 sg13g2_o21ai_1 _18564_ (.B1(_04878_),
    .Y(_04984_),
    .A1(_04852_),
    .A2(_04876_));
 sg13g2_nor2_1 _18565_ (.A(net7206),
    .B(net7148),
    .Y(_04985_));
 sg13g2_nor2_1 _18566_ (.A(net7196),
    .B(net7159),
    .Y(_04986_));
 sg13g2_nor2_1 _18567_ (.A(net7202),
    .B(net7156),
    .Y(_04987_));
 sg13g2_xnor2_1 _18568_ (.Y(_04988_),
    .A(_04986_),
    .B(_04987_));
 sg13g2_xnor2_1 _18569_ (.Y(_04989_),
    .A(_04985_),
    .B(_04988_));
 sg13g2_a21oi_1 _18570_ (.A1(_04881_),
    .A2(_04883_),
    .Y(_04990_),
    .B1(_04882_));
 sg13g2_nor2_1 _18571_ (.A(_04881_),
    .B(_04883_),
    .Y(_04991_));
 sg13g2_nor2_1 _18572_ (.A(_04990_),
    .B(_04991_),
    .Y(_04992_));
 sg13g2_nor2_1 _18573_ (.A(net7219),
    .B(net7132),
    .Y(_04993_));
 sg13g2_nor2_1 _18574_ (.A(net7215),
    .B(net7137),
    .Y(_04994_));
 sg13g2_nor2_1 _18575_ (.A(net7227),
    .B(net7116),
    .Y(_04995_));
 sg13g2_xnor2_1 _18576_ (.Y(_04996_),
    .A(_04993_),
    .B(_04995_));
 sg13g2_xnor2_1 _18577_ (.Y(_04997_),
    .A(_04994_),
    .B(_04996_));
 sg13g2_nor2_1 _18578_ (.A(_04992_),
    .B(_04997_),
    .Y(_04998_));
 sg13g2_xnor2_1 _18579_ (.Y(_04999_),
    .A(_04992_),
    .B(_04997_));
 sg13g2_xnor2_1 _18580_ (.Y(_05000_),
    .A(_04989_),
    .B(_04999_));
 sg13g2_o21ai_1 _18581_ (.B1(_04885_),
    .Y(_05001_),
    .A1(_04888_),
    .A2(_04893_));
 sg13g2_nand4_1 _18582_ (.B(_04866_),
    .C(_04868_),
    .A(_04864_),
    .Y(_05002_),
    .D(_04870_));
 sg13g2_a22oi_1 _18583_ (.Y(_05003_),
    .B1(_04868_),
    .B2(_04870_),
    .A2(_04866_),
    .A1(_04864_));
 sg13g2_o21ai_1 _18584_ (.B1(_05002_),
    .Y(_05004_),
    .A1(_04863_),
    .A2(_05003_));
 sg13g2_and3_1 _18585_ (.X(_05005_),
    .A(_04894_),
    .B(_05001_),
    .C(_05004_));
 sg13g2_nand3_1 _18586_ (.B(_05001_),
    .C(_05004_),
    .A(_04894_),
    .Y(_05006_));
 sg13g2_a21oi_1 _18587_ (.A1(_04894_),
    .A2(_05001_),
    .Y(_05007_),
    .B1(_05004_));
 sg13g2_nor2_1 _18588_ (.A(_05005_),
    .B(_05007_),
    .Y(_05008_));
 sg13g2_xnor2_1 _18589_ (.Y(_05009_),
    .A(_05000_),
    .B(_05008_));
 sg13g2_xnor2_1 _18590_ (.Y(_05010_),
    .A(_04984_),
    .B(_05009_));
 sg13g2_xor2_1 _18591_ (.B(_05010_),
    .A(_04983_),
    .X(_05011_));
 sg13g2_o21ai_1 _18592_ (.B1(_04908_),
    .Y(_05012_),
    .A1(_04834_),
    .A2(_04909_));
 sg13g2_nand2_1 _18593_ (.Y(_05013_),
    .A(_04890_),
    .B(_04891_));
 sg13g2_o21ai_1 _18594_ (.B1(_04889_),
    .Y(_05014_),
    .A1(_04890_),
    .A2(_04891_));
 sg13g2_nand2_1 _18595_ (.Y(_05015_),
    .A(_05013_),
    .B(_05014_));
 sg13g2_and3_1 _18596_ (.X(_05016_),
    .A(_01668_),
    .B(_00538_),
    .C(_04791_));
 sg13g2_a21oi_1 _18597_ (.A1(_01652_),
    .A2(net7325),
    .Y(_05017_),
    .B1(_05016_));
 sg13g2_and4_1 _18598_ (.A(_01668_),
    .B(_00538_),
    .C(_08249_),
    .D(_04790_),
    .X(_05018_));
 sg13g2_inv_1 _18599_ (.Y(_05019_),
    .A(net7314));
 sg13g2_a21oi_1 _18600_ (.A1(_01652_),
    .A2(net7320),
    .Y(_05020_),
    .B1(net7315));
 sg13g2_nand3_1 _18601_ (.B(_05014_),
    .C(_05017_),
    .A(_05013_),
    .Y(_05021_));
 sg13g2_xnor2_1 _18602_ (.Y(_05022_),
    .A(_05015_),
    .B(_05017_));
 sg13g2_nor2_1 _18603_ (.A(_04914_),
    .B(_04918_),
    .Y(_05023_));
 sg13g2_nor2_1 _18604_ (.A(net7245),
    .B(net7240),
    .Y(_05024_));
 sg13g2_nor3_1 _18605_ (.A(net7245),
    .B(net7237),
    .C(_04794_),
    .Y(_05025_));
 sg13g2_nor3_1 _18606_ (.A(net7245),
    .B(net7240),
    .C(_04798_),
    .Y(_05026_));
 sg13g2_nand2_1 _18607_ (.Y(_05027_),
    .A(_04797_),
    .B(_05024_));
 sg13g2_and2_1 _18608_ (.A(_04914_),
    .B(net7004),
    .X(_05028_));
 sg13g2_a21oi_1 _18609_ (.A1(_04914_),
    .A2(_04918_),
    .Y(_05029_),
    .B1(_04927_));
 sg13g2_o21ai_1 _18610_ (.B1(_04923_),
    .Y(_05030_),
    .A1(_05023_),
    .A2(_05029_));
 sg13g2_nand2b_1 _18611_ (.Y(_05031_),
    .B(_05023_),
    .A_N(_04927_));
 sg13g2_a21oi_1 _18612_ (.A1(_05030_),
    .A2(_05031_),
    .Y(_05032_),
    .B1(net7053));
 sg13g2_o21ai_1 _18613_ (.B1(_04929_),
    .Y(_05033_),
    .A1(_04920_),
    .A2(_04930_));
 sg13g2_a221oi_1 _18614_ (.B2(net7053),
    .C1(_05032_),
    .B1(_05033_),
    .A1(_04928_),
    .Y(_05034_),
    .A2(_05028_));
 sg13g2_xnor2_1 _18615_ (.Y(_05035_),
    .A(_05022_),
    .B(_05034_));
 sg13g2_o21ai_1 _18616_ (.B1(_04904_),
    .Y(_05036_),
    .A1(_04897_),
    .A2(_04902_));
 sg13g2_xnor2_1 _18617_ (.Y(_05037_),
    .A(_04936_),
    .B(_05036_));
 sg13g2_xnor2_1 _18618_ (.Y(_05038_),
    .A(_05035_),
    .B(_05037_));
 sg13g2_nor2_1 _18619_ (.A(_05012_),
    .B(_05038_),
    .Y(_05039_));
 sg13g2_nand2_1 _18620_ (.Y(_05040_),
    .A(_05012_),
    .B(_05038_));
 sg13g2_nand2b_1 _18621_ (.Y(_05041_),
    .B(_05040_),
    .A_N(_05039_));
 sg13g2_xor2_1 _18622_ (.B(_05041_),
    .A(_05011_),
    .X(_05042_));
 sg13g2_o21ai_1 _18623_ (.B1(_04911_),
    .Y(_05043_),
    .A1(_04912_),
    .A2(_04940_));
 sg13g2_nand2_1 _18624_ (.Y(_05044_),
    .A(_04941_),
    .B(_05043_));
 sg13g2_nand2_1 _18625_ (.Y(_05045_),
    .A(_04913_),
    .B(_04937_));
 sg13g2_nor2_1 _18626_ (.A(_04913_),
    .B(_04937_),
    .Y(_05046_));
 sg13g2_a21oi_1 _18627_ (.A1(_04938_),
    .A2(_05045_),
    .Y(_05047_),
    .B1(_05046_));
 sg13g2_a21oi_1 _18628_ (.A1(_04941_),
    .A2(_05043_),
    .Y(_05048_),
    .B1(_05047_));
 sg13g2_nand3_1 _18629_ (.B(_05043_),
    .C(_05047_),
    .A(_04941_),
    .Y(_05049_));
 sg13g2_xnor2_1 _18630_ (.Y(_05050_),
    .A(_05042_),
    .B(_05047_));
 sg13g2_xor2_1 _18631_ (.B(_05050_),
    .A(_05044_),
    .X(_05051_));
 sg13g2_nor2_1 _18632_ (.A(net7210),
    .B(net7140),
    .Y(_05052_));
 sg13g2_nor2_1 _18633_ (.A(net7212),
    .B(net7135),
    .Y(_05053_));
 sg13g2_xnor2_1 _18634_ (.Y(_05054_),
    .A(_05052_),
    .B(_05053_));
 sg13g2_nand2_1 _18635_ (.Y(_05055_),
    .A(net7222),
    .B(net7064));
 sg13g2_xnor2_1 _18636_ (.Y(_05056_),
    .A(_05054_),
    .B(_05055_));
 sg13g2_nor2_1 _18637_ (.A(_04955_),
    .B(_04956_),
    .Y(_05057_));
 sg13g2_a22oi_1 _18638_ (.Y(_05058_),
    .B1(_04955_),
    .B2(_04956_),
    .A2(net7064),
    .A1(net7231));
 sg13g2_or2_1 _18639_ (.X(_05059_),
    .B(_05058_),
    .A(_05057_));
 sg13g2_or2_1 _18640_ (.X(_05060_),
    .B(net7147),
    .A(net7200));
 sg13g2_or2_1 _18641_ (.X(_05061_),
    .B(net7163),
    .A(net7189));
 sg13g2_or2_1 _18642_ (.X(_05062_),
    .B(net7152),
    .A(_04041_));
 sg13g2_xnor2_1 _18643_ (.Y(_05063_),
    .A(_05060_),
    .B(_05062_));
 sg13g2_xnor2_1 _18644_ (.Y(_05064_),
    .A(_05061_),
    .B(_05063_));
 sg13g2_xor2_1 _18645_ (.B(_05064_),
    .A(_05059_),
    .X(_05065_));
 sg13g2_xnor2_1 _18646_ (.Y(_05066_),
    .A(_05056_),
    .B(_05065_));
 sg13g2_and2_1 _18647_ (.A(_04959_),
    .B(_04964_),
    .X(_05067_));
 sg13g2_or2_1 _18648_ (.X(_05068_),
    .B(_04964_),
    .A(_04959_));
 sg13g2_a21oi_1 _18649_ (.A1(_04954_),
    .A2(_05068_),
    .Y(_05069_),
    .B1(_05067_));
 sg13g2_nor2_1 _18650_ (.A(net7186),
    .B(net7159),
    .Y(_05070_));
 sg13g2_nor2_1 _18651_ (.A(net7177),
    .B(net7175),
    .Y(_05071_));
 sg13g2_nor2_1 _18652_ (.A(net7183),
    .B(net7169),
    .Y(_05072_));
 sg13g2_xnor2_1 _18653_ (.Y(_05073_),
    .A(_05070_),
    .B(_05072_));
 sg13g2_xnor2_1 _18654_ (.Y(_05074_),
    .A(_05071_),
    .B(_05073_));
 sg13g2_nor2_1 _18655_ (.A(_04961_),
    .B(_04962_),
    .Y(_05075_));
 sg13g2_a21oi_1 _18656_ (.A1(_04961_),
    .A2(_04962_),
    .Y(_05076_),
    .B1(_04960_));
 sg13g2_nor2_1 _18657_ (.A(_05075_),
    .B(_05076_),
    .Y(_05077_));
 sg13g2_nor2_1 _18658_ (.A(_04968_),
    .B(_04969_),
    .Y(_05078_));
 sg13g2_a21oi_1 _18659_ (.A1(_04968_),
    .A2(_04969_),
    .Y(_05079_),
    .B1(_04967_));
 sg13g2_nor2_1 _18660_ (.A(_05078_),
    .B(_05079_),
    .Y(_05080_));
 sg13g2_xor2_1 _18661_ (.B(_05080_),
    .A(_05077_),
    .X(_05081_));
 sg13g2_xnor2_1 _18662_ (.Y(_05082_),
    .A(_05074_),
    .B(_05081_));
 sg13g2_nor2_1 _18663_ (.A(_05069_),
    .B(_05082_),
    .Y(_05083_));
 sg13g2_nand2_1 _18664_ (.Y(_05084_),
    .A(_05069_),
    .B(_05082_));
 sg13g2_nand2b_1 _18665_ (.Y(_05085_),
    .B(_05084_),
    .A_N(_05083_));
 sg13g2_xnor2_1 _18666_ (.Y(_05086_),
    .A(_05066_),
    .B(_05085_));
 sg13g2_o21ai_1 _18667_ (.B1(_04966_),
    .Y(_05087_),
    .A1(_04979_),
    .A2(_04980_));
 sg13g2_nand2_1 _18668_ (.Y(_05088_),
    .A(_04981_),
    .B(_05087_));
 sg13g2_nand3b_1 _18669_ (.B(_04677_),
    .C(net7219),
    .Y(_05089_),
    .A_N(net7216));
 sg13g2_nand2b_1 _18670_ (.Y(_05090_),
    .B(net7216),
    .A_N(net7219));
 sg13g2_o21ai_1 _18671_ (.B1(net7220),
    .Y(_05091_),
    .A1(_03904_),
    .A2(_04678_));
 sg13g2_nor2_1 _18672_ (.A(net7220),
    .B(net7216),
    .Y(_05092_));
 sg13g2_and2_1 _18673_ (.A(_05089_),
    .B(_05090_),
    .X(_05093_));
 sg13g2_nor3_1 _18674_ (.A(net7216),
    .B(net7130),
    .C(net7118),
    .Y(_05094_));
 sg13g2_o21ai_1 _18675_ (.B1(_05089_),
    .Y(_05095_),
    .A1(net7116),
    .A2(_05090_));
 sg13g2_a221oi_1 _18676_ (.B2(net7227),
    .C1(_05094_),
    .B1(_05095_),
    .A1(_04995_),
    .Y(_05096_),
    .A2(_05093_));
 sg13g2_nor2_1 _18677_ (.A(_04986_),
    .B(_04987_),
    .Y(_05097_));
 sg13g2_a21oi_1 _18678_ (.A1(_04986_),
    .A2(_04987_),
    .Y(_05098_),
    .B1(_04985_));
 sg13g2_nor2_1 _18679_ (.A(_05097_),
    .B(_05098_),
    .Y(_05099_));
 sg13g2_or2_1 _18680_ (.X(_05100_),
    .B(net7137),
    .A(net7206));
 sg13g2_nor2_1 _18681_ (.A(net7196),
    .B(net7158),
    .Y(_05101_));
 sg13g2_nor2_1 _18682_ (.A(net7202),
    .B(net7149),
    .Y(_05102_));
 sg13g2_xnor2_1 _18683_ (.Y(_05103_),
    .A(_05101_),
    .B(_05102_));
 sg13g2_xnor2_1 _18684_ (.Y(_05104_),
    .A(_05100_),
    .B(_05103_));
 sg13g2_nand2b_1 _18685_ (.Y(_05105_),
    .B(_05099_),
    .A_N(_05104_));
 sg13g2_nor2b_1 _18686_ (.A(_05099_),
    .B_N(_05104_),
    .Y(_05106_));
 sg13g2_xnor2_1 _18687_ (.Y(_05107_),
    .A(_05099_),
    .B(_05104_));
 sg13g2_xnor2_1 _18688_ (.Y(_05108_),
    .A(_05096_),
    .B(_05107_));
 sg13g2_nand4_1 _18689_ (.B(_04973_),
    .C(_04975_),
    .A(_04972_),
    .Y(_05109_),
    .D(_04976_));
 sg13g2_a22oi_1 _18690_ (.Y(_05110_),
    .B1(_04975_),
    .B2(_04976_),
    .A2(_04973_),
    .A1(_04972_));
 sg13g2_o21ai_1 _18691_ (.B1(_05109_),
    .Y(_05111_),
    .A1(_04971_),
    .A2(_05110_));
 sg13g2_a21oi_1 _18692_ (.A1(_04992_),
    .A2(_04997_),
    .Y(_05112_),
    .B1(_04989_));
 sg13g2_inv_1 _18693_ (.Y(_05113_),
    .A(_00556_));
 sg13g2_nor3_1 _18694_ (.A(_04998_),
    .B(_05111_),
    .C(_05112_),
    .Y(_05114_));
 sg13g2_o21ai_1 _18695_ (.B1(_05111_),
    .Y(_05115_),
    .A1(_04998_),
    .A2(_05112_));
 sg13g2_nand2b_1 _18696_ (.Y(_05116_),
    .B(_05115_),
    .A_N(_05114_));
 sg13g2_xnor2_1 _18697_ (.Y(_05117_),
    .A(_05108_),
    .B(_05116_));
 sg13g2_nor2b_1 _18698_ (.A(_05088_),
    .B_N(_05117_),
    .Y(_05118_));
 sg13g2_a21o_1 _18699_ (.A2(_05087_),
    .A1(_04981_),
    .B1(_05117_),
    .X(_05119_));
 sg13g2_xnor2_1 _18700_ (.Y(_05120_),
    .A(_05088_),
    .B(_05117_));
 sg13g2_xnor2_1 _18701_ (.Y(_05121_),
    .A(_05086_),
    .B(_05120_));
 sg13g2_nor2_1 _18702_ (.A(_04984_),
    .B(_05009_),
    .Y(_05122_));
 sg13g2_nand2_1 _18703_ (.Y(_05123_),
    .A(_04984_),
    .B(_05009_));
 sg13g2_a21oi_1 _18704_ (.A1(_04983_),
    .A2(_05123_),
    .Y(_05124_),
    .B1(_05122_));
 sg13g2_nor2_1 _18705_ (.A(_04917_),
    .B(_05017_),
    .Y(_05125_));
 sg13g2_or2_1 _18706_ (.X(_05126_),
    .B(_05125_),
    .A(_05025_));
 sg13g2_nor2_1 _18707_ (.A(_04993_),
    .B(_04994_),
    .Y(_05127_));
 sg13g2_a21oi_1 _18708_ (.A1(_04993_),
    .A2(_04994_),
    .Y(_05128_),
    .B1(_04995_));
 sg13g2_nor2_1 _18709_ (.A(_05127_),
    .B(_05128_),
    .Y(_05129_));
 sg13g2_a21oi_1 _18710_ (.A1(_01653_),
    .A2(net7325),
    .Y(_05130_),
    .B1(_05016_));
 sg13g2_xnor2_1 _18711_ (.Y(_05131_),
    .A(_04916_),
    .B(_05130_));
 sg13g2_and2_1 _18712_ (.A(_05129_),
    .B(_05131_),
    .X(_05132_));
 sg13g2_inv_1 _18713_ (.Y(_05133_),
    .A(_05132_));
 sg13g2_a21oi_1 _18714_ (.A1(_01653_),
    .A2(net7320),
    .Y(_05134_),
    .B1(net7315));
 sg13g2_xnor2_1 _18715_ (.Y(_05135_),
    .A(net7004),
    .B(_05134_));
 sg13g2_nor2_1 _18716_ (.A(_05129_),
    .B(_05135_),
    .Y(_05136_));
 sg13g2_nor2_1 _18717_ (.A(_05132_),
    .B(_05136_),
    .Y(_05137_));
 sg13g2_nor2_1 _18718_ (.A(_04919_),
    .B(_05020_),
    .Y(_05138_));
 sg13g2_nor2_1 _18719_ (.A(net7053),
    .B(_05138_),
    .Y(_05139_));
 sg13g2_o21ai_1 _18720_ (.B1(_05027_),
    .Y(_05140_),
    .A1(_04919_),
    .A2(_05020_));
 sg13g2_xnor2_1 _18721_ (.Y(_05141_),
    .A(_05126_),
    .B(_05137_));
 sg13g2_nand2_1 _18722_ (.Y(_05142_),
    .A(_04914_),
    .B(_05027_));
 sg13g2_nor2_1 _18723_ (.A(_05015_),
    .B(_05142_),
    .Y(_05143_));
 sg13g2_nand2_1 _18724_ (.Y(_05144_),
    .A(_05015_),
    .B(_05142_));
 sg13g2_a21oi_1 _18725_ (.A1(_05013_),
    .A2(_05014_),
    .Y(_05145_),
    .B1(_05017_));
 sg13g2_o21ai_1 _18726_ (.B1(_05021_),
    .Y(_05146_),
    .A1(_05025_),
    .A2(_05145_));
 sg13g2_a221oi_1 _18727_ (.B2(_04917_),
    .C1(_05143_),
    .B1(_05146_),
    .A1(_05125_),
    .Y(_05147_),
    .A2(_05144_));
 sg13g2_nand2_1 _18728_ (.Y(_05148_),
    .A(_05015_),
    .B(net7053));
 sg13g2_nand2_1 _18729_ (.Y(_05149_),
    .A(_05020_),
    .B(_05148_));
 sg13g2_o21ai_1 _18730_ (.B1(_05149_),
    .Y(_05150_),
    .A1(_05015_),
    .A2(net7053));
 sg13g2_a221oi_1 _18731_ (.B2(_04919_),
    .C1(_05143_),
    .B1(_05150_),
    .A1(_05125_),
    .Y(_05151_),
    .A2(_05144_));
 sg13g2_xnor2_1 _18732_ (.Y(_05152_),
    .A(_05141_),
    .B(_05151_));
 sg13g2_a21oi_1 _18733_ (.A1(_05000_),
    .A2(_05006_),
    .Y(_05153_),
    .B1(_05007_));
 sg13g2_a21o_1 _18734_ (.A2(net7005),
    .A1(_04914_),
    .B1(_05025_),
    .X(_05154_));
 sg13g2_a21oi_1 _18735_ (.A1(_05022_),
    .A2(_05154_),
    .Y(_05155_),
    .B1(_05033_));
 sg13g2_o21ai_1 _18736_ (.B1(_05155_),
    .Y(_05156_),
    .A1(_05022_),
    .A2(_05154_));
 sg13g2_nand2_1 _18737_ (.Y(_05157_),
    .A(_05153_),
    .B(_05156_));
 sg13g2_xor2_1 _18738_ (.B(_05156_),
    .A(_05153_),
    .X(_05158_));
 sg13g2_inv_1 _18739_ (.Y(_05159_),
    .A(_00544_));
 sg13g2_xnor2_1 _18740_ (.Y(_05160_),
    .A(_05152_),
    .B(_05158_));
 sg13g2_nand2_1 _18741_ (.Y(_05161_),
    .A(_05124_),
    .B(_05160_));
 sg13g2_inv_1 _18742_ (.Y(_05162_),
    .A(_00543_));
 sg13g2_xnor2_1 _18743_ (.Y(_05163_),
    .A(_05124_),
    .B(_05160_));
 sg13g2_xnor2_1 _18744_ (.Y(_05164_),
    .A(_05121_),
    .B(_05163_));
 sg13g2_a21oi_1 _18745_ (.A1(_05011_),
    .A2(_05040_),
    .Y(_05165_),
    .B1(_05039_));
 sg13g2_nand2b_1 _18746_ (.Y(_05166_),
    .B(_05035_),
    .A_N(_05036_));
 sg13g2_nor2b_1 _18747_ (.A(_05035_),
    .B_N(_05036_),
    .Y(_05167_));
 sg13g2_o21ai_1 _18748_ (.B1(_05166_),
    .Y(_05168_),
    .A1(_04936_),
    .A2(_05167_));
 sg13g2_nor2_1 _18749_ (.A(_05165_),
    .B(_05168_),
    .Y(_05169_));
 sg13g2_nand2_1 _18750_ (.Y(_05170_),
    .A(_05165_),
    .B(_05168_));
 sg13g2_nor2b_1 _18751_ (.A(_05169_),
    .B_N(_05170_),
    .Y(_05171_));
 sg13g2_xnor2_1 _18752_ (.Y(_05172_),
    .A(_05164_),
    .B(_05171_));
 sg13g2_a21oi_1 _18753_ (.A1(_05108_),
    .A2(_05115_),
    .Y(_05173_),
    .B1(_05114_));
 sg13g2_inv_1 _18754_ (.Y(_05174_),
    .A(_00540_));
 sg13g2_o21ai_1 _18755_ (.B1(net7228),
    .Y(_05175_),
    .A1(net7220),
    .A2(net7215));
 sg13g2_nand3_1 _18756_ (.B(_05091_),
    .C(_05175_),
    .A(net7061),
    .Y(_05176_));
 sg13g2_a21oi_1 _18757_ (.A1(_01654_),
    .A2(net7325),
    .Y(_05177_),
    .B1(_05016_));
 sg13g2_a21oi_1 _18758_ (.A1(net7005),
    .A2(_05130_),
    .Y(_05178_),
    .B1(net7059));
 sg13g2_xnor2_1 _18759_ (.Y(_05179_),
    .A(_05177_),
    .B(_05178_));
 sg13g2_inv_1 _18760_ (.Y(_05180_),
    .A(_00539_));
 sg13g2_xnor2_1 _18761_ (.Y(_05181_),
    .A(net6992),
    .B(_05179_));
 sg13g2_a21oi_1 _18762_ (.A1(_03863_),
    .A2(_05091_),
    .Y(_05182_),
    .B1(_05092_));
 sg13g2_a21o_1 _18763_ (.A2(_05091_),
    .A1(_03863_),
    .B1(_05092_),
    .X(_05183_));
 sg13g2_nor2_1 _18764_ (.A(_04798_),
    .B(_05182_),
    .Y(_05184_));
 sg13g2_nand2_1 _18765_ (.Y(_05185_),
    .A(net7119),
    .B(_05183_));
 sg13g2_inv_1 _18766_ (.Y(_05186_),
    .A(_00005_));
 sg13g2_a21oi_1 _18767_ (.A1(_01654_),
    .A2(net7320),
    .Y(_05187_),
    .B1(net7315));
 sg13g2_a21o_1 _18768_ (.A2(net7320),
    .A1(_01654_),
    .B1(net7315),
    .X(_05188_));
 sg13g2_a21oi_1 _18769_ (.A1(net7004),
    .A2(_05134_),
    .Y(_05189_),
    .B1(_05026_));
 sg13g2_xnor2_1 _18770_ (.Y(_05190_),
    .A(_05187_),
    .B(_05189_));
 sg13g2_xnor2_1 _18771_ (.Y(_05191_),
    .A(_05184_),
    .B(_05190_));
 sg13g2_xnor2_1 _18772_ (.Y(_05192_),
    .A(_05173_),
    .B(_05191_));
 sg13g2_and3_1 _18773_ (.X(_05193_),
    .A(_05126_),
    .B(_05129_),
    .C(_05131_));
 sg13g2_a22oi_1 _18774_ (.Y(_05194_),
    .B1(_05147_),
    .B2(_05193_),
    .A2(_05139_),
    .A1(_05136_));
 sg13g2_inv_1 _18775_ (.Y(_05195_),
    .A(_00536_));
 sg13g2_a21oi_1 _18776_ (.A1(_05129_),
    .A2(_05135_),
    .Y(_05196_),
    .B1(_05140_));
 sg13g2_inv_1 _18777_ (.Y(_05197_),
    .A(_05198_));
 sg13g2_or2_1 _18778_ (.X(_05198_),
    .B(_05196_),
    .A(_05136_));
 sg13g2_inv_1 _18779_ (.Y(_05199_),
    .A(_00534_));
 sg13g2_o21ai_1 _18780_ (.B1(_05194_),
    .Y(_05200_),
    .A1(_05151_),
    .A2(_05197_));
 sg13g2_inv_1 _18781_ (.Y(_05201_),
    .A(_00533_));
 sg13g2_xor2_1 _18782_ (.B(_05200_),
    .A(_05192_),
    .X(_05202_));
 sg13g2_nor2_1 _18783_ (.A(net7206),
    .B(net7130),
    .Y(_05203_));
 sg13g2_nor2_1 _18784_ (.A(net7196),
    .B(net7150),
    .Y(_05204_));
 sg13g2_nor2_1 _18785_ (.A(net7203),
    .B(net7137),
    .Y(_05205_));
 sg13g2_xnor2_1 _18786_ (.Y(_05206_),
    .A(_05204_),
    .B(_05205_));
 sg13g2_xnor2_1 _18787_ (.Y(_05207_),
    .A(_05203_),
    .B(_05206_));
 sg13g2_nand2_1 _18788_ (.Y(_05208_),
    .A(_05101_),
    .B(_05102_));
 sg13g2_nor2_1 _18789_ (.A(_05101_),
    .B(_05102_),
    .Y(_05209_));
 sg13g2_o21ai_1 _18790_ (.B1(_05208_),
    .Y(_05210_),
    .A1(_05100_),
    .A2(_05209_));
 sg13g2_nand2_1 _18791_ (.Y(_05211_),
    .A(_05207_),
    .B(_05210_));
 sg13g2_xor2_1 _18792_ (.B(_05210_),
    .A(_05207_),
    .X(_05212_));
 sg13g2_inv_1 _18793_ (.Y(_05213_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_by_zero_q ));
 sg13g2_nand3_1 _18794_ (.B(_05089_),
    .C(_05090_),
    .A(_03863_),
    .Y(_05214_));
 sg13g2_xor2_1 _18795_ (.B(net7216),
    .A(net7219),
    .X(_05215_));
 sg13g2_nand2_1 _18796_ (.Y(_05216_),
    .A(net7227),
    .B(_05215_));
 sg13g2_a21oi_1 _18797_ (.A1(_05214_),
    .A2(_05216_),
    .Y(_05217_),
    .B1(net7120));
 sg13g2_inv_1 _18798_ (.Y(_05218_),
    .A(_05217_));
 sg13g2_xnor2_1 _18799_ (.Y(_05219_),
    .A(_05212_),
    .B(_05217_));
 sg13g2_a21oi_1 _18800_ (.A1(_05096_),
    .A2(_05105_),
    .Y(_05220_),
    .B1(_05106_));
 sg13g2_nand2_1 _18801_ (.Y(_05221_),
    .A(_05077_),
    .B(_05080_));
 sg13g2_o21ai_1 _18802_ (.B1(_05074_),
    .Y(_05222_),
    .A1(_05077_),
    .A2(_05080_));
 sg13g2_nand2_1 _18803_ (.Y(_05223_),
    .A(_05221_),
    .B(_05222_));
 sg13g2_xnor2_1 _18804_ (.Y(_05224_),
    .A(_05220_),
    .B(_05223_));
 sg13g2_xnor2_1 _18805_ (.Y(_05225_),
    .A(_05219_),
    .B(_05224_));
 sg13g2_o21ai_1 _18806_ (.B1(_05084_),
    .Y(_05226_),
    .A1(_05066_),
    .A2(_05083_));
 sg13g2_nor2_1 _18807_ (.A(net7200),
    .B(net7140),
    .Y(_05227_));
 sg13g2_nor2_1 _18808_ (.A(net7210),
    .B(net7135),
    .Y(_05228_));
 sg13g2_xnor2_1 _18809_ (.Y(_05229_),
    .A(_05227_),
    .B(_05228_));
 sg13g2_nand2_1 _18810_ (.Y(_05230_),
    .A(net7212),
    .B(_04737_));
 sg13g2_xnor2_1 _18811_ (.Y(_05231_),
    .A(_05229_),
    .B(_05230_));
 sg13g2_nor2_1 _18812_ (.A(_05052_),
    .B(_05053_),
    .Y(_05232_));
 sg13g2_a22oi_1 _18813_ (.Y(_05233_),
    .B1(_05052_),
    .B2(_05053_),
    .A2(net7064),
    .A1(net7222));
 sg13g2_or2_1 _18814_ (.X(_05234_),
    .B(_05233_),
    .A(_05232_));
 sg13g2_or2_1 _18815_ (.X(_05235_),
    .B(net7147),
    .A(_04041_));
 sg13g2_or2_1 _18816_ (.X(_05236_),
    .B(net7163),
    .A(net7183));
 sg13g2_or2_1 _18817_ (.X(_05237_),
    .B(net7152),
    .A(net7189));
 sg13g2_xnor2_1 _18818_ (.Y(_05238_),
    .A(_05235_),
    .B(_05237_));
 sg13g2_xnor2_1 _18819_ (.Y(_05239_),
    .A(_05236_),
    .B(_05238_));
 sg13g2_or2_1 _18820_ (.X(_05240_),
    .B(_05239_),
    .A(_05234_));
 sg13g2_nand2_1 _18821_ (.Y(_05241_),
    .A(_05234_),
    .B(_05239_));
 sg13g2_xor2_1 _18822_ (.B(_05239_),
    .A(_05234_),
    .X(_05242_));
 sg13g2_xnor2_1 _18823_ (.Y(_05243_),
    .A(_05231_),
    .B(_05242_));
 sg13g2_a21o_1 _18824_ (.A2(_05064_),
    .A1(_05059_),
    .B1(_05056_),
    .X(_05244_));
 sg13g2_o21ai_1 _18825_ (.B1(_05244_),
    .Y(_05245_),
    .A1(_05059_),
    .A2(_05064_));
 sg13g2_nor2_1 _18826_ (.A(net7186),
    .B(net7158),
    .Y(_05246_));
 sg13g2_nor2_1 _18827_ (.A(net7175),
    .B(net7172),
    .Y(_05247_));
 sg13g2_nor2_1 _18828_ (.A(net7180),
    .B(net7161),
    .Y(_05248_));
 sg13g2_xnor2_1 _18829_ (.Y(_05249_),
    .A(_05247_),
    .B(_05248_));
 sg13g2_xnor2_1 _18830_ (.Y(_05250_),
    .A(_05246_),
    .B(_05249_));
 sg13g2_or2_1 _18831_ (.X(_05251_),
    .B(_05062_),
    .A(_05061_));
 sg13g2_a21o_1 _18832_ (.A2(_05062_),
    .A1(_05061_),
    .B1(_05060_),
    .X(_05252_));
 sg13g2_nand2_1 _18833_ (.Y(_05253_),
    .A(_05251_),
    .B(_05252_));
 sg13g2_nand2_1 _18834_ (.Y(_05254_),
    .A(_05071_),
    .B(_05072_));
 sg13g2_o21ai_1 _18835_ (.B1(_05070_),
    .Y(_05255_),
    .A1(_05071_),
    .A2(_05072_));
 sg13g2_nand2_1 _18836_ (.Y(_05256_),
    .A(_05254_),
    .B(_05255_));
 sg13g2_xnor2_1 _18837_ (.Y(_05257_),
    .A(_05253_),
    .B(_05256_));
 sg13g2_xnor2_1 _18838_ (.Y(_05258_),
    .A(_05250_),
    .B(_05257_));
 sg13g2_or2_1 _18839_ (.X(_05259_),
    .B(_05258_),
    .A(_05245_));
 sg13g2_xor2_1 _18840_ (.B(_05258_),
    .A(_05245_),
    .X(_05260_));
 sg13g2_xnor2_1 _18841_ (.Y(_05261_),
    .A(_05243_),
    .B(_05260_));
 sg13g2_nand2_1 _18842_ (.Y(_05262_),
    .A(_05226_),
    .B(_05261_));
 sg13g2_xnor2_1 _18843_ (.Y(_05263_),
    .A(_05226_),
    .B(_05261_));
 sg13g2_xnor2_1 _18844_ (.Y(_05264_),
    .A(_05225_),
    .B(_05263_));
 sg13g2_a21oi_1 _18845_ (.A1(_05086_),
    .A2(_05119_),
    .Y(_05265_),
    .B1(_05118_));
 sg13g2_nand2_1 _18846_ (.Y(_05266_),
    .A(net6716),
    .B(_05265_));
 sg13g2_xnor2_1 _18847_ (.Y(_05267_),
    .A(_05264_),
    .B(_05265_));
 sg13g2_xnor2_1 _18848_ (.Y(_05268_),
    .A(_05202_),
    .B(_05267_));
 sg13g2_o21ai_1 _18849_ (.B1(_05121_),
    .Y(_05269_),
    .A1(_05124_),
    .A2(_05160_));
 sg13g2_nand2_1 _18850_ (.Y(_05270_),
    .A(_05152_),
    .B(_05157_));
 sg13g2_o21ai_1 _18851_ (.B1(_05270_),
    .Y(_05271_),
    .A1(_05153_),
    .A2(_05156_));
 sg13g2_a21oi_1 _18852_ (.A1(_05161_),
    .A2(_05269_),
    .Y(_05272_),
    .B1(_05271_));
 sg13g2_nand3_1 _18853_ (.B(_05269_),
    .C(_05271_),
    .A(_05161_),
    .Y(_05273_));
 sg13g2_nor2b_1 _18854_ (.A(_05272_),
    .B_N(_05273_),
    .Y(_05274_));
 sg13g2_xnor2_1 _18855_ (.Y(_05275_),
    .A(_05268_),
    .B(_05274_));
 sg13g2_nand2_1 _18856_ (.Y(_05276_),
    .A(_05220_),
    .B(_05223_));
 sg13g2_nor2_1 _18857_ (.A(_05220_),
    .B(_05223_),
    .Y(_05277_));
 sg13g2_nand2_1 _18858_ (.Y(_05278_),
    .A(_05219_),
    .B(_05276_));
 sg13g2_o21ai_1 _18859_ (.B1(_05276_),
    .Y(_05279_),
    .A1(_05219_),
    .A2(_05277_));
 sg13g2_nand2b_1 _18860_ (.Y(_05280_),
    .B(_05278_),
    .A_N(_05277_));
 sg13g2_a21oi_1 _18861_ (.A1(_01655_),
    .A2(net7325),
    .Y(_05281_),
    .B1(_05016_));
 sg13g2_a21o_1 _18862_ (.A2(net7325),
    .A1(_01655_),
    .B1(_05016_),
    .X(_05282_));
 sg13g2_nor2_1 _18863_ (.A(net7005),
    .B(net6992),
    .Y(_05283_));
 sg13g2_a21oi_1 _18864_ (.A1(_01655_),
    .A2(net7320),
    .Y(_05284_),
    .B1(net7315));
 sg13g2_a21o_1 _18865_ (.A2(net7320),
    .A1(_01655_),
    .B1(net7315),
    .X(_05285_));
 sg13g2_nand2_1 _18866_ (.Y(_05286_),
    .A(net6939),
    .B(_05188_));
 sg13g2_nor2_1 _18867_ (.A(net7002),
    .B(net6939),
    .Y(_05287_));
 sg13g2_inv_1 _18868_ (.Y(_05288_),
    .A(_00506_));
 sg13g2_inv_1 _18869_ (.Y(_05289_),
    .A(_00505_));
 sg13g2_nand2_1 _18870_ (.Y(_05290_),
    .A(_05191_),
    .B(_05197_));
 sg13g2_o21ai_1 _18871_ (.B1(_05189_),
    .Y(_05291_),
    .A1(net6939),
    .A2(_05188_));
 sg13g2_inv_1 _18872_ (.Y(_05292_),
    .A(_00504_));
 sg13g2_nand2_1 _18873_ (.Y(_05293_),
    .A(_05286_),
    .B(_05291_));
 sg13g2_xnor2_1 _18874_ (.Y(_05294_),
    .A(_05285_),
    .B(_05293_));
 sg13g2_xnor2_1 _18875_ (.Y(_05295_),
    .A(_05279_),
    .B(_05294_));
 sg13g2_inv_1 _18876_ (.Y(_05296_),
    .A(_00503_));
 sg13g2_xnor2_1 _18877_ (.Y(_05297_),
    .A(_05290_),
    .B(_05295_));
 sg13g2_o21ai_1 _18878_ (.B1(_05225_),
    .Y(_05298_),
    .A1(_05226_),
    .A2(_05261_));
 sg13g2_nand2_1 _18879_ (.Y(_05299_),
    .A(_05262_),
    .B(_05298_));
 sg13g2_nor2_1 _18880_ (.A(_05204_),
    .B(_05205_),
    .Y(_05300_));
 sg13g2_inv_1 _18881_ (.Y(_05301_),
    .A(_00502_));
 sg13g2_a21oi_1 _18882_ (.A1(_05204_),
    .A2(_05205_),
    .Y(_05302_),
    .B1(_05203_));
 sg13g2_nor2_1 _18883_ (.A(_05300_),
    .B(_05302_),
    .Y(_05303_));
 sg13g2_nor2_1 _18884_ (.A(net7203),
    .B(net7130),
    .Y(_05304_));
 sg13g2_nor2_1 _18885_ (.A(net7196),
    .B(net7136),
    .Y(_05305_));
 sg13g2_inv_1 _18886_ (.Y(_05306_),
    .A(_00501_));
 sg13g2_nor2_1 _18887_ (.A(net7207),
    .B(net7115),
    .Y(_05307_));
 sg13g2_inv_1 _18888_ (.Y(_05308_),
    .A(_00500_));
 sg13g2_xor2_1 _18889_ (.B(_05307_),
    .A(_05304_),
    .X(_05309_));
 sg13g2_xnor2_1 _18890_ (.Y(_05310_),
    .A(_05305_),
    .B(_05309_));
 sg13g2_nand2b_1 _18891_ (.Y(_05311_),
    .B(_05303_),
    .A_N(_05310_));
 sg13g2_nor2b_1 _18892_ (.A(_05303_),
    .B_N(_05310_),
    .Y(_05312_));
 sg13g2_xor2_1 _18893_ (.B(_05310_),
    .A(_05303_),
    .X(_05313_));
 sg13g2_inv_1 _18894_ (.Y(_05314_),
    .A(_00499_));
 sg13g2_xnor2_1 _18895_ (.Y(_05315_),
    .A(_05217_),
    .B(_05313_));
 sg13g2_o21ai_1 _18896_ (.B1(_05217_),
    .Y(_05316_),
    .A1(_05207_),
    .A2(_05210_));
 sg13g2_inv_1 _18897_ (.Y(_05317_),
    .A(_00498_));
 sg13g2_nand4_1 _18898_ (.B(_05252_),
    .C(_05254_),
    .A(_05251_),
    .Y(_05318_),
    .D(_05255_));
 sg13g2_a22oi_1 _18899_ (.Y(_05319_),
    .B1(_05254_),
    .B2(_05255_),
    .A2(_05252_),
    .A1(_05251_));
 sg13g2_o21ai_1 _18900_ (.B1(_05318_),
    .Y(_05320_),
    .A1(_05250_),
    .A2(_05319_));
 sg13g2_and3_1 _18901_ (.X(_05321_),
    .A(_05211_),
    .B(_05316_),
    .C(_05320_));
 sg13g2_nand3_1 _18902_ (.B(_05316_),
    .C(_05320_),
    .A(_05211_),
    .Y(_05322_));
 sg13g2_inv_1 _18903_ (.Y(_05323_),
    .A(_00497_));
 sg13g2_a21oi_1 _18904_ (.A1(_05211_),
    .A2(_05316_),
    .Y(_05324_),
    .B1(_05320_));
 sg13g2_nor2_1 _18905_ (.A(_05321_),
    .B(_05324_),
    .Y(_05325_));
 sg13g2_inv_1 _18906_ (.Y(_05326_),
    .A(_00496_));
 sg13g2_xnor2_1 _18907_ (.Y(_05327_),
    .A(_05315_),
    .B(_05325_));
 sg13g2_a21o_1 _18908_ (.A2(_05258_),
    .A1(_05245_),
    .B1(_05243_),
    .X(_05328_));
 sg13g2_nor2_1 _18909_ (.A(_04041_),
    .B(net7140),
    .Y(_05329_));
 sg13g2_nor2_1 _18910_ (.A(net7200),
    .B(net7135),
    .Y(_05330_));
 sg13g2_inv_1 _18911_ (.Y(_05331_),
    .A(_00495_));
 sg13g2_xnor2_1 _18912_ (.Y(_05332_),
    .A(_05329_),
    .B(_05330_));
 sg13g2_nand2_1 _18913_ (.Y(_05333_),
    .A(net7210),
    .B(net7064));
 sg13g2_inv_1 _18914_ (.Y(_05334_),
    .A(_00494_));
 sg13g2_xnor2_1 _18915_ (.Y(_05335_),
    .A(_05332_),
    .B(_05333_));
 sg13g2_nor2_1 _18916_ (.A(_05227_),
    .B(_05228_),
    .Y(_05336_));
 sg13g2_a22oi_1 _18917_ (.Y(_05337_),
    .B1(_05227_),
    .B2(_05228_),
    .A2(net7064),
    .A1(net7212));
 sg13g2_or2_1 _18918_ (.X(_05338_),
    .B(_05337_),
    .A(_05336_));
 sg13g2_inv_1 _18919_ (.Y(_05339_),
    .A(_00493_));
 sg13g2_nor2_1 _18920_ (.A(net7189),
    .B(net7147),
    .Y(_05340_));
 sg13g2_nor2_1 _18921_ (.A(_04215_),
    .B(net7165),
    .Y(_05341_));
 sg13g2_nor2_1 _18922_ (.A(net7183),
    .B(net7155),
    .Y(_05342_));
 sg13g2_inv_1 _18923_ (.Y(_05343_),
    .A(_00492_));
 sg13g2_xnor2_1 _18924_ (.Y(_05344_),
    .A(_05340_),
    .B(_05342_));
 sg13g2_xor2_1 _18925_ (.B(_05344_),
    .A(_05341_),
    .X(_05345_));
 sg13g2_or2_1 _18926_ (.X(_05346_),
    .B(_05345_),
    .A(_05338_));
 sg13g2_nand2_1 _18927_ (.Y(_05347_),
    .A(_05338_),
    .B(_05345_));
 sg13g2_inv_1 _18928_ (.Y(_05348_),
    .A(_00491_));
 sg13g2_xor2_1 _18929_ (.B(_05345_),
    .A(_05338_),
    .X(_05349_));
 sg13g2_inv_1 _18930_ (.Y(_05350_),
    .A(_00490_));
 sg13g2_xnor2_1 _18931_ (.Y(_05351_),
    .A(_05335_),
    .B(_05349_));
 sg13g2_a21o_1 _18932_ (.A2(_05239_),
    .A1(_05234_),
    .B1(_05231_),
    .X(_05352_));
 sg13g2_o21ai_1 _18933_ (.B1(_05231_),
    .Y(_05353_),
    .A1(_05234_),
    .A2(_05239_));
 sg13g2_inv_1 _18934_ (.Y(_05354_),
    .A(_00489_));
 sg13g2_nor2_1 _18935_ (.A(net7186),
    .B(net7151),
    .Y(_05355_));
 sg13g2_nor2_1 _18936_ (.A(net7180),
    .B(net7158),
    .Y(_05356_));
 sg13g2_nor2_1 _18937_ (.A(net7172),
    .B(net7161),
    .Y(_05357_));
 sg13g2_inv_1 _18938_ (.Y(_05358_),
    .A(_00488_));
 sg13g2_xnor2_1 _18939_ (.Y(_05359_),
    .A(net7052),
    .B(_05357_));
 sg13g2_xor2_1 _18940_ (.B(_05359_),
    .A(_05356_),
    .X(_05360_));
 sg13g2_xnor2_1 _18941_ (.Y(_05361_),
    .A(_05356_),
    .B(_05359_));
 sg13g2_or2_1 _18942_ (.X(_05362_),
    .B(_05237_),
    .A(_05236_));
 sg13g2_nand2_1 _18943_ (.Y(_05363_),
    .A(_05236_),
    .B(_05237_));
 sg13g2_inv_1 _18944_ (.Y(_05364_),
    .A(_00487_));
 sg13g2_a21o_1 _18945_ (.A2(_05237_),
    .A1(_05236_),
    .B1(_05235_),
    .X(_05365_));
 sg13g2_o21ai_1 _18946_ (.B1(_05235_),
    .Y(_05366_),
    .A1(_05236_),
    .A2(_05237_));
 sg13g2_nand2_1 _18947_ (.Y(_05367_),
    .A(_05362_),
    .B(_05365_));
 sg13g2_o21ai_1 _18948_ (.B1(_05246_),
    .Y(_05368_),
    .A1(_05247_),
    .A2(_05248_));
 sg13g2_nand2_1 _18949_ (.Y(_05369_),
    .A(_05247_),
    .B(_05248_));
 sg13g2_a21o_1 _18950_ (.A2(_05247_),
    .A1(_05246_),
    .B1(_05248_),
    .X(_05370_));
 sg13g2_inv_1 _18951_ (.Y(_05371_),
    .A(_00486_));
 sg13g2_or2_1 _18952_ (.X(_05372_),
    .B(_05247_),
    .A(_05246_));
 sg13g2_nand2_1 _18953_ (.Y(_05373_),
    .A(_05368_),
    .B(_05369_));
 sg13g2_a22oi_1 _18954_ (.Y(_05374_),
    .B1(_05370_),
    .B2(_05372_),
    .A2(_05365_),
    .A1(_05362_));
 sg13g2_nand4_1 _18955_ (.B(_05366_),
    .C(_05368_),
    .A(_05363_),
    .Y(_05375_),
    .D(_05369_));
 sg13g2_a22oi_1 _18956_ (.Y(_05376_),
    .B1(_05368_),
    .B2(_05369_),
    .A2(_05366_),
    .A1(_05363_));
 sg13g2_nand4_1 _18957_ (.B(_05365_),
    .C(_05370_),
    .A(_05362_),
    .Y(_05377_),
    .D(_05372_));
 sg13g2_nand3_1 _18958_ (.B(_05375_),
    .C(_05377_),
    .A(_05360_),
    .Y(_05378_));
 sg13g2_o21ai_1 _18959_ (.B1(_05361_),
    .Y(_05379_),
    .A1(_05374_),
    .A2(_05376_));
 sg13g2_nand3_1 _18960_ (.B(_05375_),
    .C(_05377_),
    .A(_05361_),
    .Y(_05380_));
 sg13g2_o21ai_1 _18961_ (.B1(_05360_),
    .Y(_05381_),
    .A1(_05374_),
    .A2(_05376_));
 sg13g2_inv_1 _18962_ (.Y(_05382_),
    .A(_00485_));
 sg13g2_a22oi_1 _18963_ (.Y(_05383_),
    .B1(_05380_),
    .B2(_05381_),
    .A2(_05352_),
    .A1(_05240_));
 sg13g2_nand4_1 _18964_ (.B(_05353_),
    .C(_05378_),
    .A(_05241_),
    .Y(_05384_),
    .D(_05379_));
 sg13g2_nand4_1 _18965_ (.B(_05352_),
    .C(_05380_),
    .A(_05240_),
    .Y(_05385_),
    .D(_05381_));
 sg13g2_a21o_1 _18966_ (.A2(_05385_),
    .A1(_05384_),
    .B1(_05351_),
    .X(_05386_));
 sg13g2_nand3_1 _18967_ (.B(_05384_),
    .C(_05385_),
    .A(_05351_),
    .Y(_05387_));
 sg13g2_inv_1 _18968_ (.Y(_05388_),
    .A(_00484_));
 sg13g2_and4_1 _18969_ (.A(_05259_),
    .B(_05328_),
    .C(_05386_),
    .D(_05387_),
    .X(_05389_));
 sg13g2_nand4_1 _18970_ (.B(_05328_),
    .C(_05386_),
    .A(_05259_),
    .Y(_05390_),
    .D(_05387_));
 sg13g2_a22oi_1 _18971_ (.Y(_05391_),
    .B1(_05386_),
    .B2(_05387_),
    .A2(_05328_),
    .A1(_05259_));
 sg13g2_nor2_1 _18972_ (.A(_05389_),
    .B(_05391_),
    .Y(_05392_));
 sg13g2_xor2_1 _18973_ (.B(_05392_),
    .A(_05327_),
    .X(_05393_));
 sg13g2_nand2_1 _18974_ (.Y(_05394_),
    .A(_05299_),
    .B(_05393_));
 sg13g2_xnor2_1 _18975_ (.Y(_05395_),
    .A(_05299_),
    .B(_05393_));
 sg13g2_xnor2_1 _18976_ (.Y(_05396_),
    .A(_05297_),
    .B(_05395_));
 sg13g2_a21oi_1 _18977_ (.A1(net6716),
    .A2(_05265_),
    .Y(_05397_),
    .B1(_05202_));
 sg13g2_nor2_1 _18978_ (.A(_05126_),
    .B(_05147_),
    .Y(_05398_));
 sg13g2_o21ai_1 _18979_ (.B1(_05133_),
    .Y(_05399_),
    .A1(_05173_),
    .A2(_05398_));
 sg13g2_nand2_1 _18980_ (.Y(_05400_),
    .A(_05126_),
    .B(_05147_));
 sg13g2_nand2_1 _18981_ (.Y(_05401_),
    .A(_05136_),
    .B(_05400_));
 sg13g2_o21ai_1 _18982_ (.B1(_05147_),
    .Y(_05402_),
    .A1(_05126_),
    .A2(_05137_));
 sg13g2_nand2_1 _18983_ (.Y(_05403_),
    .A(_05173_),
    .B(_05402_));
 sg13g2_nand4_1 _18984_ (.B(_05399_),
    .C(_05401_),
    .A(_05181_),
    .Y(_05404_),
    .D(_05403_));
 sg13g2_o21ai_1 _18985_ (.B1(_05132_),
    .Y(_05405_),
    .A1(_05173_),
    .A2(_05400_));
 sg13g2_a21oi_1 _18986_ (.A1(_05126_),
    .A2(_05137_),
    .Y(_05406_),
    .B1(_05181_));
 sg13g2_nand3_1 _18987_ (.B(_05405_),
    .C(_05406_),
    .A(_05403_),
    .Y(_05407_));
 sg13g2_and2_1 _18988_ (.A(_05404_),
    .B(_05407_),
    .X(_05408_));
 sg13g2_o21ai_1 _18989_ (.B1(_05408_),
    .Y(_05409_),
    .A1(net6716),
    .A2(_05265_));
 sg13g2_nor2_1 _18990_ (.A(_05397_),
    .B(_05409_),
    .Y(_05410_));
 sg13g2_or2_1 _18991_ (.X(_05411_),
    .B(_05409_),
    .A(_05397_));
 sg13g2_nor3_1 _18992_ (.A(net6716),
    .B(_05265_),
    .C(_05408_),
    .Y(_05412_));
 sg13g2_nor2_1 _18993_ (.A(_05202_),
    .B(_05408_),
    .Y(_05413_));
 sg13g2_a21oi_1 _18994_ (.A1(_05266_),
    .A2(_05413_),
    .Y(_05414_),
    .B1(_05412_));
 sg13g2_nand3_1 _18995_ (.B(_05411_),
    .C(_05414_),
    .A(_05396_),
    .Y(_05415_));
 sg13g2_a21o_1 _18996_ (.A2(_05414_),
    .A1(_05411_),
    .B1(_05396_),
    .X(_05416_));
 sg13g2_nand2_1 _18997_ (.Y(_05417_),
    .A(_05415_),
    .B(_05416_));
 sg13g2_nor2_1 _18998_ (.A(_05026_),
    .B(_05185_),
    .Y(_05418_));
 sg13g2_inv_1 _18999_ (.Y(_05419_),
    .A(_00003_));
 sg13g2_a21oi_1 _19000_ (.A1(_05315_),
    .A2(_05322_),
    .Y(_05420_),
    .B1(_05324_));
 sg13g2_nand3b_1 _19001_ (.B(_05176_),
    .C(_05281_),
    .Y(_05421_),
    .A_N(_05130_));
 sg13g2_o21ai_1 _19002_ (.B1(_05421_),
    .Y(_05422_),
    .A1(_05176_),
    .A2(_05281_));
 sg13g2_nor2b_1 _19003_ (.A(net7060),
    .B_N(_05177_),
    .Y(_05423_));
 sg13g2_nor2_1 _19004_ (.A(_05177_),
    .B(_05282_),
    .Y(_05424_));
 sg13g2_nor4_1 _19005_ (.A(_05130_),
    .B(_05176_),
    .C(_05177_),
    .D(_05282_),
    .Y(_05425_));
 sg13g2_a21oi_1 _19006_ (.A1(_05422_),
    .A2(_05423_),
    .Y(_05426_),
    .B1(_05425_));
 sg13g2_nor2_1 _19007_ (.A(_05025_),
    .B(net6992),
    .Y(_05427_));
 sg13g2_nand2_1 _19008_ (.Y(_05428_),
    .A(net6992),
    .B(_05424_));
 sg13g2_o21ai_1 _19009_ (.B1(_05428_),
    .Y(_05429_),
    .A1(_05176_),
    .A2(_05281_));
 sg13g2_a221oi_1 _19010_ (.B2(net7059),
    .C1(net7005),
    .B1(_05429_),
    .A1(_05424_),
    .Y(_05430_),
    .A2(_05427_));
 sg13g2_a21oi_1 _19011_ (.A1(net7005),
    .A2(_05426_),
    .Y(_05431_),
    .B1(_05430_));
 sg13g2_nand2b_1 _19012_ (.Y(_05432_),
    .B(_05420_),
    .A_N(_05431_));
 sg13g2_nor2b_1 _19013_ (.A(_05420_),
    .B_N(_05431_),
    .Y(_05433_));
 sg13g2_xnor2_1 _19014_ (.Y(_05434_),
    .A(_05420_),
    .B(_05431_));
 sg13g2_a21oi_1 _19015_ (.A1(_01656_),
    .A2(net7325),
    .Y(_05435_),
    .B1(_05016_));
 sg13g2_a21oi_1 _19016_ (.A1(net6992),
    .A2(_05281_),
    .Y(_05436_),
    .B1(_05283_));
 sg13g2_nand2_1 _19017_ (.Y(_05437_),
    .A(net7005),
    .B(_05177_));
 sg13g2_a21oi_1 _19018_ (.A1(_05176_),
    .A2(_05282_),
    .Y(_05438_),
    .B1(_05437_));
 sg13g2_nor2_1 _19019_ (.A(_05176_),
    .B(_05282_),
    .Y(_05439_));
 sg13g2_nor3_1 _19020_ (.A(net7059),
    .B(_05438_),
    .C(_05439_),
    .Y(_05440_));
 sg13g2_a21oi_1 _19021_ (.A1(net7060),
    .A2(_05436_),
    .Y(_05441_),
    .B1(_05440_));
 sg13g2_xnor2_1 _19022_ (.Y(_05442_),
    .A(_05435_),
    .B(_05441_));
 sg13g2_nand2_1 _19023_ (.Y(_05443_),
    .A(_01656_),
    .B(net7320));
 sg13g2_a21oi_1 _19024_ (.A1(_01656_),
    .A2(net7320),
    .Y(_05444_),
    .B1(net7314));
 sg13g2_nand2_1 _19025_ (.Y(_05445_),
    .A(_05019_),
    .B(_05443_));
 sg13g2_xnor2_1 _19026_ (.Y(_05446_),
    .A(_05434_),
    .B(_05442_));
 sg13g2_a21oi_1 _19027_ (.A1(_04576_),
    .A2(_04678_),
    .Y(_05447_),
    .B1(net7197));
 sg13g2_nor4_1 _19028_ (.A(_03970_),
    .B(_04019_),
    .C(_04020_),
    .D(_04677_),
    .Y(_05448_));
 sg13g2_nor4_1 _19029_ (.A(net7205),
    .B(_04794_),
    .C(_05447_),
    .D(_05448_),
    .Y(_05449_));
 sg13g2_nor2_1 _19030_ (.A(net7197),
    .B(_04678_),
    .Y(_05450_));
 sg13g2_nor2b_1 _19031_ (.A(net7205),
    .B_N(_04576_),
    .Y(_05451_));
 sg13g2_nand2_1 _19032_ (.Y(_05452_),
    .A(_04576_),
    .B(_04798_));
 sg13g2_o21ai_1 _19033_ (.B1(_05452_),
    .Y(_05453_),
    .A1(_03971_),
    .A2(_05451_));
 sg13g2_o21ai_1 _19034_ (.B1(_04022_),
    .Y(_05454_),
    .A1(_04576_),
    .A2(_04678_));
 sg13g2_and3_1 _19035_ (.X(_05455_),
    .A(net7205),
    .B(_03971_),
    .C(net7061));
 sg13g2_a221oi_1 _19036_ (.B2(_05455_),
    .C1(_05449_),
    .B1(_05454_),
    .A1(_05450_),
    .Y(_05456_),
    .A2(_05453_));
 sg13g2_nor2b_1 _19037_ (.A(_05456_),
    .B_N(_05217_),
    .Y(_05457_));
 sg13g2_xnor2_1 _19038_ (.Y(_05458_),
    .A(_05217_),
    .B(_05456_));
 sg13g2_nand2_1 _19039_ (.Y(_05459_),
    .A(_05367_),
    .B(_05373_));
 sg13g2_o21ai_1 _19040_ (.B1(_05361_),
    .Y(_05460_),
    .A1(_05367_),
    .A2(_05373_));
 sg13g2_nand2_1 _19041_ (.Y(_05461_),
    .A(_05459_),
    .B(_05460_));
 sg13g2_a21oi_1 _19042_ (.A1(_05218_),
    .A2(_05311_),
    .Y(_05462_),
    .B1(_05312_));
 sg13g2_xnor2_1 _19043_ (.Y(_05463_),
    .A(_05461_),
    .B(_05462_));
 sg13g2_inv_1 _19044_ (.Y(_05464_),
    .A(_00462_));
 sg13g2_xnor2_1 _19045_ (.Y(_05465_),
    .A(_05458_),
    .B(_05463_));
 sg13g2_nor2_1 _19046_ (.A(net7189),
    .B(net7141),
    .Y(_05466_));
 sg13g2_nor2_1 _19047_ (.A(_04041_),
    .B(_04649_),
    .Y(_05467_));
 sg13g2_xnor2_1 _19048_ (.Y(_05468_),
    .A(_05466_),
    .B(_05467_));
 sg13g2_nand2_1 _19049_ (.Y(_05469_),
    .A(net7200),
    .B(net7064));
 sg13g2_xnor2_1 _19050_ (.Y(_05470_),
    .A(_05468_),
    .B(_05469_));
 sg13g2_nor2_1 _19051_ (.A(_05329_),
    .B(_05330_),
    .Y(_05471_));
 sg13g2_a22oi_1 _19052_ (.Y(_05472_),
    .B1(_05329_),
    .B2(_05330_),
    .A2(net7064),
    .A1(net7210));
 sg13g2_nor2_1 _19053_ (.A(_05471_),
    .B(_05472_),
    .Y(_05473_));
 sg13g2_nor2_1 _19054_ (.A(net7182),
    .B(net7146),
    .Y(_05474_));
 sg13g2_nor2_1 _19055_ (.A(net7165),
    .B(net7160),
    .Y(_05475_));
 sg13g2_nor2_1 _19056_ (.A(net7176),
    .B(net7154),
    .Y(_05476_));
 sg13g2_xor2_1 _19057_ (.B(_05476_),
    .A(_05475_),
    .X(_05477_));
 sg13g2_xnor2_1 _19058_ (.Y(_05478_),
    .A(_05474_),
    .B(_05477_));
 sg13g2_nand2b_1 _19059_ (.Y(_05479_),
    .B(_05473_),
    .A_N(_05478_));
 sg13g2_nor2b_1 _19060_ (.A(_05473_),
    .B_N(_05478_),
    .Y(_05480_));
 sg13g2_xnor2_1 _19061_ (.Y(_05481_),
    .A(_05473_),
    .B(_05478_));
 sg13g2_xnor2_1 _19062_ (.Y(_05482_),
    .A(_05470_),
    .B(_05481_));
 sg13g2_a21o_1 _19063_ (.A2(_05345_),
    .A1(_05338_),
    .B1(_05335_),
    .X(_05483_));
 sg13g2_o21ai_1 _19064_ (.B1(_05335_),
    .Y(_05484_),
    .A1(_05338_),
    .A2(_05345_));
 sg13g2_nor2_1 _19065_ (.A(net7186),
    .B(net7138),
    .Y(_05485_));
 sg13g2_nor2_1 _19066_ (.A(net7171),
    .B(net7158),
    .Y(_05486_));
 sg13g2_nor2_1 _19067_ (.A(net7180),
    .B(net7151),
    .Y(_05487_));
 sg13g2_xnor2_1 _19068_ (.Y(_05488_),
    .A(_05485_),
    .B(_05487_));
 sg13g2_xor2_1 _19069_ (.B(_05488_),
    .A(_05486_),
    .X(_05489_));
 sg13g2_xnor2_1 _19070_ (.Y(_05490_),
    .A(_05486_),
    .B(net6990));
 sg13g2_nand2_1 _19071_ (.Y(_05491_),
    .A(_05341_),
    .B(_05342_));
 sg13g2_or2_1 _19072_ (.X(_05492_),
    .B(_05342_),
    .A(_05341_));
 sg13g2_o21ai_1 _19073_ (.B1(_05340_),
    .Y(_05493_),
    .A1(_05341_),
    .A2(_05342_));
 sg13g2_a21o_1 _19074_ (.A2(_05342_),
    .A1(_05341_),
    .B1(_05340_),
    .X(_05494_));
 sg13g2_or2_1 _19075_ (.X(_05495_),
    .B(_05357_),
    .A(_05356_));
 sg13g2_a21o_1 _19076_ (.A2(_05357_),
    .A1(_05356_),
    .B1(_05355_),
    .X(_05496_));
 sg13g2_a22oi_1 _19077_ (.Y(_05497_),
    .B1(_05495_),
    .B2(_05496_),
    .A2(_05493_),
    .A1(_05491_));
 sg13g2_and4_1 _19078_ (.A(_05491_),
    .B(_05493_),
    .C(_05495_),
    .D(_05496_),
    .X(_05498_));
 sg13g2_or3_1 _19079_ (.A(_05490_),
    .B(_05497_),
    .C(_05498_),
    .X(_05499_));
 sg13g2_o21ai_1 _19080_ (.B1(_05490_),
    .Y(_05500_),
    .A1(_05497_),
    .A2(net6934));
 sg13g2_or3_1 _19081_ (.A(_05489_),
    .B(_05497_),
    .C(_05498_),
    .X(_05501_));
 sg13g2_o21ai_1 _19082_ (.B1(_05489_),
    .Y(_05502_),
    .A1(_05497_),
    .A2(net6934));
 sg13g2_a22oi_1 _19083_ (.Y(_05503_),
    .B1(_05501_),
    .B2(_05502_),
    .A2(_05483_),
    .A1(_05346_));
 sg13g2_nand4_1 _19084_ (.B(_05484_),
    .C(_05499_),
    .A(_05347_),
    .Y(_05504_),
    .D(_05500_));
 sg13g2_nand4_1 _19085_ (.B(_05483_),
    .C(_05501_),
    .A(_05346_),
    .Y(_05505_),
    .D(_05502_));
 sg13g2_a21oi_1 _19086_ (.A1(_05504_),
    .A2(_05505_),
    .Y(_05506_),
    .B1(_05482_));
 sg13g2_and3_1 _19087_ (.X(_05507_),
    .A(_05482_),
    .B(_05504_),
    .C(_05505_));
 sg13g2_o21ai_1 _19088_ (.B1(_05385_),
    .Y(_05508_),
    .A1(_05351_),
    .A2(_05383_));
 sg13g2_o21ai_1 _19089_ (.B1(_05508_),
    .Y(_05509_),
    .A1(_05506_),
    .A2(_05507_));
 sg13g2_nor3_1 _19090_ (.A(_05506_),
    .B(net6830),
    .C(_05508_),
    .Y(_05510_));
 sg13g2_or3_1 _19091_ (.A(_05506_),
    .B(_05507_),
    .C(_05508_),
    .X(_05511_));
 sg13g2_nand2_1 _19092_ (.Y(_05512_),
    .A(net6782),
    .B(_05511_));
 sg13g2_xnor2_1 _19093_ (.Y(_05513_),
    .A(_05465_),
    .B(_05512_));
 sg13g2_o21ai_1 _19094_ (.B1(_05390_),
    .Y(_05514_),
    .A1(_05327_),
    .A2(_05391_));
 sg13g2_nand2_1 _19095_ (.Y(_05515_),
    .A(net6715),
    .B(_05514_));
 sg13g2_nor2_1 _19096_ (.A(net6715),
    .B(_05514_),
    .Y(_05516_));
 sg13g2_xnor2_1 _19097_ (.Y(_05517_),
    .A(_05446_),
    .B(_05514_));
 sg13g2_xor2_1 _19098_ (.B(_05517_),
    .A(net6715),
    .X(_05518_));
 sg13g2_xnor2_1 _19099_ (.Y(_05519_),
    .A(net6715),
    .B(_05517_));
 sg13g2_nand2_1 _19100_ (.Y(_05520_),
    .A(_05280_),
    .B(_05290_));
 sg13g2_o21ai_1 _19101_ (.B1(_05297_),
    .Y(_05521_),
    .A1(_05299_),
    .A2(_05393_));
 sg13g2_nand2_1 _19102_ (.Y(_05522_),
    .A(_05394_),
    .B(_05521_));
 sg13g2_nor2_1 _19103_ (.A(_05280_),
    .B(_05290_),
    .Y(_05523_));
 sg13g2_a21oi_1 _19104_ (.A1(_05294_),
    .A2(_05520_),
    .Y(_05524_),
    .B1(_05523_));
 sg13g2_a21o_1 _19105_ (.A2(_05520_),
    .A1(_05294_),
    .B1(_05523_),
    .X(_05525_));
 sg13g2_xnor2_1 _19106_ (.Y(_05526_),
    .A(_05518_),
    .B(_05524_));
 sg13g2_xnor2_1 _19107_ (.Y(_05527_),
    .A(_05522_),
    .B(_05526_));
 sg13g2_a21o_1 _19108_ (.A2(_05515_),
    .A1(_05446_),
    .B1(_05516_),
    .X(_05528_));
 sg13g2_nor2_1 _19109_ (.A(net7182),
    .B(net7142),
    .Y(_05529_));
 sg13g2_nor2_1 _19110_ (.A(net7189),
    .B(_04649_),
    .Y(_05530_));
 sg13g2_xnor2_1 _19111_ (.Y(_05531_),
    .A(_05529_),
    .B(_05530_));
 sg13g2_nand2_1 _19112_ (.Y(_05532_),
    .A(_04041_),
    .B(_04737_));
 sg13g2_xnor2_1 _19113_ (.Y(_05533_),
    .A(_05531_),
    .B(_05532_));
 sg13g2_nor2_1 _19114_ (.A(_05466_),
    .B(_05467_),
    .Y(_05534_));
 sg13g2_a22oi_1 _19115_ (.Y(_05535_),
    .B1(_05466_),
    .B2(_05467_),
    .A2(net7064),
    .A1(net7200));
 sg13g2_or2_1 _19116_ (.X(_05536_),
    .B(_05535_),
    .A(_05534_));
 sg13g2_nor2_1 _19117_ (.A(net7160),
    .B(net7155),
    .Y(_05537_));
 sg13g2_nor2_1 _19118_ (.A(net7166),
    .B(net7157),
    .Y(_05538_));
 sg13g2_nor2_1 _19119_ (.A(net7176),
    .B(net7146),
    .Y(_05539_));
 sg13g2_xor2_1 _19120_ (.B(_05539_),
    .A(_05537_),
    .X(_05540_));
 sg13g2_xnor2_1 _19121_ (.Y(_05541_),
    .A(_05538_),
    .B(_05540_));
 sg13g2_or2_1 _19122_ (.X(_05542_),
    .B(_05541_),
    .A(_05536_));
 sg13g2_nand2_1 _19123_ (.Y(_05543_),
    .A(_05536_),
    .B(_05541_));
 sg13g2_nand2_1 _19124_ (.Y(_05544_),
    .A(_05542_),
    .B(_05543_));
 sg13g2_xnor2_1 _19125_ (.Y(_05545_),
    .A(_05533_),
    .B(_05544_));
 sg13g2_o21ai_1 _19126_ (.B1(_05479_),
    .Y(_05546_),
    .A1(_05470_),
    .A2(_05480_));
 sg13g2_nand2b_1 _19127_ (.Y(_05547_),
    .B(net7133),
    .A_N(net7185));
 sg13g2_or2_1 _19128_ (.X(_05548_),
    .B(net7151),
    .A(net7171));
 sg13g2_or2_1 _19129_ (.X(_05549_),
    .B(net7138),
    .A(net7179));
 sg13g2_xor2_1 _19130_ (.B(_05549_),
    .A(_05548_),
    .X(_05550_));
 sg13g2_xnor2_1 _19131_ (.Y(_05551_),
    .A(_05547_),
    .B(_05550_));
 sg13g2_inv_1 _19132_ (.Y(_05552_),
    .A(_00434_));
 sg13g2_nor2_1 _19133_ (.A(_05475_),
    .B(_05476_),
    .Y(_05553_));
 sg13g2_a21oi_1 _19134_ (.A1(_05475_),
    .A2(_05476_),
    .Y(_05554_),
    .B1(_05474_));
 sg13g2_nor2_1 _19135_ (.A(_05553_),
    .B(_05554_),
    .Y(_05555_));
 sg13g2_nor2_1 _19136_ (.A(_05486_),
    .B(_05487_),
    .Y(_05556_));
 sg13g2_a21oi_1 _19137_ (.A1(_05486_),
    .A2(_05487_),
    .Y(_05557_),
    .B1(_05485_));
 sg13g2_nor2_1 _19138_ (.A(_05556_),
    .B(_05557_),
    .Y(_05558_));
 sg13g2_xor2_1 _19139_ (.B(_05558_),
    .A(_05555_),
    .X(_05559_));
 sg13g2_xnor2_1 _19140_ (.Y(_05560_),
    .A(_05551_),
    .B(_05559_));
 sg13g2_nand2b_1 _19141_ (.Y(_05561_),
    .B(_05546_),
    .A_N(_05560_));
 sg13g2_nor2b_1 _19142_ (.A(_05546_),
    .B_N(_05560_),
    .Y(_05562_));
 sg13g2_xnor2_1 _19143_ (.Y(_05563_),
    .A(_05546_),
    .B(_05560_));
 sg13g2_xnor2_1 _19144_ (.Y(_05564_),
    .A(_05545_),
    .B(_05563_));
 sg13g2_nand3_1 _19145_ (.B(net7115),
    .C(_05205_),
    .A(net7133),
    .Y(_05565_));
 sg13g2_nor2_1 _19146_ (.A(net7136),
    .B(net7133),
    .Y(_05566_));
 sg13g2_o21ai_1 _19147_ (.B1(_05307_),
    .Y(_05567_),
    .A1(_05304_),
    .A2(_05566_));
 sg13g2_a21oi_1 _19148_ (.A1(_05565_),
    .A2(_05567_),
    .Y(_05568_),
    .B1(net7196));
 sg13g2_nor2_1 _19149_ (.A(_05457_),
    .B(_05568_),
    .Y(_05569_));
 sg13g2_a22oi_1 _19150_ (.Y(_05570_),
    .B1(_05495_),
    .B2(_05496_),
    .A2(_05494_),
    .A1(_05492_));
 sg13g2_nand4_1 _19151_ (.B(_05494_),
    .C(_05495_),
    .A(_05492_),
    .Y(_05571_),
    .D(_05496_));
 sg13g2_a21oi_1 _19152_ (.A1(_05489_),
    .A2(_05571_),
    .Y(_05572_),
    .B1(_05570_));
 sg13g2_nor3_1 _19153_ (.A(net7208),
    .B(_03970_),
    .C(_04021_),
    .Y(_05573_));
 sg13g2_and3_1 _19154_ (.X(_05574_),
    .A(net7207),
    .B(net7203),
    .C(net7196));
 sg13g2_or2_1 _19155_ (.X(_05575_),
    .B(_05574_),
    .A(_05573_));
 sg13g2_a21oi_1 _19156_ (.A1(_05214_),
    .A2(_05216_),
    .Y(_05576_),
    .B1(_05575_));
 sg13g2_and3_1 _19157_ (.X(_05577_),
    .A(_05214_),
    .B(_05216_),
    .C(_05575_));
 sg13g2_nor3_1 _19158_ (.A(net7116),
    .B(_05576_),
    .C(_05577_),
    .Y(_05578_));
 sg13g2_or3_1 _19159_ (.A(net7114),
    .B(_05576_),
    .C(_05577_),
    .X(_05579_));
 sg13g2_nor2_1 _19160_ (.A(net6896),
    .B(net6895),
    .Y(_05580_));
 sg13g2_nand2_1 _19161_ (.Y(_05581_),
    .A(net6896),
    .B(net6895));
 sg13g2_xnor2_1 _19162_ (.Y(_05582_),
    .A(_05572_),
    .B(_05578_));
 sg13g2_xnor2_1 _19163_ (.Y(_05583_),
    .A(_05569_),
    .B(_05582_));
 sg13g2_nand2_1 _19164_ (.Y(_05584_),
    .A(_05482_),
    .B(net6861));
 sg13g2_o21ai_1 _19165_ (.B1(_05505_),
    .Y(_05585_),
    .A1(_05482_),
    .A2(_05503_));
 sg13g2_nand2_1 _19166_ (.Y(_05586_),
    .A(_05504_),
    .B(_05584_));
 sg13g2_nand2_1 _19167_ (.Y(_05587_),
    .A(_05564_),
    .B(_05586_));
 sg13g2_nor2_1 _19168_ (.A(_05564_),
    .B(_05586_),
    .Y(_05588_));
 sg13g2_xor2_1 _19169_ (.B(_05585_),
    .A(_05583_),
    .X(_05589_));
 sg13g2_xnor2_1 _19170_ (.Y(_05590_),
    .A(_05564_),
    .B(_05589_));
 sg13g2_a21oi_1 _19171_ (.A1(_05465_),
    .A2(_05509_),
    .Y(_05591_),
    .B1(_05510_));
 sg13g2_xnor2_1 _19172_ (.Y(_05592_),
    .A(_05590_),
    .B(net6740));
 sg13g2_xor2_1 _19173_ (.B(_05591_),
    .A(_05590_),
    .X(_05593_));
 sg13g2_a21o_1 _19174_ (.A2(_05462_),
    .A1(_05461_),
    .B1(_05458_),
    .X(_05594_));
 sg13g2_o21ai_1 _19175_ (.B1(_05594_),
    .Y(_05595_),
    .A1(_05461_),
    .A2(_05462_));
 sg13g2_nand2_1 _19176_ (.Y(_05596_),
    .A(_05184_),
    .B(_05445_));
 sg13g2_nor2_1 _19177_ (.A(_05284_),
    .B(_05445_),
    .Y(_05597_));
 sg13g2_nand2_1 _19178_ (.Y(_05598_),
    .A(_05285_),
    .B(_05444_));
 sg13g2_o21ai_1 _19179_ (.B1(_05596_),
    .Y(_05599_),
    .A1(_05184_),
    .A2(_05598_));
 sg13g2_a22oi_1 _19180_ (.Y(_05600_),
    .B1(_05599_),
    .B2(_05026_),
    .A2(_05597_),
    .A1(_05418_));
 sg13g2_o21ai_1 _19181_ (.B1(_05596_),
    .Y(_05601_),
    .A1(_05286_),
    .A2(_05445_));
 sg13g2_nor2_1 _19182_ (.A(_05026_),
    .B(_05285_),
    .Y(_05602_));
 sg13g2_nor2_1 _19183_ (.A(_05187_),
    .B(_05598_),
    .Y(_05603_));
 sg13g2_a22oi_1 _19184_ (.Y(_05604_),
    .B1(_05603_),
    .B2(_05184_),
    .A2(_05602_),
    .A1(_05601_));
 sg13g2_mux2_1 _19185_ (.A0(_05600_),
    .A1(_05604_),
    .S(net7004),
    .X(_05605_));
 sg13g2_xor2_1 _19186_ (.B(_05605_),
    .A(_05595_),
    .X(_05606_));
 sg13g2_a21oi_1 _19187_ (.A1(_01657_),
    .A2(net7325),
    .Y(_05607_),
    .B1(_05016_));
 sg13g2_inv_1 _19188_ (.Y(_05608_),
    .A(_05607_));
 sg13g2_a21oi_1 _19189_ (.A1(_01657_),
    .A2(net7323),
    .Y(_05609_),
    .B1(net7314));
 sg13g2_a21o_1 _19190_ (.A2(net7323),
    .A1(_01657_),
    .B1(net7314),
    .X(_05610_));
 sg13g2_nor2_1 _19191_ (.A(net6943),
    .B(_05444_),
    .Y(_05611_));
 sg13g2_nand2_1 _19192_ (.Y(_05612_),
    .A(net7002),
    .B(_05284_));
 sg13g2_nand2_1 _19193_ (.Y(_05613_),
    .A(net6943),
    .B(_05444_));
 sg13g2_o21ai_1 _19194_ (.B1(_05613_),
    .Y(_05614_),
    .A1(_05611_),
    .A2(_05612_));
 sg13g2_nor2_1 _19195_ (.A(net7058),
    .B(_05614_),
    .Y(_05615_));
 sg13g2_a21oi_1 _19196_ (.A1(net6936),
    .A2(_05444_),
    .Y(_05616_),
    .B1(_05287_));
 sg13g2_a21oi_1 _19197_ (.A1(net7058),
    .A2(_05616_),
    .Y(_05617_),
    .B1(_05615_));
 sg13g2_xnor2_1 _19198_ (.Y(_05618_),
    .A(_05609_),
    .B(_05617_));
 sg13g2_mux2_1 _19199_ (.A0(_05600_),
    .A1(_05604_),
    .S(net7004),
    .X(_05619_));
 sg13g2_nor2_1 _19200_ (.A(net6993),
    .B(_05616_),
    .Y(_05620_));
 sg13g2_a21oi_1 _19201_ (.A1(net6993),
    .A2(_05614_),
    .Y(_05621_),
    .B1(_05620_));
 sg13g2_xnor2_1 _19202_ (.Y(_05622_),
    .A(_05610_),
    .B(_05621_));
 sg13g2_xnor2_1 _19203_ (.Y(_05623_),
    .A(_05606_),
    .B(_05618_));
 sg13g2_a21oi_1 _19204_ (.A1(_05432_),
    .A2(_05442_),
    .Y(_05624_),
    .B1(_05433_));
 sg13g2_nand3_1 _19205_ (.B(_05623_),
    .C(_05624_),
    .A(_05593_),
    .Y(_05625_));
 sg13g2_nand3b_1 _19206_ (.B(_05624_),
    .C(_05592_),
    .Y(_05626_),
    .A_N(_05623_));
 sg13g2_xnor2_1 _19207_ (.Y(_05627_),
    .A(_05593_),
    .B(_05623_));
 sg13g2_or3_1 _19208_ (.A(_05592_),
    .B(_05623_),
    .C(_05624_),
    .X(_05628_));
 sg13g2_nand3b_1 _19209_ (.B(_05623_),
    .C(_05592_),
    .Y(_05629_),
    .A_N(_05624_));
 sg13g2_nand4_1 _19210_ (.B(_05626_),
    .C(_05628_),
    .A(_05625_),
    .Y(_05630_),
    .D(_05629_));
 sg13g2_xnor2_1 _19211_ (.Y(_05631_),
    .A(_05528_),
    .B(_05630_));
 sg13g2_a21oi_1 _19212_ (.A1(_05569_),
    .A2(_05581_),
    .Y(_05632_),
    .B1(_05580_));
 sg13g2_a21o_1 _19213_ (.A2(_05608_),
    .A1(_05435_),
    .B1(net7060),
    .X(_05633_));
 sg13g2_a22oi_1 _19214_ (.Y(_05634_),
    .B1(_05633_),
    .B2(net7005),
    .A2(_05608_),
    .A1(net7060));
 sg13g2_xor2_1 _19215_ (.B(net6992),
    .A(net7060),
    .X(_05635_));
 sg13g2_nor3_1 _19216_ (.A(net7005),
    .B(_05435_),
    .C(_05635_),
    .Y(_05636_));
 sg13g2_xor2_1 _19217_ (.B(_05435_),
    .A(net6992),
    .X(_05637_));
 sg13g2_nor3_1 _19218_ (.A(_04917_),
    .B(_05281_),
    .C(_05637_),
    .Y(_05638_));
 sg13g2_o21ai_1 _19219_ (.B1(_05607_),
    .Y(_05639_),
    .A1(_05636_),
    .A2(_05638_));
 sg13g2_o21ai_1 _19220_ (.B1(_05639_),
    .Y(_05640_),
    .A1(net6992),
    .A2(_05634_));
 sg13g2_xnor2_1 _19221_ (.Y(_05641_),
    .A(net6939),
    .B(_05444_));
 sg13g2_nand3_1 _19222_ (.B(_05285_),
    .C(_05641_),
    .A(net7002),
    .Y(_05642_));
 sg13g2_nor2_1 _19223_ (.A(net6994),
    .B(net6945),
    .Y(_05643_));
 sg13g2_xnor2_1 _19224_ (.Y(_05644_),
    .A(net6996),
    .B(net6945));
 sg13g2_nand3_1 _19225_ (.B(_05445_),
    .C(_05644_),
    .A(net6997),
    .Y(_05645_));
 sg13g2_a21oi_1 _19226_ (.A1(_05642_),
    .A2(_05645_),
    .Y(_05646_),
    .B1(_05610_));
 sg13g2_o21ai_1 _19227_ (.B1(net6993),
    .Y(_05647_),
    .A1(_05445_),
    .A2(_05609_));
 sg13g2_a22oi_1 _19228_ (.Y(_05648_),
    .B1(_05647_),
    .B2(net7000),
    .A2(_05610_),
    .A1(net7058));
 sg13g2_nor2_1 _19229_ (.A(net6939),
    .B(_05648_),
    .Y(_05649_));
 sg13g2_o21ai_1 _19230_ (.B1(_05632_),
    .Y(_05650_),
    .A1(_05646_),
    .A2(_05649_));
 sg13g2_nor2_1 _19231_ (.A(_05632_),
    .B(_05640_),
    .Y(_05651_));
 sg13g2_xor2_1 _19232_ (.B(_05640_),
    .A(_05632_),
    .X(_05652_));
 sg13g2_a21oi_1 _19233_ (.A1(_01658_),
    .A2(net7322),
    .Y(_05653_),
    .B1(_05018_));
 sg13g2_a21o_1 _19234_ (.A2(net7323),
    .A1(_01658_),
    .B1(net7314),
    .X(_05654_));
 sg13g2_o21ai_1 _19235_ (.B1(_05610_),
    .Y(_05655_),
    .A1(net7117),
    .A2(net6991));
 sg13g2_a21oi_1 _19236_ (.A1(_05445_),
    .A2(_05610_),
    .Y(_05656_),
    .B1(net6936));
 sg13g2_o21ai_1 _19237_ (.B1(net6993),
    .Y(_05657_),
    .A1(_05611_),
    .A2(_05656_));
 sg13g2_nor2_1 _19238_ (.A(net6943),
    .B(_05610_),
    .Y(_05658_));
 sg13g2_nor2_1 _19239_ (.A(net6938),
    .B(_05609_),
    .Y(_05659_));
 sg13g2_mux2_1 _19240_ (.A0(_05658_),
    .A1(_05659_),
    .S(net6993),
    .X(_05660_));
 sg13g2_nand3_1 _19241_ (.B(_05655_),
    .C(_05657_),
    .A(net7000),
    .Y(_05661_));
 sg13g2_o21ai_1 _19242_ (.B1(_05661_),
    .Y(_05662_),
    .A1(net7000),
    .A2(_05660_));
 sg13g2_xnor2_1 _19243_ (.Y(_05663_),
    .A(_05654_),
    .B(_05662_));
 sg13g2_xnor2_1 _19244_ (.Y(_05664_),
    .A(_05652_),
    .B(_05663_));
 sg13g2_nor2_1 _19245_ (.A(net7176),
    .B(net7141),
    .Y(_05665_));
 sg13g2_nor2_1 _19246_ (.A(net7182),
    .B(_04649_),
    .Y(_05666_));
 sg13g2_xor2_1 _19247_ (.B(_05666_),
    .A(_05665_),
    .X(_05667_));
 sg13g2_nand2_1 _19248_ (.Y(_05668_),
    .A(net7189),
    .B(net7062));
 sg13g2_xnor2_1 _19249_ (.Y(_05669_),
    .A(_05667_),
    .B(_05668_));
 sg13g2_nand2_1 _19250_ (.Y(_05670_),
    .A(_05529_),
    .B(_05530_));
 sg13g2_nor2_1 _19251_ (.A(_05529_),
    .B(_05530_),
    .Y(_05671_));
 sg13g2_o21ai_1 _19252_ (.B1(_05670_),
    .Y(_05672_),
    .A1(_05532_),
    .A2(_05671_));
 sg13g2_nor2_1 _19253_ (.A(net7160),
    .B(net7146),
    .Y(_05673_));
 sg13g2_nor2_1 _19254_ (.A(_04297_),
    .B(net7150),
    .Y(_05674_));
 sg13g2_nor2_1 _19255_ (.A(net7157),
    .B(net7155),
    .Y(_05675_));
 sg13g2_xnor2_1 _19256_ (.Y(_05676_),
    .A(_05674_),
    .B(_05675_));
 sg13g2_xnor2_1 _19257_ (.Y(_05677_),
    .A(_05673_),
    .B(_05676_));
 sg13g2_nand2_1 _19258_ (.Y(_05678_),
    .A(_05672_),
    .B(_05677_));
 sg13g2_or2_1 _19259_ (.X(_05679_),
    .B(_05677_),
    .A(_05672_));
 sg13g2_xor2_1 _19260_ (.B(_05677_),
    .A(_05672_),
    .X(_05680_));
 sg13g2_xnor2_1 _19261_ (.Y(_05681_),
    .A(_05669_),
    .B(_05680_));
 sg13g2_xor2_1 _19262_ (.B(_05680_),
    .A(_05669_),
    .X(_05682_));
 sg13g2_a21o_1 _19263_ (.A2(_05541_),
    .A1(_05536_),
    .B1(_05533_),
    .X(_05683_));
 sg13g2_o21ai_1 _19264_ (.B1(_05533_),
    .Y(_05684_),
    .A1(_05536_),
    .A2(_05541_));
 sg13g2_nor2_1 _19265_ (.A(net7179),
    .B(net7131),
    .Y(_05685_));
 sg13g2_nor2_1 _19266_ (.A(net7170),
    .B(net7138),
    .Y(_05686_));
 sg13g2_nor2_1 _19267_ (.A(net7185),
    .B(net7115),
    .Y(_05687_));
 sg13g2_xnor2_1 _19268_ (.Y(_05688_),
    .A(_05686_),
    .B(_05687_));
 sg13g2_xor2_1 _19269_ (.B(_05688_),
    .A(_05685_),
    .X(_05689_));
 sg13g2_xnor2_1 _19270_ (.Y(_05690_),
    .A(_05685_),
    .B(_05688_));
 sg13g2_or2_1 _19271_ (.X(_05691_),
    .B(_05549_),
    .A(_05548_));
 sg13g2_nand2_1 _19272_ (.Y(_05692_),
    .A(_05548_),
    .B(_05549_));
 sg13g2_a21o_1 _19273_ (.A2(_05549_),
    .A1(_05548_),
    .B1(_05547_),
    .X(_05693_));
 sg13g2_o21ai_1 _19274_ (.B1(_05547_),
    .Y(_05694_),
    .A1(_05548_),
    .A2(_05549_));
 sg13g2_nand2_1 _19275_ (.Y(_05695_),
    .A(_05691_),
    .B(_05693_));
 sg13g2_nand2_1 _19276_ (.Y(_05696_),
    .A(_05537_),
    .B(_05538_));
 sg13g2_or2_1 _19277_ (.X(_05697_),
    .B(_05538_),
    .A(_05537_));
 sg13g2_o21ai_1 _19278_ (.B1(_05539_),
    .Y(_05698_),
    .A1(_05537_),
    .A2(_05538_));
 sg13g2_a21o_1 _19279_ (.A2(_05538_),
    .A1(_05537_),
    .B1(_05539_),
    .X(_05699_));
 sg13g2_nand2_1 _19280_ (.Y(_05700_),
    .A(_05696_),
    .B(_05698_));
 sg13g2_a22oi_1 _19281_ (.Y(_05701_),
    .B1(_05697_),
    .B2(_05699_),
    .A2(_05693_),
    .A1(_05691_));
 sg13g2_nand4_1 _19282_ (.B(_05694_),
    .C(_05696_),
    .A(_05692_),
    .Y(_05702_),
    .D(_05698_));
 sg13g2_a22oi_1 _19283_ (.Y(_05703_),
    .B1(_05696_),
    .B2(_05698_),
    .A2(_05694_),
    .A1(_05692_));
 sg13g2_nand4_1 _19284_ (.B(_05693_),
    .C(_05697_),
    .A(_05691_),
    .Y(_05704_),
    .D(_05699_));
 sg13g2_nand3_1 _19285_ (.B(_05702_),
    .C(_05704_),
    .A(_05689_),
    .Y(_05705_));
 sg13g2_o21ai_1 _19286_ (.B1(_05690_),
    .Y(_05706_),
    .A1(_05701_),
    .A2(_05703_));
 sg13g2_nand3_1 _19287_ (.B(_05702_),
    .C(_05704_),
    .A(_05690_),
    .Y(_05707_));
 sg13g2_o21ai_1 _19288_ (.B1(_05689_),
    .Y(_05708_),
    .A1(_05701_),
    .A2(_05703_));
 sg13g2_a22oi_1 _19289_ (.Y(_05709_),
    .B1(_05707_),
    .B2(_05708_),
    .A2(_05683_),
    .A1(_05542_));
 sg13g2_nand4_1 _19290_ (.B(_05684_),
    .C(_05705_),
    .A(_05543_),
    .Y(_05710_),
    .D(_05706_));
 sg13g2_a22oi_1 _19291_ (.Y(_05711_),
    .B1(_05705_),
    .B2(_05706_),
    .A2(_05684_),
    .A1(_05543_));
 sg13g2_nand4_1 _19292_ (.B(_05683_),
    .C(_05707_),
    .A(_05542_),
    .Y(_05712_),
    .D(_05708_));
 sg13g2_a21oi_1 _19293_ (.A1(_05710_),
    .A2(_05712_),
    .Y(_05713_),
    .B1(_05682_));
 sg13g2_nor3_1 _19294_ (.A(_05681_),
    .B(_05709_),
    .C(_05711_),
    .Y(_05714_));
 sg13g2_or2_1 _19295_ (.X(_05715_),
    .B(_05714_),
    .A(_05713_));
 sg13g2_a21oi_1 _19296_ (.A1(_05545_),
    .A2(_05561_),
    .Y(_05716_),
    .B1(_05562_));
 sg13g2_xnor2_1 _19297_ (.Y(_05717_),
    .A(_05715_),
    .B(_05716_));
 sg13g2_nand2_1 _19298_ (.Y(_05718_),
    .A(_05555_),
    .B(_05558_));
 sg13g2_o21ai_1 _19299_ (.B1(_05551_),
    .Y(_05719_),
    .A1(_05555_),
    .A2(_05558_));
 sg13g2_nand2_1 _19300_ (.Y(_05720_),
    .A(_05718_),
    .B(_05719_));
 sg13g2_nand3_1 _19301_ (.B(_05215_),
    .C(_05573_),
    .A(net7227),
    .Y(_05721_));
 sg13g2_nand4_1 _19302_ (.B(_05089_),
    .C(_05090_),
    .A(_03863_),
    .Y(_05722_),
    .D(_05573_));
 sg13g2_nand3_1 _19303_ (.B(_05216_),
    .C(_05574_),
    .A(_05214_),
    .Y(_05723_));
 sg13g2_inv_1 _19304_ (.Y(_05724_),
    .A(_05725_));
 sg13g2_nand4_1 _19305_ (.B(_05721_),
    .C(_05722_),
    .A(_04797_),
    .Y(_05725_),
    .D(_05723_));
 sg13g2_xnor2_1 _19306_ (.Y(_05726_),
    .A(net7004),
    .B(_05184_));
 sg13g2_xnor2_1 _19307_ (.Y(_05727_),
    .A(net6894),
    .B(_05726_));
 sg13g2_xor2_1 _19308_ (.B(_05727_),
    .A(_05720_),
    .X(_05728_));
 sg13g2_xnor2_1 _19309_ (.Y(_05729_),
    .A(_05717_),
    .B(_05728_));
 sg13g2_o21ai_1 _19310_ (.B1(_05587_),
    .Y(_05730_),
    .A1(_05583_),
    .A2(_05588_));
 sg13g2_xnor2_1 _19311_ (.Y(_05731_),
    .A(_05729_),
    .B(_05730_));
 sg13g2_xnor2_1 _19312_ (.Y(_05732_),
    .A(_05664_),
    .B(_05731_));
 sg13g2_and2_1 _19313_ (.A(_05590_),
    .B(_05591_),
    .X(_05733_));
 sg13g2_or2_1 _19314_ (.X(_05734_),
    .B(_05591_),
    .A(_05590_));
 sg13g2_a21oi_1 _19315_ (.A1(_05623_),
    .A2(_05734_),
    .Y(_05735_),
    .B1(_05733_));
 sg13g2_nor2_1 _19316_ (.A(_05595_),
    .B(_05619_),
    .Y(_05736_));
 sg13g2_nor2_1 _19317_ (.A(_05622_),
    .B(_05736_),
    .Y(_05737_));
 sg13g2_a21oi_1 _19318_ (.A1(_05595_),
    .A2(_05619_),
    .Y(_05738_),
    .B1(_05737_));
 sg13g2_nor2_1 _19319_ (.A(_05735_),
    .B(_05738_),
    .Y(_05739_));
 sg13g2_xor2_1 _19320_ (.B(_05738_),
    .A(_05732_),
    .X(_05740_));
 sg13g2_xnor2_1 _19321_ (.Y(_05741_),
    .A(_05735_),
    .B(_05740_));
 sg13g2_inv_1 _19322_ (.Y(_05742_),
    .A(_00376_));
 sg13g2_xnor2_1 _19323_ (.Y(_05743_),
    .A(_05720_),
    .B(_05724_));
 sg13g2_inv_1 _19324_ (.Y(_05744_),
    .A(_00375_));
 sg13g2_xnor2_1 _19325_ (.Y(_05745_),
    .A(_05717_),
    .B(net6829));
 sg13g2_or2_1 _19326_ (.X(_05746_),
    .B(_05745_),
    .A(_05730_));
 sg13g2_and2_1 _19327_ (.A(_05730_),
    .B(_05745_),
    .X(_05747_));
 sg13g2_xor2_1 _19328_ (.B(net6892),
    .A(_05664_),
    .X(_05748_));
 sg13g2_o21ai_1 _19329_ (.B1(_05746_),
    .Y(_05749_),
    .A1(_05747_),
    .A2(_05748_));
 sg13g2_nor3_1 _19330_ (.A(_05713_),
    .B(_05714_),
    .C(_05743_),
    .Y(_05750_));
 sg13g2_o21ai_1 _19331_ (.B1(net6829),
    .Y(_05751_),
    .A1(_05713_),
    .A2(_05714_));
 sg13g2_inv_1 _19332_ (.Y(_05752_),
    .A(_00372_));
 sg13g2_o21ai_1 _19333_ (.B1(_05751_),
    .Y(_05753_),
    .A1(_05716_),
    .A2(_05750_));
 sg13g2_a21oi_1 _19334_ (.A1(_01659_),
    .A2(net7323),
    .Y(_05754_),
    .B1(net7314));
 sg13g2_a21o_1 _19335_ (.A2(net7323),
    .A1(_01659_),
    .B1(net7314),
    .X(_05755_));
 sg13g2_o21ai_1 _19336_ (.B1(_05653_),
    .Y(_05756_),
    .A1(net7117),
    .A2(net6991));
 sg13g2_nor2_1 _19337_ (.A(net6994),
    .B(_05756_),
    .Y(_05757_));
 sg13g2_nor3_1 _19338_ (.A(_04798_),
    .B(_05182_),
    .C(_05653_),
    .Y(_05758_));
 sg13g2_a21oi_1 _19339_ (.A1(net6994),
    .A2(_05758_),
    .Y(_05759_),
    .B1(_05757_));
 sg13g2_nor2_1 _19340_ (.A(_05609_),
    .B(_05653_),
    .Y(_05760_));
 sg13g2_o21ai_1 _19341_ (.B1(_05655_),
    .Y(_05761_),
    .A1(net6938),
    .A2(_05760_));
 sg13g2_a221oi_1 _19342_ (.B2(net6994),
    .C1(net6999),
    .B1(_05761_),
    .A1(net6938),
    .Y(_05762_),
    .A2(_05654_));
 sg13g2_a21oi_1 _19343_ (.A1(net6999),
    .A2(_05759_),
    .Y(_05763_),
    .B1(_05762_));
 sg13g2_xnor2_1 _19344_ (.Y(_05764_),
    .A(net7113),
    .B(_05763_));
 sg13g2_xnor2_1 _19345_ (.Y(_05765_),
    .A(_05753_),
    .B(_05764_));
 sg13g2_nor2_1 _19346_ (.A(net7160),
    .B(net7141),
    .Y(_05766_));
 sg13g2_nor2_1 _19347_ (.A(net7176),
    .B(_04649_),
    .Y(_05767_));
 sg13g2_xnor2_1 _19348_ (.Y(_05768_),
    .A(_05766_),
    .B(_05767_));
 sg13g2_and2_1 _19349_ (.A(net7182),
    .B(_04737_),
    .X(_05769_));
 sg13g2_xnor2_1 _19350_ (.Y(_05770_),
    .A(_05768_),
    .B(_05769_));
 sg13g2_nor2_1 _19351_ (.A(_05665_),
    .B(_05666_),
    .Y(_05771_));
 sg13g2_a22oi_1 _19352_ (.Y(_05772_),
    .B1(_05665_),
    .B2(_05666_),
    .A2(net7062),
    .A1(net7189));
 sg13g2_nor2_1 _19353_ (.A(_05771_),
    .B(_05772_),
    .Y(_05773_));
 sg13g2_or2_1 _19354_ (.X(_05774_),
    .B(_05772_),
    .A(_05771_));
 sg13g2_nor2_1 _19355_ (.A(net7154),
    .B(net7150),
    .Y(_05775_));
 sg13g2_nor2_1 _19356_ (.A(net7166),
    .B(net7138),
    .Y(_05776_));
 sg13g2_nor2_1 _19357_ (.A(net7157),
    .B(net7146),
    .Y(_05777_));
 sg13g2_xnor2_1 _19358_ (.Y(_05778_),
    .A(_05775_),
    .B(_05777_));
 sg13g2_xor2_1 _19359_ (.B(_05778_),
    .A(_05776_),
    .X(_05779_));
 sg13g2_xnor2_1 _19360_ (.Y(_05780_),
    .A(_05776_),
    .B(_05778_));
 sg13g2_xnor2_1 _19361_ (.Y(_05781_),
    .A(_05773_),
    .B(_05779_));
 sg13g2_xnor2_1 _19362_ (.Y(_05782_),
    .A(_05770_),
    .B(_05781_));
 sg13g2_xor2_1 _19363_ (.B(_05781_),
    .A(_05770_),
    .X(_05783_));
 sg13g2_nor2_1 _19364_ (.A(net7171),
    .B(net7061),
    .Y(_05784_));
 sg13g2_nand3b_1 _19365_ (.B(net7133),
    .C(net7179),
    .Y(_05785_),
    .A_N(net7171));
 sg13g2_nand3b_1 _19366_ (.B(net7171),
    .C(_04797_),
    .Y(_05786_),
    .A_N(net7179));
 sg13g2_a21oi_1 _19367_ (.A1(_05785_),
    .A2(_05786_),
    .Y(_05787_),
    .B1(_04130_));
 sg13g2_inv_1 _19368_ (.Y(_05788_),
    .A(_05789_));
 sg13g2_or2_1 _19369_ (.X(_05789_),
    .B(net7170),
    .A(net7179));
 sg13g2_o21ai_1 _19370_ (.B1(net7178),
    .Y(_05790_),
    .A1(net7170),
    .A2(net7131));
 sg13g2_nand2_1 _19371_ (.Y(_05791_),
    .A(_05789_),
    .B(_05790_));
 sg13g2_a221oi_1 _19372_ (.B2(_05687_),
    .C1(_05787_),
    .B1(_05791_),
    .A1(net7133),
    .Y(_05792_),
    .A2(_05784_));
 sg13g2_o21ai_1 _19373_ (.B1(_05674_),
    .Y(_05793_),
    .A1(_05673_),
    .A2(_05675_));
 sg13g2_nand2_1 _19374_ (.Y(_05794_),
    .A(_05673_),
    .B(_05675_));
 sg13g2_nor4_1 _19375_ (.A(net7178),
    .B(net7170),
    .C(net7138),
    .D(net7131),
    .Y(_05795_));
 sg13g2_nor4_1 _19376_ (.A(net7185),
    .B(net7179),
    .C(net7131),
    .D(net7120),
    .Y(_05796_));
 sg13g2_a21oi_1 _19377_ (.A1(_05674_),
    .A2(_05675_),
    .Y(_05797_),
    .B1(_05673_));
 sg13g2_nor2_1 _19378_ (.A(_05674_),
    .B(_05675_),
    .Y(_05798_));
 sg13g2_nor4_1 _19379_ (.A(net7185),
    .B(net7171),
    .C(net7138),
    .D(net7115),
    .Y(_05799_));
 sg13g2_nor3_1 _19380_ (.A(_05795_),
    .B(_05796_),
    .C(_05799_),
    .Y(_05800_));
 sg13g2_and3_1 _19381_ (.X(_05801_),
    .A(_05793_),
    .B(_05794_),
    .C(_05800_));
 sg13g2_o21ai_1 _19382_ (.B1(_05800_),
    .Y(_05802_),
    .A1(_05797_),
    .A2(_05798_));
 sg13g2_nor3_1 _19383_ (.A(_05797_),
    .B(_05798_),
    .C(_05800_),
    .Y(_05803_));
 sg13g2_or3_1 _19384_ (.A(_05797_),
    .B(_05798_),
    .C(_05800_),
    .X(_05804_));
 sg13g2_nand3_1 _19385_ (.B(_05802_),
    .C(_05804_),
    .A(_05792_),
    .Y(_05805_));
 sg13g2_a21o_1 _19386_ (.A2(_05804_),
    .A1(_05802_),
    .B1(_05792_),
    .X(_05806_));
 sg13g2_nand3b_1 _19387_ (.B(_05802_),
    .C(_05804_),
    .Y(_05807_),
    .A_N(_05792_));
 sg13g2_o21ai_1 _19388_ (.B1(net6933),
    .Y(_05808_),
    .A1(_05801_),
    .A2(_05803_));
 sg13g2_nand2_1 _19389_ (.Y(_05809_),
    .A(_05805_),
    .B(_05806_));
 sg13g2_o21ai_1 _19390_ (.B1(_05669_),
    .Y(_05810_),
    .A1(_05672_),
    .A2(_05677_));
 sg13g2_a21o_1 _19391_ (.A2(_05677_),
    .A1(_05672_),
    .B1(_05669_),
    .X(_05811_));
 sg13g2_nand2_1 _19392_ (.Y(_05812_),
    .A(_05678_),
    .B(_05810_));
 sg13g2_nand2_1 _19393_ (.Y(_05813_),
    .A(_05679_),
    .B(_05811_));
 sg13g2_nand4_1 _19394_ (.B(_05805_),
    .C(_05806_),
    .A(_05679_),
    .Y(_05814_),
    .D(_05811_));
 sg13g2_nand4_1 _19395_ (.B(_05807_),
    .C(_05808_),
    .A(_05678_),
    .Y(_05815_),
    .D(_05810_));
 sg13g2_nand3_1 _19396_ (.B(_05814_),
    .C(_05815_),
    .A(_05783_),
    .Y(_05816_));
 sg13g2_a21o_1 _19397_ (.A2(_05815_),
    .A1(_05814_),
    .B1(_05783_),
    .X(_05817_));
 sg13g2_nand2_1 _19398_ (.Y(_05818_),
    .A(_05695_),
    .B(_05700_));
 sg13g2_o21ai_1 _19399_ (.B1(_05690_),
    .Y(_05819_),
    .A1(_05695_),
    .A2(_05700_));
 sg13g2_nand2_1 _19400_ (.Y(_05820_),
    .A(_05818_),
    .B(_05819_));
 sg13g2_xor2_1 _19401_ (.B(net6859),
    .A(_05727_),
    .X(_05821_));
 sg13g2_o21ai_1 _19402_ (.B1(_05712_),
    .Y(_05822_),
    .A1(_05682_),
    .A2(_05709_));
 sg13g2_a21oi_1 _19403_ (.A1(_05681_),
    .A2(_05710_),
    .Y(_05823_),
    .B1(_05711_));
 sg13g2_a21oi_1 _19404_ (.A1(_05816_),
    .A2(_05817_),
    .Y(_05824_),
    .B1(_05822_));
 sg13g2_and3_1 _19405_ (.X(_05825_),
    .A(_05816_),
    .B(_05817_),
    .C(_05822_));
 sg13g2_nor2_1 _19406_ (.A(_05824_),
    .B(_05825_),
    .Y(_05826_));
 sg13g2_inv_1 _19407_ (.Y(_05827_),
    .A(_00348_));
 sg13g2_inv_1 _19408_ (.Y(_05828_),
    .A(\load_store_unit_i.lsu_err_q ));
 sg13g2_inv_1 _19409_ (.Y(_05829_),
    .A(_00347_));
 sg13g2_inv_1 _19410_ (.Y(_05830_),
    .A(_00346_));
 sg13g2_a22oi_1 _19411_ (.Y(_05831_),
    .B1(_05214_),
    .B2(_05216_),
    .A2(net7196),
    .A1(net7203));
 sg13g2_a22oi_1 _19412_ (.Y(_05832_),
    .B1(_05215_),
    .B2(net7227),
    .A2(_04022_),
    .A1(_03971_));
 sg13g2_a21oi_1 _19413_ (.A1(_05214_),
    .A2(_05832_),
    .Y(_05833_),
    .B1(net7207));
 sg13g2_inv_1 _19414_ (.Y(_05834_),
    .A(net6891));
 sg13g2_o21ai_1 _19415_ (.B1(net7118),
    .Y(_05835_),
    .A1(_05831_),
    .A2(_05833_));
 sg13g2_nand3_1 _19416_ (.B(_05719_),
    .C(_05835_),
    .A(_05718_),
    .Y(_05836_));
 sg13g2_a221oi_1 _19417_ (.B2(_05019_),
    .C1(_05654_),
    .B1(_05443_),
    .A1(net7119),
    .Y(_05837_),
    .A2(_05183_));
 sg13g2_nor2_1 _19418_ (.A(net7058),
    .B(_05610_),
    .Y(_05838_));
 sg13g2_o21ai_1 _19419_ (.B1(_05838_),
    .Y(_05839_),
    .A1(_05758_),
    .A2(_05837_));
 sg13g2_nand2_1 _19420_ (.Y(_05840_),
    .A(_05609_),
    .B(_05654_));
 sg13g2_a21oi_1 _19421_ (.A1(net7119),
    .A2(_05183_),
    .Y(_05841_),
    .B1(_05840_));
 sg13g2_nor3_1 _19422_ (.A(net7117),
    .B(_05182_),
    .C(_05654_),
    .Y(_05842_));
 sg13g2_o21ai_1 _19423_ (.B1(net7057),
    .Y(_05843_),
    .A1(_05841_),
    .A2(_05842_));
 sg13g2_nor2_1 _19424_ (.A(_05609_),
    .B(_05654_),
    .Y(_05844_));
 sg13g2_nand3_1 _19425_ (.B(_05445_),
    .C(_05844_),
    .A(_05184_),
    .Y(_05845_));
 sg13g2_and3_1 _19426_ (.X(_05846_),
    .A(_05839_),
    .B(_05843_),
    .C(_05845_));
 sg13g2_a21o_1 _19427_ (.A2(_05844_),
    .A1(net6939),
    .B1(_05758_),
    .X(_05847_));
 sg13g2_a221oi_1 _19428_ (.B2(net7057),
    .C1(net7002),
    .B1(_05847_),
    .A1(_05418_),
    .Y(_05848_),
    .A2(_05844_));
 sg13g2_a21oi_1 _19429_ (.A1(net7003),
    .A2(_05846_),
    .Y(_05849_),
    .B1(_05848_));
 sg13g2_a21oi_1 _19430_ (.A1(_05718_),
    .A2(_05719_),
    .Y(_05850_),
    .B1(_05835_));
 sg13g2_o21ai_1 _19431_ (.B1(_05836_),
    .Y(_05851_),
    .A1(net6895),
    .A2(_05850_));
 sg13g2_xnor2_1 _19432_ (.Y(_05852_),
    .A(_05849_),
    .B(_05851_));
 sg13g2_xnor2_1 _19433_ (.Y(_05853_),
    .A(_05821_),
    .B(_05852_));
 sg13g2_xnor2_1 _19434_ (.Y(_05854_),
    .A(_05826_),
    .B(_05853_));
 sg13g2_xnor2_1 _19435_ (.Y(_05855_),
    .A(_05765_),
    .B(_05854_));
 sg13g2_xor2_1 _19436_ (.B(net6892),
    .A(_05663_),
    .X(_05856_));
 sg13g2_o21ai_1 _19437_ (.B1(_05650_),
    .Y(_05857_),
    .A1(_05651_),
    .A2(_05856_));
 sg13g2_inv_1 _19438_ (.Y(_05858_),
    .A(net7657));
 sg13g2_nor2_1 _19439_ (.A(_05855_),
    .B(_05857_),
    .Y(_05859_));
 sg13g2_xor2_1 _19440_ (.B(_05857_),
    .A(_05855_),
    .X(_05860_));
 sg13g2_xnor2_1 _19441_ (.Y(_05861_),
    .A(_05749_),
    .B(_05860_));
 sg13g2_xnor2_1 _19442_ (.Y(_05862_),
    .A(_05724_),
    .B(_05820_));
 sg13g2_xor2_1 _19443_ (.B(_05862_),
    .A(_05826_),
    .X(_05863_));
 sg13g2_xnor2_1 _19444_ (.Y(_05864_),
    .A(net6893),
    .B(_05764_));
 sg13g2_xnor2_1 _19445_ (.Y(_05865_),
    .A(_05852_),
    .B(_05864_));
 sg13g2_o21ai_1 _19446_ (.B1(_05753_),
    .Y(_05866_),
    .A1(_05863_),
    .A2(_05865_));
 sg13g2_nand2_1 _19447_ (.Y(_05867_),
    .A(_05863_),
    .B(_05865_));
 sg13g2_nand2_1 _19448_ (.Y(_05868_),
    .A(_05866_),
    .B(_05867_));
 sg13g2_nand2_1 _19449_ (.Y(_05869_),
    .A(net6943),
    .B(_05755_));
 sg13g2_nor2_1 _19450_ (.A(_05653_),
    .B(_05755_),
    .Y(_05870_));
 sg13g2_nand2_1 _19451_ (.Y(_05871_),
    .A(net6938),
    .B(_05870_));
 sg13g2_nand2_1 _19452_ (.Y(_05872_),
    .A(_05869_),
    .B(_05871_));
 sg13g2_a221oi_1 _19453_ (.B2(net7055),
    .C1(net7001),
    .B1(_05872_),
    .A1(net6897),
    .Y(_05873_),
    .A2(_05870_));
 sg13g2_o21ai_1 _19454_ (.B1(_05869_),
    .Y(_05874_),
    .A1(_05655_),
    .A2(_05755_));
 sg13g2_nor2_1 _19455_ (.A(net7055),
    .B(_05654_),
    .Y(_05875_));
 sg13g2_a22oi_1 _19456_ (.Y(_05876_),
    .B1(_05874_),
    .B2(_05875_),
    .A2(_05870_),
    .A1(_05659_));
 sg13g2_a21o_1 _19457_ (.A2(_05876_),
    .A1(net7001),
    .B1(_05873_),
    .X(_05877_));
 sg13g2_a21o_1 _19458_ (.A2(_05834_),
    .A1(net6859),
    .B1(net6895),
    .X(_05878_));
 sg13g2_o21ai_1 _19459_ (.B1(_05878_),
    .Y(_05879_),
    .A1(net6859),
    .A2(_05834_));
 sg13g2_xor2_1 _19460_ (.B(_05879_),
    .A(_05877_),
    .X(_05880_));
 sg13g2_a21oi_1 _19461_ (.A1(_01661_),
    .A2(net7323),
    .Y(_05881_),
    .B1(_05018_));
 sg13g2_a21o_1 _19462_ (.A2(net7322),
    .A1(_01661_),
    .B1(net7317),
    .X(_05882_));
 sg13g2_nand3_1 _19463_ (.B(net7113),
    .C(_05756_),
    .A(net6994),
    .Y(_05883_));
 sg13g2_nand2_1 _19464_ (.Y(_05884_),
    .A(_05653_),
    .B(_05755_));
 sg13g2_nor2_1 _19465_ (.A(_05091_),
    .B(_05754_),
    .Y(_05885_));
 sg13g2_nor3_1 _19466_ (.A(_03863_),
    .B(_05092_),
    .C(_05754_),
    .Y(_05886_));
 sg13g2_nor2_1 _19467_ (.A(_05885_),
    .B(_05886_),
    .Y(_05887_));
 sg13g2_nand4_1 _19468_ (.B(_05883_),
    .C(_05884_),
    .A(net7003),
    .Y(_05888_),
    .D(_05887_));
 sg13g2_mux2_1 _19469_ (.A0(_05418_),
    .A1(_05643_),
    .S(net7113),
    .X(_05889_));
 sg13g2_o21ai_1 _19470_ (.B1(_05888_),
    .Y(_05890_),
    .A1(net7003),
    .A2(_05889_));
 sg13g2_xnor2_1 _19471_ (.Y(_05891_),
    .A(_05882_),
    .B(_05890_));
 sg13g2_xnor2_1 _19472_ (.Y(_05892_),
    .A(_05880_),
    .B(_05891_));
 sg13g2_nor2_1 _19473_ (.A(_05783_),
    .B(_05812_),
    .Y(_05893_));
 sg13g2_nand2_1 _19474_ (.Y(_05894_),
    .A(_05783_),
    .B(_05812_));
 sg13g2_a21oi_1 _19475_ (.A1(_05783_),
    .A2(_05812_),
    .Y(_05895_),
    .B1(_05809_));
 sg13g2_a21o_1 _19476_ (.A2(_05812_),
    .A1(_05783_),
    .B1(_05809_),
    .X(_05896_));
 sg13g2_o21ai_1 _19477_ (.B1(_05809_),
    .Y(_05897_),
    .A1(_05783_),
    .A2(_05812_));
 sg13g2_nor2_1 _19478_ (.A(net7157),
    .B(net7141),
    .Y(_05898_));
 sg13g2_nor2_1 _19479_ (.A(net7160),
    .B(_04649_),
    .Y(_05899_));
 sg13g2_xor2_1 _19480_ (.B(_05899_),
    .A(_05898_),
    .X(_05900_));
 sg13g2_nand2_1 _19481_ (.Y(_05901_),
    .A(net7176),
    .B(net7062));
 sg13g2_xnor2_1 _19482_ (.Y(_05902_),
    .A(_05900_),
    .B(_05901_));
 sg13g2_and2_1 _19483_ (.A(_05766_),
    .B(_05767_),
    .X(_05903_));
 sg13g2_or2_1 _19484_ (.X(_05904_),
    .B(_05767_),
    .A(_05766_));
 sg13g2_a21o_1 _19485_ (.A2(_05904_),
    .A1(_05769_),
    .B1(_05903_),
    .X(_05905_));
 sg13g2_a21oi_1 _19486_ (.A1(_05769_),
    .A2(_05904_),
    .Y(_05906_),
    .B1(_05903_));
 sg13g2_nor2_1 _19487_ (.A(net7165),
    .B(net7132),
    .Y(_05907_));
 sg13g2_nor2_1 _19488_ (.A(net7150),
    .B(net7146),
    .Y(_05908_));
 sg13g2_nor2_1 _19489_ (.A(net7154),
    .B(net7138),
    .Y(_05909_));
 sg13g2_xnor2_1 _19490_ (.Y(_05910_),
    .A(_05908_),
    .B(_05909_));
 sg13g2_xor2_1 _19491_ (.B(_05910_),
    .A(_05907_),
    .X(_05911_));
 sg13g2_xnor2_1 _19492_ (.Y(_05912_),
    .A(_05907_),
    .B(_05910_));
 sg13g2_xnor2_1 _19493_ (.Y(_05913_),
    .A(_05905_),
    .B(_05911_));
 sg13g2_xnor2_1 _19494_ (.Y(_05914_),
    .A(_05902_),
    .B(_05913_));
 sg13g2_a21o_1 _19495_ (.A2(_05780_),
    .A1(_05773_),
    .B1(_05770_),
    .X(_05915_));
 sg13g2_nand2_1 _19496_ (.Y(_05916_),
    .A(_05775_),
    .B(_05777_));
 sg13g2_o21ai_1 _19497_ (.B1(_05776_),
    .Y(_05917_),
    .A1(_05775_),
    .A2(_05777_));
 sg13g2_nand2_1 _19498_ (.Y(_05918_),
    .A(_05916_),
    .B(_05917_));
 sg13g2_nor3_1 _19499_ (.A(net7185),
    .B(net7178),
    .C(net7170),
    .Y(_05919_));
 sg13g2_nand2_1 _19500_ (.Y(_05920_),
    .A(net7178),
    .B(net7170));
 sg13g2_and3_1 _19501_ (.X(_05921_),
    .A(net7185),
    .B(net7178),
    .C(net7170));
 sg13g2_nor3_1 _19502_ (.A(net7120),
    .B(_05919_),
    .C(_05921_),
    .Y(_05922_));
 sg13g2_or3_1 _19503_ (.A(net7120),
    .B(_05919_),
    .C(_05921_),
    .X(_05923_));
 sg13g2_nor3_1 _19504_ (.A(net7115),
    .B(_05919_),
    .C(_05921_),
    .Y(_05924_));
 sg13g2_a21o_1 _19505_ (.A2(_05917_),
    .A1(_05916_),
    .B1(_05922_),
    .X(_05925_));
 sg13g2_nand3_1 _19506_ (.B(_05917_),
    .C(_05922_),
    .A(_05916_),
    .Y(_05926_));
 sg13g2_nand3_1 _19507_ (.B(_05917_),
    .C(_05923_),
    .A(_05916_),
    .Y(_05927_));
 sg13g2_a21o_1 _19508_ (.A2(_05917_),
    .A1(_05916_),
    .B1(_05923_),
    .X(_05928_));
 sg13g2_a22oi_1 _19509_ (.Y(_05929_),
    .B1(_05925_),
    .B2(_05926_),
    .A2(_05779_),
    .A1(_05774_));
 sg13g2_o21ai_1 _19510_ (.B1(_05770_),
    .Y(_05930_),
    .A1(_05773_),
    .A2(_05780_));
 sg13g2_nand2_1 _19511_ (.Y(_05931_),
    .A(_05915_),
    .B(_05929_));
 sg13g2_a22oi_1 _19512_ (.Y(_05932_),
    .B1(_05927_),
    .B2(_05928_),
    .A2(_05780_),
    .A1(_05773_));
 sg13g2_a22oi_1 _19513_ (.Y(_05933_),
    .B1(_05930_),
    .B2(_05932_),
    .A2(_05929_),
    .A1(_05915_));
 sg13g2_xnor2_1 _19514_ (.Y(_05934_),
    .A(_05914_),
    .B(_05933_));
 sg13g2_nor3_1 _19515_ (.A(_05893_),
    .B(_05895_),
    .C(_05934_),
    .Y(_05935_));
 sg13g2_and3_1 _19516_ (.X(_05936_),
    .A(_05894_),
    .B(_05897_),
    .C(_05934_));
 sg13g2_nor2_1 _19517_ (.A(_05935_),
    .B(_05936_),
    .Y(_05937_));
 sg13g2_a21oi_1 _19518_ (.A1(_05792_),
    .A2(_05804_),
    .Y(_05938_),
    .B1(_05801_));
 sg13g2_xnor2_1 _19519_ (.Y(_05939_),
    .A(_05727_),
    .B(net6890));
 sg13g2_o21ai_1 _19520_ (.B1(_05939_),
    .Y(_05940_),
    .A1(_05935_),
    .A2(_05936_));
 sg13g2_or3_1 _19521_ (.A(_05935_),
    .B(_05936_),
    .C(_05939_),
    .X(_05941_));
 sg13g2_a21oi_1 _19522_ (.A1(_05816_),
    .A2(_05817_),
    .Y(_05942_),
    .B1(_05862_));
 sg13g2_nand3_1 _19523_ (.B(_05817_),
    .C(_05862_),
    .A(_05816_),
    .Y(_05943_));
 sg13g2_a21oi_1 _19524_ (.A1(_05823_),
    .A2(_05943_),
    .Y(_05944_),
    .B1(_05942_));
 sg13g2_nand3_1 _19525_ (.B(_05941_),
    .C(_05944_),
    .A(_05940_),
    .Y(_05945_));
 sg13g2_a21o_1 _19526_ (.A2(_05941_),
    .A1(_05940_),
    .B1(_05944_),
    .X(_05946_));
 sg13g2_nand3_1 _19527_ (.B(_05945_),
    .C(_05946_),
    .A(_05892_),
    .Y(_05947_));
 sg13g2_a21o_1 _19528_ (.A2(_05946_),
    .A1(_05945_),
    .B1(_05892_),
    .X(_05948_));
 sg13g2_nor2_1 _19529_ (.A(_05849_),
    .B(_05864_),
    .Y(_05949_));
 sg13g2_nand2_1 _19530_ (.Y(_05950_),
    .A(_05849_),
    .B(_05864_));
 sg13g2_o21ai_1 _19531_ (.B1(_05950_),
    .Y(_05951_),
    .A1(_05851_),
    .A2(_05949_));
 sg13g2_a21oi_1 _19532_ (.A1(_05947_),
    .A2(_05948_),
    .Y(_05952_),
    .B1(_05951_));
 sg13g2_nand3_1 _19533_ (.B(_05948_),
    .C(_05951_),
    .A(_05947_),
    .Y(_05953_));
 sg13g2_nor2b_1 _19534_ (.A(_05952_),
    .B_N(_05953_),
    .Y(_05954_));
 sg13g2_xnor2_1 _19535_ (.Y(_05955_),
    .A(_05868_),
    .B(_05954_));
 sg13g2_xor2_1 _19536_ (.B(_05938_),
    .A(net6894),
    .X(_05956_));
 sg13g2_inv_1 _19537_ (.Y(_05957_),
    .A(\load_store_unit_i.handle_misaligned_q ));
 sg13g2_xnor2_1 _19538_ (.Y(_05958_),
    .A(_05937_),
    .B(net6858));
 sg13g2_xor2_1 _19539_ (.B(_05891_),
    .A(net6893),
    .X(_05959_));
 sg13g2_xor2_1 _19540_ (.B(_05959_),
    .A(_05880_),
    .X(_05960_));
 sg13g2_nand2_1 _19541_ (.Y(_05961_),
    .A(_05958_),
    .B(_05960_));
 sg13g2_o21ai_1 _19542_ (.B1(_05944_),
    .Y(_05962_),
    .A1(_05958_),
    .A2(_05960_));
 sg13g2_nand2_1 _19543_ (.Y(_05963_),
    .A(_05961_),
    .B(_05962_));
 sg13g2_a22oi_1 _19544_ (.Y(_05964_),
    .B1(_05932_),
    .B2(_05930_),
    .A2(_05931_),
    .A1(_05914_));
 sg13g2_nor2_1 _19545_ (.A(net7154),
    .B(net7132),
    .Y(_05965_));
 sg13g2_nor2_1 _19546_ (.A(net7145),
    .B(net7138),
    .Y(_05966_));
 sg13g2_nor2_1 _19547_ (.A(net7164),
    .B(net7115),
    .Y(_05967_));
 sg13g2_xor2_1 _19548_ (.B(_05967_),
    .A(_05965_),
    .X(_05968_));
 sg13g2_xnor2_1 _19549_ (.Y(_05969_),
    .A(_05966_),
    .B(_05968_));
 sg13g2_nor2_1 _19550_ (.A(_05898_),
    .B(_05899_),
    .Y(_05970_));
 sg13g2_a22oi_1 _19551_ (.Y(_05971_),
    .B1(_05898_),
    .B2(_05899_),
    .A2(net7062),
    .A1(net7176));
 sg13g2_or2_1 _19552_ (.X(_05972_),
    .B(_05971_),
    .A(_05970_));
 sg13g2_nor2_1 _19553_ (.A(net7150),
    .B(net7141),
    .Y(_05973_));
 sg13g2_nor2_1 _19554_ (.A(net7157),
    .B(net7134),
    .Y(_05974_));
 sg13g2_and2_1 _19555_ (.A(net7160),
    .B(_04737_),
    .X(_05975_));
 sg13g2_and2_1 _19556_ (.A(net7160),
    .B(net7062),
    .X(_05976_));
 sg13g2_xor2_1 _19557_ (.B(_05974_),
    .A(_05973_),
    .X(_05977_));
 sg13g2_xnor2_1 _19558_ (.Y(_05978_),
    .A(_05976_),
    .B(_05977_));
 sg13g2_nor2_1 _19559_ (.A(_05972_),
    .B(_05978_),
    .Y(_05979_));
 sg13g2_xnor2_1 _19560_ (.Y(_05980_),
    .A(_05972_),
    .B(_05978_));
 sg13g2_xnor2_1 _19561_ (.Y(_05981_),
    .A(_05969_),
    .B(_05980_));
 sg13g2_a21o_1 _19562_ (.A2(_05912_),
    .A1(_05905_),
    .B1(_05902_),
    .X(_05982_));
 sg13g2_nand2_1 _19563_ (.Y(_05983_),
    .A(_05908_),
    .B(_05909_));
 sg13g2_o21ai_1 _19564_ (.B1(_05907_),
    .Y(_05984_),
    .A1(_05908_),
    .A2(_05909_));
 sg13g2_nand2_1 _19565_ (.Y(_05985_),
    .A(_05983_),
    .B(_05984_));
 sg13g2_a21o_1 _19566_ (.A2(_05984_),
    .A1(_05983_),
    .B1(_05923_),
    .X(_05986_));
 sg13g2_nand3_1 _19567_ (.B(_05983_),
    .C(_05984_),
    .A(_05923_),
    .Y(_05987_));
 sg13g2_nand3_1 _19568_ (.B(_05983_),
    .C(_05984_),
    .A(_05924_),
    .Y(_05988_));
 sg13g2_a21o_1 _19569_ (.A2(_05984_),
    .A1(_05983_),
    .B1(_05924_),
    .X(_05989_));
 sg13g2_a22oi_1 _19570_ (.Y(_05990_),
    .B1(_05988_),
    .B2(_05989_),
    .A2(_05911_),
    .A1(_05906_));
 sg13g2_o21ai_1 _19571_ (.B1(_05902_),
    .Y(_05991_),
    .A1(_05905_),
    .A2(_05912_));
 sg13g2_nand2_1 _19572_ (.Y(_05992_),
    .A(_05982_),
    .B(_05990_));
 sg13g2_a22oi_1 _19573_ (.Y(_05993_),
    .B1(_05986_),
    .B2(_05987_),
    .A2(_05912_),
    .A1(_05905_));
 sg13g2_a22oi_1 _19574_ (.Y(_05994_),
    .B1(_05991_),
    .B2(_05993_),
    .A2(_05990_),
    .A1(_05982_));
 sg13g2_xnor2_1 _19575_ (.Y(_05995_),
    .A(_05981_),
    .B(_05994_));
 sg13g2_xor2_1 _19576_ (.B(_05994_),
    .A(_05981_),
    .X(_05996_));
 sg13g2_nand3_1 _19577_ (.B(_05916_),
    .C(_05917_),
    .A(_05789_),
    .Y(_05997_));
 sg13g2_a22oi_1 _19578_ (.Y(_05998_),
    .B1(_05997_),
    .B2(net7067),
    .A2(_05920_),
    .A1(_05918_));
 sg13g2_nand2b_1 _19579_ (.Y(_05999_),
    .B(net7118),
    .A_N(_05998_));
 sg13g2_xnor2_1 _19580_ (.Y(_06000_),
    .A(_05995_),
    .B(_05999_));
 sg13g2_xnor2_1 _19581_ (.Y(_06001_),
    .A(_05964_),
    .B(_06000_));
 sg13g2_a21oi_1 _19582_ (.A1(_05782_),
    .A2(_05813_),
    .Y(_06002_),
    .B1(_05956_));
 sg13g2_a21o_1 _19583_ (.A2(_06002_),
    .A1(_05896_),
    .B1(_05934_),
    .X(_06003_));
 sg13g2_o21ai_1 _19584_ (.B1(_05956_),
    .Y(_06004_),
    .A1(_05893_),
    .A2(_05895_));
 sg13g2_nand2_1 _19585_ (.Y(_06005_),
    .A(_06003_),
    .B(_06004_));
 sg13g2_nand3_1 _19586_ (.B(_06003_),
    .C(_06004_),
    .A(_05727_),
    .Y(_06006_));
 sg13g2_a21o_1 _19587_ (.A2(_06004_),
    .A1(_06003_),
    .B1(_05727_),
    .X(_06007_));
 sg13g2_and3_1 _19588_ (.X(_06008_),
    .A(_06001_),
    .B(_06006_),
    .C(_06007_));
 sg13g2_a21oi_1 _19589_ (.A1(_06006_),
    .A2(_06007_),
    .Y(_06009_),
    .B1(_06001_));
 sg13g2_a21oi_1 _19590_ (.A1(_01662_),
    .A2(net7322),
    .Y(_06010_),
    .B1(net7317));
 sg13g2_a21o_1 _19591_ (.A2(net7322),
    .A1(_01662_),
    .B1(net7317),
    .X(_06011_));
 sg13g2_o21ai_1 _19592_ (.B1(_05881_),
    .Y(_06012_),
    .A1(net7117),
    .A2(net6991));
 sg13g2_or2_1 _19593_ (.X(_06013_),
    .B(_06012_),
    .A(net6994));
 sg13g2_nor2_1 _19594_ (.A(net6938),
    .B(_05881_),
    .Y(_06014_));
 sg13g2_nand3_1 _19595_ (.B(_05183_),
    .C(_05882_),
    .A(net7119),
    .Y(_06015_));
 sg13g2_o21ai_1 _19596_ (.B1(_06013_),
    .Y(_06016_),
    .A1(net7057),
    .A2(_06015_));
 sg13g2_nor2_1 _19597_ (.A(net7003),
    .B(_06016_),
    .Y(_06017_));
 sg13g2_nand2_1 _19598_ (.Y(_06018_),
    .A(net6937),
    .B(_05882_));
 sg13g2_nor2_1 _19599_ (.A(net6945),
    .B(_05755_),
    .Y(_06019_));
 sg13g2_nor2_1 _19600_ (.A(net7113),
    .B(_05881_),
    .Y(_06020_));
 sg13g2_a21oi_1 _19601_ (.A1(net6945),
    .A2(_06020_),
    .Y(_06021_),
    .B1(_06019_));
 sg13g2_a22oi_1 _19602_ (.Y(_06022_),
    .B1(_06021_),
    .B2(net6996),
    .A2(_05882_),
    .A1(net6937));
 sg13g2_a21oi_1 _19603_ (.A1(net7003),
    .A2(_06022_),
    .Y(_06023_),
    .B1(_06017_));
 sg13g2_xnor2_1 _19604_ (.Y(_06024_),
    .A(net7112),
    .B(_06023_));
 sg13g2_nand2b_1 _19605_ (.Y(_06025_),
    .B(net6890),
    .A_N(net6891));
 sg13g2_nor2b_1 _19606_ (.A(net6890),
    .B_N(net6891),
    .Y(_06026_));
 sg13g2_a21oi_1 _19607_ (.A1(_05579_),
    .A2(_06025_),
    .Y(_06027_),
    .B1(_06026_));
 sg13g2_nor2_1 _19608_ (.A(net7113),
    .B(_05882_),
    .Y(_06028_));
 sg13g2_o21ai_1 _19609_ (.B1(_06028_),
    .Y(_06029_),
    .A1(net7117),
    .A2(net6991));
 sg13g2_a21oi_1 _19610_ (.A1(_06015_),
    .A2(_06029_),
    .Y(_06030_),
    .B1(net6994));
 sg13g2_nor4_1 _19611_ (.A(net7057),
    .B(net6938),
    .C(net7113),
    .D(_05882_),
    .Y(_06031_));
 sg13g2_o21ai_1 _19612_ (.B1(net6999),
    .Y(_06032_),
    .A1(_06030_),
    .A2(_06031_));
 sg13g2_a21oi_1 _19613_ (.A1(net6994),
    .A2(net6938),
    .Y(_06033_),
    .B1(_05755_));
 sg13g2_a21oi_1 _19614_ (.A1(_05654_),
    .A2(_05887_),
    .Y(_06034_),
    .B1(_06033_));
 sg13g2_nand3_1 _19615_ (.B(_05183_),
    .C(_05881_),
    .A(net7119),
    .Y(_06035_));
 sg13g2_or4_1 _19616_ (.A(_04798_),
    .B(_04915_),
    .C(_05183_),
    .D(_05881_),
    .X(_06036_));
 sg13g2_a221oi_1 _19617_ (.B2(_06036_),
    .C1(_05754_),
    .B1(_06035_),
    .A1(net7119),
    .Y(_06037_),
    .A2(_05024_));
 sg13g2_nand2_1 _19618_ (.Y(_06038_),
    .A(_06012_),
    .B(_06015_));
 sg13g2_nor2_1 _19619_ (.A(net6999),
    .B(_05755_),
    .Y(_06039_));
 sg13g2_a221oi_1 _19620_ (.B2(_06039_),
    .C1(_06037_),
    .B1(_06038_),
    .A1(net7057),
    .Y(_06040_),
    .A2(_06014_));
 sg13g2_o21ai_1 _19621_ (.B1(_06032_),
    .Y(_06041_),
    .A1(_06034_),
    .A2(_06040_));
 sg13g2_xor2_1 _19622_ (.B(_06041_),
    .A(_06027_),
    .X(_06042_));
 sg13g2_xnor2_1 _19623_ (.Y(_06043_),
    .A(_06024_),
    .B(_06042_));
 sg13g2_mux2_1 _19624_ (.A0(net7113),
    .A1(_06020_),
    .S(net6945),
    .X(_06044_));
 sg13g2_o21ai_1 _19625_ (.B1(_06018_),
    .Y(_06045_),
    .A1(net7057),
    .A2(_06044_));
 sg13g2_mux2_1 _19626_ (.A0(_06016_),
    .A1(_06045_),
    .S(net7003),
    .X(_06046_));
 sg13g2_xnor2_1 _19627_ (.Y(_06047_),
    .A(_06011_),
    .B(_06046_));
 sg13g2_a21oi_1 _19628_ (.A1(_06012_),
    .A2(_06015_),
    .Y(_06048_),
    .B1(net6999));
 sg13g2_a221oi_1 _19629_ (.B2(net7113),
    .C1(_06037_),
    .B1(_06048_),
    .A1(net7057),
    .Y(_06049_),
    .A2(_06014_));
 sg13g2_a21oi_1 _19630_ (.A1(net6991),
    .A2(_05755_),
    .Y(_06050_),
    .B1(_05653_));
 sg13g2_nor2_1 _19631_ (.A(_06033_),
    .B(_06050_),
    .Y(_06051_));
 sg13g2_o21ai_1 _19632_ (.B1(_06032_),
    .Y(_06052_),
    .A1(_06049_),
    .A2(_06051_));
 sg13g2_nor2_1 _19633_ (.A(net6827),
    .B(_06052_),
    .Y(_06053_));
 sg13g2_nand2_1 _19634_ (.Y(_06054_),
    .A(net6827),
    .B(_06052_));
 sg13g2_xnor2_1 _19635_ (.Y(_06055_),
    .A(net6827),
    .B(_06052_));
 sg13g2_xnor2_1 _19636_ (.Y(_06056_),
    .A(_06047_),
    .B(_06055_));
 sg13g2_o21ai_1 _19637_ (.B1(_06043_),
    .Y(_06057_),
    .A1(_06008_),
    .A2(_06009_));
 sg13g2_or3_1 _19638_ (.A(_06008_),
    .B(_06009_),
    .C(_06043_),
    .X(_06058_));
 sg13g2_a21o_1 _19639_ (.A2(_05959_),
    .A1(_05877_),
    .B1(_05879_),
    .X(_06059_));
 sg13g2_o21ai_1 _19640_ (.B1(_06059_),
    .Y(_06060_),
    .A1(_05877_),
    .A2(_05959_));
 sg13g2_a21oi_1 _19641_ (.A1(_06057_),
    .A2(_06058_),
    .Y(_06061_),
    .B1(_06060_));
 sg13g2_nand3_1 _19642_ (.B(_06058_),
    .C(_06060_),
    .A(_06057_),
    .Y(_06062_));
 sg13g2_nand2b_1 _19643_ (.Y(_06063_),
    .B(_06062_),
    .A_N(_06061_));
 sg13g2_xor2_1 _19644_ (.B(_06063_),
    .A(_05963_),
    .X(_06064_));
 sg13g2_xnor2_1 _19645_ (.Y(_06065_),
    .A(net6894),
    .B(_06001_));
 sg13g2_nor2_1 _19646_ (.A(_06005_),
    .B(_06065_),
    .Y(_06066_));
 sg13g2_inv_1 _19647_ (.Y(_06067_),
    .A(_00275_));
 sg13g2_xnor2_1 _19648_ (.Y(_06068_),
    .A(net6893),
    .B(_06056_));
 sg13g2_a21oi_1 _19649_ (.A1(_06005_),
    .A2(_06065_),
    .Y(_06069_),
    .B1(_06068_));
 sg13g2_nor2_1 _19650_ (.A(_06066_),
    .B(_06069_),
    .Y(_06070_));
 sg13g2_nor3_1 _19651_ (.A(net7145),
    .B(net7132),
    .C(net7118),
    .Y(_06071_));
 sg13g2_nand2b_1 _19652_ (.Y(_06072_),
    .B(net7145),
    .A_N(net7154));
 sg13g2_xnor2_1 _19653_ (.Y(_06073_),
    .A(net7154),
    .B(net7145));
 sg13g2_nand3b_1 _19654_ (.B(net7133),
    .C(net7154),
    .Y(_06074_),
    .A_N(net7145));
 sg13g2_o21ai_1 _19655_ (.B1(_06074_),
    .Y(_06075_),
    .A1(net7115),
    .A2(_06072_));
 sg13g2_a221oi_1 _19656_ (.B2(net7164),
    .C1(_06071_),
    .B1(_06075_),
    .A1(_05967_),
    .Y(_06076_),
    .A2(_06073_));
 sg13g2_inv_1 _19657_ (.Y(_06077_),
    .A(_00007_));
 sg13g2_nor2_1 _19658_ (.A(net7141),
    .B(net7136),
    .Y(_06078_));
 sg13g2_nor2_1 _19659_ (.A(net7150),
    .B(net7134),
    .Y(_06079_));
 sg13g2_xnor2_1 _19660_ (.Y(_06080_),
    .A(_06078_),
    .B(_06079_));
 sg13g2_and2_1 _19661_ (.A(net7157),
    .B(net7063),
    .X(_06081_));
 sg13g2_xor2_1 _19662_ (.B(_06081_),
    .A(_06080_),
    .X(_06082_));
 sg13g2_xnor2_1 _19663_ (.Y(_06083_),
    .A(_06080_),
    .B(_06081_));
 sg13g2_and2_1 _19664_ (.A(_05973_),
    .B(_05974_),
    .X(_06084_));
 sg13g2_or2_1 _19665_ (.X(_06085_),
    .B(_05974_),
    .A(_05973_));
 sg13g2_a21o_1 _19666_ (.A2(_06085_),
    .A1(_05975_),
    .B1(_06084_),
    .X(_06086_));
 sg13g2_o21ai_1 _19667_ (.B1(_06085_),
    .Y(_06087_),
    .A1(_05976_),
    .A2(_06084_));
 sg13g2_nand2_1 _19668_ (.Y(_06088_),
    .A(_06083_),
    .B(_06086_));
 sg13g2_xnor2_1 _19669_ (.Y(_06089_),
    .A(_06083_),
    .B(_06086_));
 sg13g2_xnor2_1 _19670_ (.Y(_06090_),
    .A(_06076_),
    .B(_06089_));
 sg13g2_a21oi_1 _19671_ (.A1(_05972_),
    .A2(_05978_),
    .Y(_06091_),
    .B1(_05969_));
 sg13g2_nor2_1 _19672_ (.A(_05965_),
    .B(_05966_),
    .Y(_06092_));
 sg13g2_a21oi_1 _19673_ (.A1(_05965_),
    .A2(_05966_),
    .Y(_06093_),
    .B1(_05967_));
 sg13g2_nor2_1 _19674_ (.A(_06092_),
    .B(_06093_),
    .Y(_06094_));
 sg13g2_xnor2_1 _19675_ (.Y(_06095_),
    .A(_05923_),
    .B(_06094_));
 sg13g2_nor3_1 _19676_ (.A(_05979_),
    .B(_06091_),
    .C(_06095_),
    .Y(_06096_));
 sg13g2_o21ai_1 _19677_ (.B1(_06095_),
    .Y(_06097_),
    .A1(_05979_),
    .A2(_06091_));
 sg13g2_nor2b_1 _19678_ (.A(_06096_),
    .B_N(_06097_),
    .Y(_06098_));
 sg13g2_xnor2_1 _19679_ (.Y(_06099_),
    .A(_06090_),
    .B(_06098_));
 sg13g2_a22oi_1 _19680_ (.Y(_06100_),
    .B1(_05993_),
    .B2(_05991_),
    .A2(_05992_),
    .A1(_05981_));
 sg13g2_nand3_1 _19681_ (.B(_05983_),
    .C(_05984_),
    .A(_05789_),
    .Y(_06101_));
 sg13g2_a22oi_1 _19682_ (.Y(_06102_),
    .B1(_06101_),
    .B2(net7067),
    .A2(_05985_),
    .A1(_05920_));
 sg13g2_nand2b_1 _19683_ (.Y(_06103_),
    .B(net7118),
    .A_N(_06102_));
 sg13g2_xnor2_1 _19684_ (.Y(_06104_),
    .A(_06100_),
    .B(_06103_));
 sg13g2_xor2_1 _19685_ (.B(_06104_),
    .A(_06099_),
    .X(_06105_));
 sg13g2_xnor2_1 _19686_ (.Y(_06106_),
    .A(_06099_),
    .B(_06104_));
 sg13g2_nand3_1 _19687_ (.B(_05996_),
    .C(_05999_),
    .A(_05964_),
    .Y(_06107_));
 sg13g2_nand3b_1 _19688_ (.B(net6828),
    .C(_05999_),
    .Y(_06108_),
    .A_N(_05964_));
 sg13g2_nand3_1 _19689_ (.B(_05964_),
    .C(net6828),
    .A(net6860),
    .Y(_06109_));
 sg13g2_nand3b_1 _19690_ (.B(_05996_),
    .C(net6894),
    .Y(_06110_),
    .A_N(_05964_));
 sg13g2_nand4_1 _19691_ (.B(_06108_),
    .C(_06109_),
    .A(_06107_),
    .Y(_06111_),
    .D(_06110_));
 sg13g2_xnor2_1 _19692_ (.Y(_06112_),
    .A(_06105_),
    .B(_06111_));
 sg13g2_nand4_1 _19693_ (.B(net6937),
    .C(_06010_),
    .A(net6996),
    .Y(_06113_),
    .D(_06028_));
 sg13g2_xnor2_1 _19694_ (.Y(_06114_),
    .A(_05024_),
    .B(_05182_));
 sg13g2_nand4_1 _19695_ (.B(_05881_),
    .C(_06011_),
    .A(net7119),
    .Y(_06115_),
    .D(_06114_));
 sg13g2_nand3_1 _19696_ (.B(_06010_),
    .C(_06020_),
    .A(net6944),
    .Y(_06116_));
 sg13g2_o21ai_1 _19697_ (.B1(_05579_),
    .Y(_06117_),
    .A1(net6891),
    .A2(_05999_));
 sg13g2_nand2_1 _19698_ (.Y(_06118_),
    .A(net6891),
    .B(_05999_));
 sg13g2_nand2_1 _19699_ (.Y(_06119_),
    .A(_06117_),
    .B(_06118_));
 sg13g2_a21oi_1 _19700_ (.A1(_01663_),
    .A2(net7322),
    .Y(_06120_),
    .B1(net7317));
 sg13g2_a21o_1 _19701_ (.A2(net7321),
    .A1(_01663_),
    .B1(net7317),
    .X(_06121_));
 sg13g2_a21oi_1 _19702_ (.A1(net6937),
    .A2(net7112),
    .Y(_06122_),
    .B1(_05287_));
 sg13g2_nand2_1 _19703_ (.Y(_06123_),
    .A(net6937),
    .B(_06011_));
 sg13g2_nand3_1 _19704_ (.B(_05881_),
    .C(_06123_),
    .A(net7001),
    .Y(_06124_));
 sg13g2_nand3_1 _19705_ (.B(net6944),
    .C(_06011_),
    .A(net7055),
    .Y(_06125_));
 sg13g2_nand3_1 _19706_ (.B(_05882_),
    .C(_06010_),
    .A(_05644_),
    .Y(_06126_));
 sg13g2_nand3_1 _19707_ (.B(_06125_),
    .C(_06126_),
    .A(net6998),
    .Y(_06127_));
 sg13g2_nand3_1 _19708_ (.B(_06115_),
    .C(_06116_),
    .A(_06113_),
    .Y(_06128_));
 sg13g2_o21ai_1 _19709_ (.B1(_06127_),
    .Y(_06129_),
    .A1(net6998),
    .A2(_06128_));
 sg13g2_a21oi_1 _19710_ (.A1(net6944),
    .A2(net7112),
    .Y(_06130_),
    .B1(net7055));
 sg13g2_a22oi_1 _19711_ (.Y(_06131_),
    .B1(_06124_),
    .B2(_06130_),
    .A2(_06122_),
    .A1(net7055));
 sg13g2_xnor2_1 _19712_ (.Y(_06132_),
    .A(net7111),
    .B(_06131_));
 sg13g2_xnor2_1 _19713_ (.Y(_06133_),
    .A(_06129_),
    .B(_06132_));
 sg13g2_xnor2_1 _19714_ (.Y(_06134_),
    .A(_06119_),
    .B(_06133_));
 sg13g2_inv_1 _19715_ (.Y(_06135_),
    .A(_00248_));
 sg13g2_xnor2_1 _19716_ (.Y(_06136_),
    .A(_06112_),
    .B(_06134_));
 sg13g2_xnor2_1 _19717_ (.Y(_06137_),
    .A(net6892),
    .B(_06047_));
 sg13g2_o21ai_1 _19718_ (.B1(_06054_),
    .Y(_06138_),
    .A1(_06053_),
    .A2(_06137_));
 sg13g2_xor2_1 _19719_ (.B(_06138_),
    .A(_06136_),
    .X(_06139_));
 sg13g2_inv_1 _19720_ (.Y(_06140_),
    .A(_00246_));
 sg13g2_xnor2_1 _19721_ (.Y(_06141_),
    .A(_06070_),
    .B(_06139_));
 sg13g2_nor2_1 _19722_ (.A(net6894),
    .B(_05999_),
    .Y(_06142_));
 sg13g2_o21ai_1 _19723_ (.B1(_06142_),
    .Y(_06143_),
    .A1(_06105_),
    .A2(net6714));
 sg13g2_and2_1 _19724_ (.A(net6894),
    .B(_05999_),
    .X(_06144_));
 sg13g2_inv_1 _19725_ (.Y(_06145_),
    .A(_00001_));
 sg13g2_o21ai_1 _19726_ (.B1(_06144_),
    .Y(_06146_),
    .A1(_06106_),
    .A2(net6714));
 sg13g2_a22oi_1 _19727_ (.Y(_06147_),
    .B1(_06143_),
    .B2(_06146_),
    .A2(net6828),
    .A1(_05964_));
 sg13g2_nor2_1 _19728_ (.A(_05964_),
    .B(net6828),
    .Y(_06148_));
 sg13g2_inv_1 _19729_ (.Y(_06149_),
    .A(_00000_));
 sg13g2_xnor2_1 _19730_ (.Y(_06150_),
    .A(net6860),
    .B(_06105_));
 sg13g2_o21ai_1 _19731_ (.B1(_06150_),
    .Y(_06151_),
    .A1(net6714),
    .A2(_06148_));
 sg13g2_inv_1 _19732_ (.Y(_06152_),
    .A(_00243_));
 sg13g2_nand2_1 _19733_ (.Y(_06153_),
    .A(net6714),
    .B(_06148_));
 sg13g2_nand2_1 _19734_ (.Y(_06154_),
    .A(_06151_),
    .B(_06153_));
 sg13g2_nor2_1 _19735_ (.A(_06147_),
    .B(_06154_),
    .Y(_06155_));
 sg13g2_inv_1 _19736_ (.Y(_06156_),
    .A(_06157_));
 sg13g2_o21ai_1 _19737_ (.B1(_06119_),
    .Y(_06157_),
    .A1(_06129_),
    .A2(_06132_));
 sg13g2_a21oi_1 _19738_ (.A1(_06129_),
    .A2(_06132_),
    .Y(_06158_),
    .B1(_06156_));
 sg13g2_inv_1 _19739_ (.Y(_06159_),
    .A(_06158_));
 sg13g2_a21oi_1 _19740_ (.A1(_01664_),
    .A2(net7321),
    .Y(_06160_),
    .B1(net7316));
 sg13g2_a21o_1 _19741_ (.A2(net7321),
    .A1(_01664_),
    .B1(net7316),
    .X(_06161_));
 sg13g2_inv_1 _19742_ (.Y(_06162_),
    .A(_00242_));
 sg13g2_nor4_1 _19743_ (.A(net7117),
    .B(net6991),
    .C(_06010_),
    .D(_06120_),
    .Y(_06163_));
 sg13g2_a21oi_1 _19744_ (.A1(net6937),
    .A2(net7112),
    .Y(_06164_),
    .B1(_06163_));
 sg13g2_a221oi_1 _19745_ (.B2(net6996),
    .C1(net6998),
    .B1(_06164_),
    .A1(net6937),
    .Y(_06165_),
    .A2(net7111));
 sg13g2_o21ai_1 _19746_ (.B1(_06120_),
    .Y(_06166_),
    .A1(net7117),
    .A2(net6991));
 sg13g2_nand3_1 _19747_ (.B(_05183_),
    .C(_06121_),
    .A(net7119),
    .Y(_06167_));
 sg13g2_inv_1 _19748_ (.Y(_06168_),
    .A(_00241_));
 sg13g2_mux2_1 _19749_ (.A0(_06166_),
    .A1(_06167_),
    .S(net6995),
    .X(_06169_));
 sg13g2_a21oi_1 _19750_ (.A1(net6998),
    .A2(_06169_),
    .Y(_06170_),
    .B1(_06165_));
 sg13g2_xnor2_1 _19751_ (.Y(_06171_),
    .A(net7110),
    .B(_06170_));
 sg13g2_o21ai_1 _19752_ (.B1(_06167_),
    .Y(_06172_),
    .A1(_05881_),
    .A2(_06166_));
 sg13g2_nor2_1 _19753_ (.A(net7055),
    .B(_06011_),
    .Y(_06173_));
 sg13g2_inv_1 _19754_ (.Y(_06174_),
    .A(_00240_));
 sg13g2_nor2_1 _19755_ (.A(net7112),
    .B(net7111),
    .Y(_06175_));
 sg13g2_a22oi_1 _19756_ (.Y(_06176_),
    .B1(_06175_),
    .B2(_06014_),
    .A2(_06173_),
    .A1(_06172_));
 sg13g2_o21ai_1 _19757_ (.B1(_06175_),
    .Y(_06177_),
    .A1(net7117),
    .A2(net6991));
 sg13g2_nand2_1 _19758_ (.Y(_06178_),
    .A(_06167_),
    .B(_06177_));
 sg13g2_a22oi_1 _19759_ (.Y(_06179_),
    .B1(_06178_),
    .B2(net7055),
    .A2(_06175_),
    .A1(_05418_));
 sg13g2_mux2_1 _19760_ (.A0(_06176_),
    .A1(_06179_),
    .S(net6998),
    .X(_06180_));
 sg13g2_nor3_1 _19761_ (.A(net7114),
    .B(net6891),
    .C(_06102_),
    .Y(_06181_));
 sg13g2_o21ai_1 _19762_ (.B1(net6891),
    .Y(_06182_),
    .A1(net7114),
    .A2(_06102_));
 sg13g2_o21ai_1 _19763_ (.B1(_06182_),
    .Y(_06183_),
    .A1(net6895),
    .A2(_06181_));
 sg13g2_xnor2_1 _19764_ (.Y(_06184_),
    .A(_06180_),
    .B(_06183_));
 sg13g2_inv_1 _19765_ (.Y(_06185_),
    .A(_00238_));
 sg13g2_xnor2_1 _19766_ (.Y(_06186_),
    .A(_06171_),
    .B(_06184_));
 sg13g2_nor2_1 _19767_ (.A(_06099_),
    .B(_06100_),
    .Y(_06187_));
 sg13g2_xnor2_1 _19768_ (.Y(_06188_),
    .A(net6860),
    .B(_06103_));
 sg13g2_a21oi_1 _19769_ (.A1(_06099_),
    .A2(_06100_),
    .Y(_06189_),
    .B1(_06188_));
 sg13g2_or2_1 _19770_ (.X(_06190_),
    .B(_06189_),
    .A(_06187_));
 sg13g2_a21oi_1 _19771_ (.A1(_06090_),
    .A2(_06097_),
    .Y(_06191_),
    .B1(_06096_));
 sg13g2_nor2_1 _19772_ (.A(net7142),
    .B(net7130),
    .Y(_06192_));
 sg13g2_nor2_1 _19773_ (.A(net7136),
    .B(net7134),
    .Y(_06193_));
 sg13g2_nand3_1 _19774_ (.B(net7149),
    .C(net7129),
    .A(net7637),
    .Y(_06194_));
 sg13g2_inv_1 _19775_ (.Y(_06195_),
    .A(_00235_));
 sg13g2_xnor2_1 _19776_ (.Y(_06196_),
    .A(_06193_),
    .B(_06194_));
 sg13g2_xnor2_1 _19777_ (.Y(_06197_),
    .A(_06192_),
    .B(_06196_));
 sg13g2_nor2_1 _19778_ (.A(_06078_),
    .B(_06079_),
    .Y(_06198_));
 sg13g2_inv_1 _19779_ (.Y(_06199_),
    .A(_00234_));
 sg13g2_a22oi_1 _19780_ (.Y(_06200_),
    .B1(_06078_),
    .B2(_06079_),
    .A2(net7063),
    .A1(net7157));
 sg13g2_or2_1 _19781_ (.X(_06201_),
    .B(_06200_),
    .A(_06198_));
 sg13g2_nand2_1 _19782_ (.Y(_06202_),
    .A(_06197_),
    .B(_06201_));
 sg13g2_nor2_1 _19783_ (.A(_06197_),
    .B(_06201_),
    .Y(_06203_));
 sg13g2_xor2_1 _19784_ (.B(_06201_),
    .A(_06197_),
    .X(_06204_));
 sg13g2_a21oi_1 _19785_ (.A1(_06072_),
    .A2(_06074_),
    .Y(_06205_),
    .B1(net7164));
 sg13g2_a21o_1 _19786_ (.A2(_06073_),
    .A1(net7164),
    .B1(_06205_),
    .X(_06206_));
 sg13g2_nor2_1 _19787_ (.A(net7120),
    .B(_06206_),
    .Y(_06207_));
 sg13g2_inv_1 _19788_ (.Y(_06208_),
    .A(_00232_));
 sg13g2_xnor2_1 _19789_ (.Y(_06209_),
    .A(_06204_),
    .B(_06207_));
 sg13g2_inv_1 _19790_ (.Y(_06210_),
    .A(_00231_));
 sg13g2_nor3_1 _19791_ (.A(net7164),
    .B(net7145),
    .C(net7131),
    .Y(_06211_));
 sg13g2_a21oi_1 _19792_ (.A1(net7164),
    .A2(net7145),
    .Y(_06212_),
    .B1(net7154));
 sg13g2_or2_1 _19793_ (.X(_06213_),
    .B(_06212_),
    .A(_06211_));
 sg13g2_nand2_1 _19794_ (.Y(_06214_),
    .A(net7118),
    .B(_06213_));
 sg13g2_xor2_1 _19795_ (.B(_06214_),
    .A(net6989),
    .X(_06215_));
 sg13g2_a21o_1 _19796_ (.A2(_06087_),
    .A1(_06082_),
    .B1(_06076_),
    .X(_06216_));
 sg13g2_nand2_1 _19797_ (.Y(_06217_),
    .A(_06088_),
    .B(_06216_));
 sg13g2_and3_1 _19798_ (.X(_06218_),
    .A(_06088_),
    .B(_06215_),
    .C(_06216_));
 sg13g2_inv_1 _19799_ (.Y(_06219_),
    .A(_00228_));
 sg13g2_xnor2_1 _19800_ (.Y(_06220_),
    .A(_06209_),
    .B(_06217_));
 sg13g2_xnor2_1 _19801_ (.Y(_06221_),
    .A(_06215_),
    .B(_06220_));
 sg13g2_o21ai_1 _19802_ (.B1(net7067),
    .Y(_06222_),
    .A1(_05788_),
    .A2(_06094_));
 sg13g2_nand2_1 _19803_ (.Y(_06223_),
    .A(_05920_),
    .B(_06094_));
 sg13g2_inv_1 _19804_ (.Y(_06224_),
    .A(_00226_));
 sg13g2_a21oi_1 _19805_ (.A1(_06222_),
    .A2(_06223_),
    .Y(_06225_),
    .B1(net7114));
 sg13g2_xnor2_1 _19806_ (.Y(_06226_),
    .A(_06191_),
    .B(_06225_));
 sg13g2_inv_1 _19807_ (.Y(_06227_),
    .A(_00225_));
 sg13g2_xnor2_1 _19808_ (.Y(_06228_),
    .A(_06221_),
    .B(_06226_));
 sg13g2_xnor2_1 _19809_ (.Y(_06229_),
    .A(_05727_),
    .B(_06228_));
 sg13g2_xnor2_1 _19810_ (.Y(_06230_),
    .A(_06190_),
    .B(_06229_));
 sg13g2_inv_1 _19811_ (.Y(_06231_),
    .A(_00224_));
 sg13g2_xnor2_1 _19812_ (.Y(_06232_),
    .A(_06186_),
    .B(_06230_));
 sg13g2_xnor2_1 _19813_ (.Y(_06233_),
    .A(_06159_),
    .B(_06232_));
 sg13g2_xnor2_1 _19814_ (.Y(_06234_),
    .A(_06155_),
    .B(_06233_));
 sg13g2_inv_1 _19815_ (.Y(_06235_),
    .A(_00223_));
 sg13g2_inv_1 _19816_ (.Y(_06236_),
    .A(_00222_));
 sg13g2_xnor2_1 _19817_ (.Y(_06237_),
    .A(_05724_),
    .B(_06228_));
 sg13g2_nand2_1 _19818_ (.Y(_06238_),
    .A(_06190_),
    .B(_06237_));
 sg13g2_inv_1 _19819_ (.Y(_06239_),
    .A(_00221_));
 sg13g2_inv_1 _19820_ (.Y(_06240_),
    .A(_00220_));
 sg13g2_inv_1 _19821_ (.Y(_06241_),
    .A(_00219_));
 sg13g2_inv_1 _19822_ (.Y(_06242_),
    .A(_00216_));
 sg13g2_mux2_1 _19823_ (.A0(_06166_),
    .A1(_06167_),
    .S(net6995),
    .X(_06243_));
 sg13g2_o21ai_1 _19824_ (.B1(net6944),
    .Y(_06244_),
    .A1(_06010_),
    .A2(_06120_));
 sg13g2_nand2_1 _19825_ (.Y(_06245_),
    .A(_06123_),
    .B(_06244_));
 sg13g2_a221oi_1 _19826_ (.B2(net6995),
    .C1(net6998),
    .B1(_06245_),
    .A1(net6937),
    .Y(_06246_),
    .A2(net7111));
 sg13g2_inv_1 _19827_ (.Y(_06247_),
    .A(_00214_));
 sg13g2_a21oi_1 _19828_ (.A1(net6998),
    .A2(_06243_),
    .Y(_06248_),
    .B1(_06246_));
 sg13g2_xnor2_1 _19829_ (.Y(_06249_),
    .A(net7110),
    .B(_06248_));
 sg13g2_mux2_1 _19830_ (.A0(_06176_),
    .A1(_06179_),
    .S(net6998),
    .X(_06250_));
 sg13g2_xor2_1 _19831_ (.B(_06186_),
    .A(net6893),
    .X(_06251_));
 sg13g2_o21ai_1 _19832_ (.B1(_06251_),
    .Y(_06252_),
    .A1(_06190_),
    .A2(_06237_));
 sg13g2_nand2_1 _19833_ (.Y(_06253_),
    .A(_06238_),
    .B(_06252_));
 sg13g2_o21ai_1 _19834_ (.B1(_04737_),
    .Y(_06254_),
    .A1(net7150),
    .A2(net7136));
 sg13g2_inv_1 _19835_ (.Y(_06255_),
    .A(_00211_));
 sg13g2_and2_1 _19836_ (.A(net7136),
    .B(net7063),
    .X(_06256_));
 sg13g2_nand2_1 _19837_ (.Y(_06257_),
    .A(net7136),
    .B(net7063));
 sg13g2_nand3b_1 _19838_ (.B(_06254_),
    .C(net7133),
    .Y(_06258_),
    .A_N(_06078_));
 sg13g2_nand3_1 _19839_ (.B(net7136),
    .C(_06192_),
    .A(net7150),
    .Y(_06259_));
 sg13g2_nand2b_1 _19840_ (.Y(_06260_),
    .B(net7130),
    .A_N(_06194_));
 sg13g2_nand2_1 _19841_ (.Y(_06261_),
    .A(net7132),
    .B(net7063));
 sg13g2_nand3_1 _19842_ (.B(_06259_),
    .C(_06260_),
    .A(_06258_),
    .Y(_06262_));
 sg13g2_inv_1 _19843_ (.Y(_06263_),
    .A(_00209_));
 sg13g2_a22oi_1 _19844_ (.Y(_06264_),
    .B1(_06262_),
    .B2(_04650_),
    .A2(_06256_),
    .A1(net7130));
 sg13g2_xnor2_1 _19845_ (.Y(_06265_),
    .A(net7142),
    .B(_06206_));
 sg13g2_inv_1 _19846_ (.Y(_06266_),
    .A(_00208_));
 sg13g2_nor2_1 _19847_ (.A(net7114),
    .B(_06265_),
    .Y(_06267_));
 sg13g2_xnor2_1 _19848_ (.Y(_06268_),
    .A(_06264_),
    .B(_06267_));
 sg13g2_a21o_1 _19849_ (.A2(_06207_),
    .A1(_06202_),
    .B1(_06203_),
    .X(_06269_));
 sg13g2_xnor2_1 _19850_ (.Y(_06270_),
    .A(_06215_),
    .B(_06269_));
 sg13g2_xnor2_1 _19851_ (.Y(_06271_),
    .A(_06268_),
    .B(_06270_));
 sg13g2_a21o_1 _19852_ (.A2(_06216_),
    .A1(_06088_),
    .B1(_06215_),
    .X(_06272_));
 sg13g2_a21oi_1 _19853_ (.A1(_06209_),
    .A2(_06272_),
    .Y(_06273_),
    .B1(_06218_));
 sg13g2_o21ai_1 _19854_ (.B1(net7067),
    .Y(_06274_),
    .A1(_05788_),
    .A2(_06213_));
 sg13g2_nand2_1 _19855_ (.Y(_06275_),
    .A(_05920_),
    .B(_06213_));
 sg13g2_a21o_1 _19856_ (.A2(_06275_),
    .A1(_06274_),
    .B1(net7114),
    .X(_06276_));
 sg13g2_inv_1 _19857_ (.Y(_06277_),
    .A(_06278_));
 sg13g2_xnor2_1 _19858_ (.Y(_06278_),
    .A(_05724_),
    .B(_06276_));
 sg13g2_nor2_1 _19859_ (.A(_06273_),
    .B(_06278_),
    .Y(_06279_));
 sg13g2_inv_1 _19860_ (.Y(_06280_),
    .A(_00203_));
 sg13g2_nand2_1 _19861_ (.Y(_06281_),
    .A(_06273_),
    .B(_06278_));
 sg13g2_xor2_1 _19862_ (.B(_06278_),
    .A(_06273_),
    .X(_06282_));
 sg13g2_xnor2_1 _19863_ (.Y(_06283_),
    .A(_06271_),
    .B(_06282_));
 sg13g2_xnor2_1 _19864_ (.Y(_06284_),
    .A(net6894),
    .B(_06225_));
 sg13g2_a21oi_1 _19865_ (.A1(_06191_),
    .A2(_06221_),
    .Y(_06285_),
    .B1(_06284_));
 sg13g2_nor2_1 _19866_ (.A(_06191_),
    .B(_06221_),
    .Y(_06286_));
 sg13g2_or2_1 _19867_ (.X(_06287_),
    .B(_06286_),
    .A(_06285_));
 sg13g2_nor2_1 _19868_ (.A(net6935),
    .B(_06161_),
    .Y(_06288_));
 sg13g2_nor2_1 _19869_ (.A(net7110),
    .B(_06166_),
    .Y(_06289_));
 sg13g2_o21ai_1 _19870_ (.B1(net7055),
    .Y(_06290_),
    .A1(_06288_),
    .A2(_06289_));
 sg13g2_nand2_1 _19871_ (.Y(_06291_),
    .A(net6941),
    .B(_06161_));
 sg13g2_nor2_1 _19872_ (.A(net6941),
    .B(_06161_),
    .Y(_06292_));
 sg13g2_nand2_1 _19873_ (.Y(_06293_),
    .A(_06011_),
    .B(_06292_));
 sg13g2_nand2_1 _19874_ (.Y(_06294_),
    .A(_06291_),
    .B(_06293_));
 sg13g2_nand3_1 _19875_ (.B(_06120_),
    .C(_06294_),
    .A(net6995),
    .Y(_06295_));
 sg13g2_nand4_1 _19876_ (.B(_06011_),
    .C(net7111),
    .A(net6944),
    .Y(_06296_),
    .D(net7110));
 sg13g2_nand4_1 _19877_ (.B(_06290_),
    .C(_06295_),
    .A(net7001),
    .Y(_06297_),
    .D(_06296_));
 sg13g2_nand3_1 _19878_ (.B(net7111),
    .C(net7110),
    .A(net6935),
    .Y(_06298_));
 sg13g2_a21oi_1 _19879_ (.A1(_06291_),
    .A2(_06298_),
    .Y(_06299_),
    .B1(net6995));
 sg13g2_nand3_1 _19880_ (.B(net7111),
    .C(net7110),
    .A(net6897),
    .Y(_06300_));
 sg13g2_nand2b_1 _19881_ (.Y(_06301_),
    .B(_06300_),
    .A_N(_06299_));
 sg13g2_o21ai_1 _19882_ (.B1(_06297_),
    .Y(_06302_),
    .A1(net7001),
    .A2(_06301_));
 sg13g2_a21o_1 _19883_ (.A2(_06225_),
    .A1(_05834_),
    .B1(net6895),
    .X(_06303_));
 sg13g2_o21ai_1 _19884_ (.B1(_06303_),
    .Y(_06304_),
    .A1(_05834_),
    .A2(_06225_));
 sg13g2_a21oi_1 _19885_ (.A1(_01665_),
    .A2(net7321),
    .Y(_06305_),
    .B1(net7316));
 sg13g2_a21o_1 _19886_ (.A2(net7321),
    .A1(_01665_),
    .B1(net7316),
    .X(_06306_));
 sg13g2_nor2_1 _19887_ (.A(net6941),
    .B(net7110),
    .Y(_06307_));
 sg13g2_nor3_1 _19888_ (.A(net6997),
    .B(net7111),
    .C(_06307_),
    .Y(_06308_));
 sg13g2_a21oi_1 _19889_ (.A1(net6944),
    .A2(net7110),
    .Y(_06309_),
    .B1(_06308_));
 sg13g2_nor3_1 _19890_ (.A(net6995),
    .B(_05287_),
    .C(_06292_),
    .Y(_06310_));
 sg13g2_a21oi_1 _19891_ (.A1(net6995),
    .A2(_06309_),
    .Y(_06311_),
    .B1(_06310_));
 sg13g2_xor2_1 _19892_ (.B(_06304_),
    .A(_06283_),
    .X(_06312_));
 sg13g2_xnor2_1 _19893_ (.Y(_06313_),
    .A(_06302_),
    .B(_06312_));
 sg13g2_xnor2_1 _19894_ (.Y(_06314_),
    .A(_06305_),
    .B(_06311_));
 sg13g2_xor2_1 _19895_ (.B(_06314_),
    .A(_06287_),
    .X(_06315_));
 sg13g2_xnor2_1 _19896_ (.Y(_06316_),
    .A(_06313_),
    .B(_06315_));
 sg13g2_nand2_1 _19897_ (.Y(_06317_),
    .A(_06183_),
    .B(_06250_));
 sg13g2_nor2_1 _19898_ (.A(_06183_),
    .B(_06250_),
    .Y(_06318_));
 sg13g2_xnor2_1 _19899_ (.Y(_06319_),
    .A(net6892),
    .B(_06249_));
 sg13g2_o21ai_1 _19900_ (.B1(_06317_),
    .Y(_06320_),
    .A1(_06318_),
    .A2(_06319_));
 sg13g2_xor2_1 _19901_ (.B(_06320_),
    .A(_06316_),
    .X(_06321_));
 sg13g2_xnor2_1 _19902_ (.Y(_06322_),
    .A(_06253_),
    .B(_06321_));
 sg13g2_nor2_1 _19903_ (.A(net7134),
    .B(net7130),
    .Y(_06323_));
 sg13g2_nor2_1 _19904_ (.A(net7142),
    .B(net7116),
    .Y(_06324_));
 sg13g2_xnor2_1 _19905_ (.Y(_06325_),
    .A(_06323_),
    .B(_06324_));
 sg13g2_xnor2_1 _19906_ (.Y(_06326_),
    .A(_06256_),
    .B(_06325_));
 sg13g2_nor2_1 _19907_ (.A(_06192_),
    .B(_06193_),
    .Y(_06327_));
 sg13g2_inv_1 _19908_ (.Y(_06328_),
    .A(_00189_));
 sg13g2_nand2_1 _19909_ (.Y(_06329_),
    .A(_06192_),
    .B(_06193_));
 sg13g2_o21ai_1 _19910_ (.B1(_06329_),
    .Y(_06330_),
    .A1(_06194_),
    .A2(_06327_));
 sg13g2_o21ai_1 _19911_ (.B1(_06330_),
    .Y(_06331_),
    .A1(_06207_),
    .A2(_06326_));
 sg13g2_nand2_1 _19912_ (.Y(_06332_),
    .A(_06207_),
    .B(_06326_));
 sg13g2_nand2_1 _19913_ (.Y(_06333_),
    .A(_06331_),
    .B(_06332_));
 sg13g2_xor2_1 _19914_ (.B(_06333_),
    .A(_06215_),
    .X(_06334_));
 sg13g2_a21oi_1 _19915_ (.A1(net7142),
    .A2(_06257_),
    .Y(_06335_),
    .B1(net7130));
 sg13g2_nor2_1 _19916_ (.A(net7114),
    .B(_06335_),
    .Y(_06336_));
 sg13g2_a21oi_1 _19917_ (.A1(net7114),
    .A2(_06256_),
    .Y(_06337_),
    .B1(_06336_));
 sg13g2_o21ai_1 _19918_ (.B1(_06261_),
    .Y(_06338_),
    .A1(net7134),
    .A2(_06337_));
 sg13g2_xor2_1 _19919_ (.B(_06338_),
    .A(_06267_),
    .X(_06339_));
 sg13g2_xnor2_1 _19920_ (.Y(_06340_),
    .A(_06334_),
    .B(_06339_));
 sg13g2_nor2_1 _19921_ (.A(_06268_),
    .B(_06269_),
    .Y(_06341_));
 sg13g2_nand2_1 _19922_ (.Y(_06342_),
    .A(_06268_),
    .B(_06269_));
 sg13g2_o21ai_1 _19923_ (.B1(_06342_),
    .Y(_06343_),
    .A1(_06215_),
    .A2(_06341_));
 sg13g2_xnor2_1 _19924_ (.Y(_06344_),
    .A(_06277_),
    .B(_06343_));
 sg13g2_inv_1 _19925_ (.Y(_06345_),
    .A(_00181_));
 sg13g2_xnor2_1 _19926_ (.Y(_06346_),
    .A(_06340_),
    .B(_06344_));
 sg13g2_a21oi_1 _19927_ (.A1(_06271_),
    .A2(_06281_),
    .Y(_06347_),
    .B1(_06279_));
 sg13g2_nor2_1 _19928_ (.A(net6935),
    .B(_06306_),
    .Y(_06348_));
 sg13g2_nor3_1 _19929_ (.A(net6942),
    .B(_06161_),
    .C(_06305_),
    .Y(_06349_));
 sg13g2_o21ai_1 _19930_ (.B1(net7054),
    .Y(_06350_),
    .A1(_06348_),
    .A2(_06349_));
 sg13g2_nor2_1 _19931_ (.A(_06160_),
    .B(_06306_),
    .Y(_06351_));
 sg13g2_nor2b_1 _19932_ (.A(_06167_),
    .B_N(_06351_),
    .Y(_06352_));
 sg13g2_nor3_1 _19933_ (.A(net6941),
    .B(_06120_),
    .C(_06306_),
    .Y(_06353_));
 sg13g2_a21oi_1 _19934_ (.A1(net6941),
    .A2(_06306_),
    .Y(_06354_),
    .B1(_06353_));
 sg13g2_nand2_1 _19935_ (.Y(_06355_),
    .A(net6995),
    .B(_06160_));
 sg13g2_mux2_1 _19936_ (.A0(_06306_),
    .A1(_06351_),
    .S(net6935),
    .X(_06356_));
 sg13g2_a22oi_1 _19937_ (.Y(_06357_),
    .B1(_06356_),
    .B2(net7054),
    .A2(_06351_),
    .A1(net6897));
 sg13g2_o21ai_1 _19938_ (.B1(_05579_),
    .Y(_06358_),
    .A1(_05835_),
    .A2(_06276_));
 sg13g2_nand2_1 _19939_ (.Y(_06359_),
    .A(_05835_),
    .B(_06276_));
 sg13g2_inv_1 _19940_ (.Y(_06360_),
    .A(_06361_));
 sg13g2_nand2_1 _19941_ (.Y(_06361_),
    .A(_06358_),
    .B(_06359_));
 sg13g2_inv_1 _19942_ (.Y(_06362_),
    .A(_00178_));
 sg13g2_a21oi_1 _19943_ (.A1(net7977),
    .A2(net7321),
    .Y(_06363_),
    .B1(net7316));
 sg13g2_a21o_1 _19944_ (.A2(net7321),
    .A1(net7977),
    .B1(net7316),
    .X(_06364_));
 sg13g2_nor2_1 _19945_ (.A(net6943),
    .B(_06305_),
    .Y(_06365_));
 sg13g2_nor3_1 _19946_ (.A(net6997),
    .B(_06161_),
    .C(_06365_),
    .Y(_06366_));
 sg13g2_nor3_1 _19947_ (.A(net7054),
    .B(_06348_),
    .C(_06366_),
    .Y(_06367_));
 sg13g2_a21oi_1 _19948_ (.A1(net6935),
    .A2(_06305_),
    .Y(_06368_),
    .B1(_05287_));
 sg13g2_inv_1 _19949_ (.Y(_06369_),
    .A(_00177_));
 sg13g2_a21oi_1 _19950_ (.A1(net7054),
    .A2(_06368_),
    .Y(_06370_),
    .B1(_06367_));
 sg13g2_o21ai_1 _19951_ (.B1(_06350_),
    .Y(_06371_),
    .A1(_06354_),
    .A2(_06355_));
 sg13g2_o21ai_1 _19952_ (.B1(net7001),
    .Y(_06372_),
    .A1(_06352_),
    .A2(_06371_));
 sg13g2_inv_1 _19953_ (.Y(_06373_),
    .A(_00175_));
 sg13g2_o21ai_1 _19954_ (.B1(_06372_),
    .Y(_06374_),
    .A1(net7001),
    .A2(_06357_));
 sg13g2_inv_1 _19955_ (.Y(_06375_),
    .A(_06376_));
 sg13g2_xnor2_1 _19956_ (.Y(_06376_),
    .A(_06363_),
    .B(_06370_));
 sg13g2_xnor2_1 _19957_ (.Y(_06377_),
    .A(_06360_),
    .B(_06376_));
 sg13g2_xnor2_1 _19958_ (.Y(_06378_),
    .A(_06374_),
    .B(_06377_));
 sg13g2_inv_1 _19959_ (.Y(_06379_),
    .A(_00174_));
 sg13g2_xor2_1 _19960_ (.B(_06347_),
    .A(_06346_),
    .X(_06380_));
 sg13g2_xnor2_1 _19961_ (.Y(_06381_),
    .A(_06378_),
    .B(_06380_));
 sg13g2_nand2b_1 _19962_ (.Y(_06382_),
    .B(_06287_),
    .A_N(_06283_));
 sg13g2_nand2b_1 _19963_ (.Y(_06383_),
    .B(_06283_),
    .A_N(_06287_));
 sg13g2_inv_1 _19964_ (.Y(_06384_),
    .A(_00173_));
 sg13g2_nor2_1 _19965_ (.A(_06302_),
    .B(_06304_),
    .Y(_06385_));
 sg13g2_inv_1 _19966_ (.Y(_06386_),
    .A(_00171_));
 sg13g2_inv_1 _19967_ (.Y(_06387_),
    .A(_00170_));
 sg13g2_inv_1 _19968_ (.Y(_06388_),
    .A(_00169_));
 sg13g2_nand2_1 _19969_ (.Y(_06389_),
    .A(_06302_),
    .B(_06304_));
 sg13g2_nor2_1 _19970_ (.A(_06382_),
    .B(_06389_),
    .Y(_06390_));
 sg13g2_inv_1 _19971_ (.Y(_06391_),
    .A(_00168_));
 sg13g2_nand2b_1 _19972_ (.Y(_06392_),
    .B(_06304_),
    .A_N(_06314_));
 sg13g2_nor2b_1 _19973_ (.A(_06392_),
    .B_N(_06302_),
    .Y(_06393_));
 sg13g2_inv_1 _19974_ (.Y(_06394_),
    .A(_00166_));
 sg13g2_mux2_1 _19975_ (.A0(_06385_),
    .A1(_06393_),
    .S(_06383_),
    .X(_06395_));
 sg13g2_nand2b_1 _19976_ (.Y(_06396_),
    .B(_06314_),
    .A_N(_06304_));
 sg13g2_nand2b_1 _19977_ (.Y(_06397_),
    .B(_06314_),
    .A_N(_06302_));
 sg13g2_a21oi_1 _19978_ (.A1(_06396_),
    .A2(_06397_),
    .Y(_06398_),
    .B1(_06383_));
 sg13g2_inv_1 _19979_ (.Y(_06399_),
    .A(_00165_));
 sg13g2_nor2_1 _19980_ (.A(_06395_),
    .B(_06398_),
    .Y(_06400_));
 sg13g2_nand2b_1 _19981_ (.Y(_06401_),
    .B(_06302_),
    .A_N(_06314_));
 sg13g2_nor2_1 _19982_ (.A(_06302_),
    .B(_06396_),
    .Y(_06402_));
 sg13g2_a21oi_1 _19983_ (.A1(_06382_),
    .A2(_06402_),
    .Y(_06403_),
    .B1(_06390_));
 sg13g2_a21o_1 _19984_ (.A2(_06401_),
    .A1(_06392_),
    .B1(_06382_),
    .X(_06404_));
 sg13g2_nand3_1 _19985_ (.B(_06403_),
    .C(_06404_),
    .A(_06400_),
    .Y(_06405_));
 sg13g2_inv_1 _19986_ (.Y(_06406_),
    .A(_00163_));
 sg13g2_xnor2_1 _19987_ (.Y(_06407_),
    .A(net6617),
    .B(_06405_));
 sg13g2_o21ai_1 _19988_ (.B1(_06374_),
    .Y(_06408_),
    .A1(_06360_),
    .A2(_06376_));
 sg13g2_o21ai_1 _19989_ (.B1(_06408_),
    .Y(_06409_),
    .A1(_06361_),
    .A2(_06375_));
 sg13g2_nor2_1 _19990_ (.A(_06305_),
    .B(_06364_),
    .Y(_06410_));
 sg13g2_nor2b_1 _19991_ (.A(_06291_),
    .B_N(_06410_),
    .Y(_06411_));
 sg13g2_nor3_1 _19992_ (.A(net6942),
    .B(_06306_),
    .C(net7109),
    .Y(_06412_));
 sg13g2_inv_1 _19993_ (.Y(_06413_),
    .A(_00162_));
 sg13g2_a21oi_1 _19994_ (.A1(net6941),
    .A2(net7109),
    .Y(_06414_),
    .B1(_06412_));
 sg13g2_nand2_1 _19995_ (.Y(_06415_),
    .A(net6942),
    .B(_06364_));
 sg13g2_nand2_1 _19996_ (.Y(_06416_),
    .A(_06307_),
    .B(net7109));
 sg13g2_a21oi_1 _19997_ (.A1(_06415_),
    .A2(_06416_),
    .Y(_06417_),
    .B1(_06306_));
 sg13g2_nor2_1 _19998_ (.A(net7054),
    .B(_06417_),
    .Y(_06418_));
 sg13g2_a21oi_1 _19999_ (.A1(net7054),
    .A2(_06414_),
    .Y(_06419_),
    .B1(_06418_));
 sg13g2_o21ai_1 _20000_ (.B1(net7000),
    .Y(_06420_),
    .A1(_06411_),
    .A2(_06419_));
 sg13g2_inv_1 _20001_ (.Y(_06421_),
    .A(_00161_));
 sg13g2_nand2_1 _20002_ (.Y(_06422_),
    .A(net6935),
    .B(_06410_));
 sg13g2_a21oi_1 _20003_ (.A1(_06415_),
    .A2(_06422_),
    .Y(_06423_),
    .B1(net6993));
 sg13g2_a21oi_1 _20004_ (.A1(net6897),
    .A2(_06410_),
    .Y(_06424_),
    .B1(_06423_));
 sg13g2_o21ai_1 _20005_ (.B1(_06420_),
    .Y(_06425_),
    .A1(net7000),
    .A2(_06424_));
 sg13g2_xnor2_1 _20006_ (.Y(_06426_),
    .A(_06360_),
    .B(_06425_));
 sg13g2_a21oi_1 _20007_ (.A1(_01667_),
    .A2(net7322),
    .Y(_06427_),
    .B1(net7317));
 sg13g2_a21o_1 _20008_ (.A2(net7322),
    .A1(_01667_),
    .B1(net7317),
    .X(_06428_));
 sg13g2_o21ai_1 _20009_ (.B1(net6942),
    .Y(_06429_),
    .A1(_06305_),
    .A2(net7109));
 sg13g2_nand2b_1 _20010_ (.Y(_06430_),
    .B(_06429_),
    .A_N(_06365_));
 sg13g2_a22oi_1 _20011_ (.Y(_06431_),
    .B1(_06430_),
    .B2(net6993),
    .A2(_06364_),
    .A1(net6935));
 sg13g2_nor2_1 _20012_ (.A(net6997),
    .B(_06431_),
    .Y(_06432_));
 sg13g2_inv_1 _20013_ (.Y(_06433_),
    .A(_00159_));
 sg13g2_nand3_1 _20014_ (.B(net6935),
    .C(net7109),
    .A(net7054),
    .Y(_06434_));
 sg13g2_o21ai_1 _20015_ (.B1(_06434_),
    .Y(_06435_),
    .A1(net7054),
    .A2(_06415_));
 sg13g2_a21oi_1 _20016_ (.A1(net6997),
    .A2(_06435_),
    .Y(_06436_),
    .B1(_06432_));
 sg13g2_xnor2_1 _20017_ (.Y(_06437_),
    .A(_06428_),
    .B(_06436_));
 sg13g2_inv_1 _20018_ (.Y(_06438_),
    .A(_00158_));
 sg13g2_xnor2_1 _20019_ (.Y(_06439_),
    .A(net6892),
    .B(_06437_));
 sg13g2_xnor2_1 _20020_ (.Y(_06440_),
    .A(_06426_),
    .B(_06439_));
 sg13g2_nor2_1 _20021_ (.A(_06333_),
    .B(_06339_),
    .Y(_06441_));
 sg13g2_nand2_1 _20022_ (.Y(_06442_),
    .A(_06333_),
    .B(_06339_));
 sg13g2_o21ai_1 _20023_ (.B1(_06442_),
    .Y(_06443_),
    .A1(net6889),
    .A2(_06441_));
 sg13g2_inv_1 _20024_ (.Y(_06444_),
    .A(_00157_));
 sg13g2_a21o_1 _20025_ (.A2(_06256_),
    .A1(net7133),
    .B1(net7134),
    .X(_06445_));
 sg13g2_nand3_1 _20026_ (.B(_06206_),
    .C(_06445_),
    .A(net7142),
    .Y(_06446_));
 sg13g2_nand2_1 _20027_ (.Y(_06447_),
    .A(net7118),
    .B(_06446_));
 sg13g2_o21ai_1 _20028_ (.B1(_06447_),
    .Y(_06448_),
    .A1(_04744_),
    .A2(net7118));
 sg13g2_inv_1 _20029_ (.Y(_06449_),
    .A(_00156_));
 sg13g2_xnor2_1 _20030_ (.Y(_06450_),
    .A(net6889),
    .B(_06448_));
 sg13g2_xnor2_1 _20031_ (.Y(_06451_),
    .A(_06277_),
    .B(_06450_));
 sg13g2_xnor2_1 _20032_ (.Y(_06452_),
    .A(_06443_),
    .B(_06451_));
 sg13g2_a21o_1 _20033_ (.A2(_06343_),
    .A1(_06340_),
    .B1(_06278_),
    .X(_06453_));
 sg13g2_inv_1 _20034_ (.Y(_06454_),
    .A(_00155_));
 sg13g2_o21ai_1 _20035_ (.B1(_06453_),
    .Y(_06455_),
    .A1(_06340_),
    .A2(_06343_));
 sg13g2_xnor2_1 _20036_ (.Y(_06456_),
    .A(_06452_),
    .B(_06455_));
 sg13g2_xnor2_1 _20037_ (.Y(_06457_),
    .A(_06440_),
    .B(_06456_));
 sg13g2_inv_1 _20038_ (.Y(_06458_),
    .A(_00152_));
 sg13g2_nor2_1 _20039_ (.A(_06347_),
    .B(_06378_),
    .Y(_06459_));
 sg13g2_nand2_1 _20040_ (.Y(_06460_),
    .A(_06347_),
    .B(_06378_));
 sg13g2_a21oi_1 _20041_ (.A1(_06346_),
    .A2(_06460_),
    .Y(_06461_),
    .B1(_06459_));
 sg13g2_xnor2_1 _20042_ (.Y(_06462_),
    .A(_06457_),
    .B(_06461_));
 sg13g2_xnor2_1 _20043_ (.Y(_06463_),
    .A(_06409_),
    .B(_06462_));
 sg13g2_nor2_1 _20044_ (.A(_06363_),
    .B(_06428_),
    .Y(_06464_));
 sg13g2_nor4_1 _20045_ (.A(net6936),
    .B(_06305_),
    .C(_06363_),
    .D(_06428_),
    .Y(_06465_));
 sg13g2_inv_1 _20046_ (.Y(_06466_),
    .A(_00148_));
 sg13g2_nor3_1 _20047_ (.A(net6940),
    .B(_06364_),
    .C(_06427_),
    .Y(_06467_));
 sg13g2_a21oi_1 _20048_ (.A1(net6940),
    .A2(_06427_),
    .Y(_06468_),
    .B1(_06467_));
 sg13g2_nand2_1 _20049_ (.Y(_06469_),
    .A(net6940),
    .B(_06428_));
 sg13g2_nand3_1 _20050_ (.B(_06306_),
    .C(_06427_),
    .A(net6936),
    .Y(_06470_));
 sg13g2_a21oi_1 _20051_ (.A1(_06469_),
    .A2(_06470_),
    .Y(_06471_),
    .B1(_06364_));
 sg13g2_inv_1 _20052_ (.Y(_06472_),
    .A(_00147_));
 sg13g2_nor2_1 _20053_ (.A(net7056),
    .B(_06471_),
    .Y(_06473_));
 sg13g2_a21oi_1 _20054_ (.A1(net7056),
    .A2(_06468_),
    .Y(_06474_),
    .B1(_06473_));
 sg13g2_o21ai_1 _20055_ (.B1(net7000),
    .Y(_06475_),
    .A1(_06465_),
    .A2(_06474_));
 sg13g2_nand2_1 _20056_ (.Y(_06476_),
    .A(net6936),
    .B(_06464_));
 sg13g2_nand2_1 _20057_ (.Y(_06477_),
    .A(_06469_),
    .B(_06476_));
 sg13g2_a22oi_1 _20058_ (.Y(_06478_),
    .B1(_06477_),
    .B2(net7056),
    .A2(_06464_),
    .A1(net6897));
 sg13g2_o21ai_1 _20059_ (.B1(_06475_),
    .Y(_06479_),
    .A1(net7000),
    .A2(_06478_));
 sg13g2_o21ai_1 _20060_ (.B1(net6940),
    .Y(_06480_),
    .A1(_06363_),
    .A2(_06427_));
 sg13g2_o21ai_1 _20061_ (.B1(_06480_),
    .Y(_06481_),
    .A1(net6940),
    .A2(_06363_));
 sg13g2_a22oi_1 _20062_ (.Y(_06482_),
    .B1(_06481_),
    .B2(net6993),
    .A2(_06428_),
    .A1(net6936));
 sg13g2_nand3_1 _20063_ (.B(net6936),
    .C(_06427_),
    .A(net7056),
    .Y(_06483_));
 sg13g2_o21ai_1 _20064_ (.B1(_06483_),
    .Y(_06484_),
    .A1(net7056),
    .A2(_06469_));
 sg13g2_nand2_1 _20065_ (.Y(_06485_),
    .A(net6997),
    .B(_06484_));
 sg13g2_o21ai_1 _20066_ (.B1(_06485_),
    .Y(_06486_),
    .A1(net6997),
    .A2(_06482_));
 sg13g2_a21oi_1 _20067_ (.A1(_01668_),
    .A2(net7321),
    .Y(_06487_),
    .B1(net7316));
 sg13g2_xor2_1 _20068_ (.B(_06487_),
    .A(_06486_),
    .X(_06488_));
 sg13g2_inv_1 _20069_ (.Y(_06489_),
    .A(_00144_));
 sg13g2_xnor2_1 _20070_ (.Y(_06490_),
    .A(_06479_),
    .B(_06488_));
 sg13g2_and2_1 _20071_ (.A(_06360_),
    .B(_06437_),
    .X(_06491_));
 sg13g2_nor2_1 _20072_ (.A(_06360_),
    .B(_06437_),
    .Y(_06492_));
 sg13g2_mux2_1 _20073_ (.A0(_06491_),
    .A1(_06492_),
    .S(_06425_),
    .X(_06493_));
 sg13g2_a21oi_1 _20074_ (.A1(net6892),
    .A2(_06426_),
    .Y(_06494_),
    .B1(_06493_));
 sg13g2_inv_1 _20075_ (.Y(_06495_),
    .A(_00143_));
 sg13g2_xnor2_1 _20076_ (.Y(_06496_),
    .A(_06490_),
    .B(_06494_));
 sg13g2_nand2b_1 _20077_ (.Y(_06497_),
    .B(_06448_),
    .A_N(_06443_));
 sg13g2_and2_1 _20078_ (.A(net6889),
    .B(_06277_),
    .X(_06498_));
 sg13g2_nor3_1 _20079_ (.A(net6889),
    .B(_06277_),
    .C(_06497_),
    .Y(_06499_));
 sg13g2_a21oi_1 _20080_ (.A1(_06497_),
    .A2(_06498_),
    .Y(_06500_),
    .B1(_06499_));
 sg13g2_xnor2_1 _20081_ (.Y(_06501_),
    .A(_06496_),
    .B(_06500_));
 sg13g2_inv_1 _20082_ (.Y(_06502_),
    .A(_00142_));
 sg13g2_nand2_1 _20083_ (.Y(_06503_),
    .A(_06452_),
    .B(_06455_));
 sg13g2_nor2_1 _20084_ (.A(_06452_),
    .B(_06455_),
    .Y(_06504_));
 sg13g2_a21oi_1 _20085_ (.A1(_06440_),
    .A2(_06503_),
    .Y(_06505_),
    .B1(_06504_));
 sg13g2_xnor2_1 _20086_ (.Y(_06506_),
    .A(_06501_),
    .B(_06505_));
 sg13g2_nor2_1 _20087_ (.A(_03928_),
    .B(_03929_),
    .Y(_06507_));
 sg13g2_inv_1 _20088_ (.Y(_06508_),
    .A(_00141_));
 sg13g2_a21oi_1 _20089_ (.A1(_04074_),
    .A2(_04139_),
    .Y(_06509_),
    .B1(_04138_));
 sg13g2_o21ai_1 _20090_ (.B1(_04209_),
    .Y(_06510_),
    .A1(_04205_),
    .A2(_04208_));
 sg13g2_a21oi_1 _20091_ (.A1(_04277_),
    .A2(_04284_),
    .Y(_06511_),
    .B1(_04285_));
 sg13g2_inv_1 _20092_ (.Y(_06512_),
    .A(_00140_));
 sg13g2_o21ai_1 _20093_ (.B1(_04361_),
    .Y(_06513_),
    .A1(_04356_),
    .A2(_04362_));
 sg13g2_a21oi_1 _20094_ (.A1(_04435_),
    .A2(_04439_),
    .Y(_06514_),
    .B1(_04440_));
 sg13g2_o21ai_1 _20095_ (.B1(_04520_),
    .Y(_06515_),
    .A1(_04516_),
    .A2(_04521_));
 sg13g2_a21oi_1 _20096_ (.A1(_04597_),
    .A2(_04602_),
    .Y(_06516_),
    .B1(_04601_));
 sg13g2_a21oi_1 _20097_ (.A1(_04701_),
    .A2(_04702_),
    .Y(_06517_),
    .B1(_04700_));
 sg13g2_nand3_1 _20098_ (.B(_04701_),
    .C(_04702_),
    .A(_04700_),
    .Y(_06518_));
 sg13g2_o21ai_1 _20099_ (.B1(_06518_),
    .Y(_06519_),
    .A1(_04699_),
    .A2(_06517_));
 sg13g2_o21ai_1 _20100_ (.B1(_04828_),
    .Y(_06520_),
    .A1(_04824_),
    .A2(_04829_));
 sg13g2_inv_1 _20101_ (.Y(_06521_),
    .A(_00138_));
 sg13g2_o21ai_1 _20102_ (.B1(_04943_),
    .Y(_06522_),
    .A1(_04945_),
    .A2(_04946_));
 sg13g2_nand2_1 _20103_ (.Y(_06523_),
    .A(_04947_),
    .B(_06522_));
 sg13g2_a21o_1 _20104_ (.A2(_05049_),
    .A1(_05042_),
    .B1(_05048_),
    .X(_06524_));
 sg13g2_a21oi_1 _20105_ (.A1(_05164_),
    .A2(_05170_),
    .Y(_06525_),
    .B1(_05169_));
 sg13g2_a21oi_1 _20106_ (.A1(_05268_),
    .A2(_05273_),
    .Y(_06526_),
    .B1(_05272_));
 sg13g2_inv_1 _20107_ (.Y(_06527_),
    .A(_00136_));
 sg13g2_a21oi_1 _20108_ (.A1(_05396_),
    .A2(_05414_),
    .Y(_06528_),
    .B1(_05410_));
 sg13g2_a22oi_1 _20109_ (.Y(_06529_),
    .B1(_05525_),
    .B2(_05518_),
    .A2(_05521_),
    .A1(_05394_));
 sg13g2_a21oi_1 _20110_ (.A1(_05519_),
    .A2(_05524_),
    .Y(_06530_),
    .B1(_06529_));
 sg13g2_nand2b_1 _20111_ (.Y(_06531_),
    .B(_05627_),
    .A_N(_05624_));
 sg13g2_inv_1 _20112_ (.Y(_06532_),
    .A(_00134_));
 sg13g2_nor2b_1 _20113_ (.A(_05627_),
    .B_N(_05624_),
    .Y(_06533_));
 sg13g2_a21oi_1 _20114_ (.A1(_05528_),
    .A2(_06531_),
    .Y(_06534_),
    .B1(_06533_));
 sg13g2_inv_1 _20115_ (.Y(_06535_),
    .A(_00133_));
 sg13g2_nand2_1 _20116_ (.Y(_06536_),
    .A(_05735_),
    .B(_05738_));
 sg13g2_a21oi_1 _20117_ (.A1(_05732_),
    .A2(_06536_),
    .Y(_06537_),
    .B1(_05739_));
 sg13g2_nand2_1 _20118_ (.Y(_06538_),
    .A(_05855_),
    .B(_05857_));
 sg13g2_a21oi_1 _20119_ (.A1(_05749_),
    .A2(_06538_),
    .Y(_06539_),
    .B1(_05859_));
 sg13g2_a21oi_1 _20120_ (.A1(_05868_),
    .A2(_05953_),
    .Y(_06540_),
    .B1(_05952_));
 sg13g2_o21ai_1 _20121_ (.B1(_06062_),
    .Y(_06541_),
    .A1(_05963_),
    .A2(_06061_));
 sg13g2_inv_1 _20122_ (.Y(_06542_),
    .A(_00131_));
 sg13g2_nand2_1 _20123_ (.Y(_06543_),
    .A(_06136_),
    .B(_06138_));
 sg13g2_nor2_1 _20124_ (.A(_06136_),
    .B(_06138_),
    .Y(_06544_));
 sg13g2_a21oi_1 _20125_ (.A1(_06070_),
    .A2(_06543_),
    .Y(_06545_),
    .B1(_06544_));
 sg13g2_nand2_1 _20126_ (.Y(_06546_),
    .A(_06159_),
    .B(_06232_));
 sg13g2_nor2_1 _20127_ (.A(_06159_),
    .B(_06232_),
    .Y(_06547_));
 sg13g2_inv_1 _20128_ (.Y(_06548_),
    .A(_00129_));
 sg13g2_a21o_1 _20129_ (.A2(_06546_),
    .A1(_06155_),
    .B1(_06547_),
    .X(_06549_));
 sg13g2_a21o_1 _20130_ (.A2(_06320_),
    .A1(_06316_),
    .B1(_06253_),
    .X(_06550_));
 sg13g2_o21ai_1 _20131_ (.B1(_06550_),
    .Y(_06551_),
    .A1(_06316_),
    .A2(_06320_));
 sg13g2_inv_1 _20132_ (.Y(_06552_),
    .A(_00128_));
 sg13g2_a21o_1 _20133_ (.A2(_06389_),
    .A1(_06381_),
    .B1(_06314_),
    .X(_06553_));
 sg13g2_o21ai_1 _20134_ (.B1(_06553_),
    .Y(_06554_),
    .A1(net6617),
    .A2(_06385_));
 sg13g2_nand2_1 _20135_ (.Y(_06555_),
    .A(net6617),
    .B(_06382_));
 sg13g2_inv_1 _20136_ (.Y(_06556_),
    .A(_00127_));
 sg13g2_o21ai_1 _20137_ (.B1(_06389_),
    .Y(_06557_),
    .A1(_06314_),
    .A2(_06385_));
 sg13g2_nor2_1 _20138_ (.A(net6617),
    .B(_06382_),
    .Y(_06558_));
 sg13g2_a221oi_1 _20139_ (.B2(_06557_),
    .C1(_06558_),
    .B1(_06555_),
    .A1(_06383_),
    .Y(_06559_),
    .A2(_06554_));
 sg13g2_a21oi_1 _20140_ (.A1(_06409_),
    .A2(_06461_),
    .Y(_06560_),
    .B1(_06457_));
 sg13g2_nor2_1 _20141_ (.A(_06409_),
    .B(_06461_),
    .Y(_06561_));
 sg13g2_nor2_1 _20142_ (.A(_06560_),
    .B(_06561_),
    .Y(_06562_));
 sg13g2_and2_1 _20143_ (.A(clknet_1_0__leaf_clk_i),
    .B(\core_clock_gate_i.en_latch ),
    .X(_06563_));
 sg13g2_nor2_1 _20144_ (.A(_05858_),
    .B(net7659),
    .Y(_06564_));
 sg13g2_or2_1 _20145_ (.X(_06565_),
    .B(_06564_),
    .A(_08623_));
 sg13g2_nor2b_1 _20146_ (.A(_01983_),
    .B_N(net348),
    .Y(_06566_));
 sg13g2_nand2_1 _20147_ (.Y(_06567_),
    .A(_06565_),
    .B(_06566_));
 sg13g2_nor2_1 _20148_ (.A(\load_store_unit_i.data_we_q ),
    .B(_06567_),
    .Y(_06568_));
 sg13g2_inv_1 _20149_ (.Y(_06569_),
    .A(_00125_));
 sg13g2_mux2_1 _20150_ (.A0(_02011_),
    .A1(net347),
    .S(net7108),
    .X(_06570_));
 sg13g2_mux2_1 _20151_ (.A0(_02010_),
    .A1(net346),
    .S(_06568_),
    .X(_06571_));
 sg13g2_mux2_1 _20152_ (.A0(_02009_),
    .A1(net340),
    .S(net7106),
    .X(_06572_));
 sg13g2_mux2_1 _20153_ (.A0(_02008_),
    .A1(net339),
    .S(net7107),
    .X(_06573_));
 sg13g2_inv_1 _20154_ (.Y(_06574_),
    .A(_00124_));
 sg13g2_mux2_1 _20155_ (.A0(_02007_),
    .A1(net337),
    .S(_06568_),
    .X(_06575_));
 sg13g2_mux2_1 _20156_ (.A0(_02006_),
    .A1(net336),
    .S(net7107),
    .X(_06576_));
 sg13g2_mux2_1 _20157_ (.A0(_02005_),
    .A1(net335),
    .S(net7107),
    .X(_06577_));
 sg13g2_mux2_1 _20158_ (.A0(_02004_),
    .A1(net334),
    .S(net7106),
    .X(_06578_));
 sg13g2_mux2_1 _20159_ (.A0(_02003_),
    .A1(net333),
    .S(net7108),
    .X(_06579_));
 sg13g2_mux2_1 _20160_ (.A0(_02002_),
    .A1(net332),
    .S(_06568_),
    .X(_06580_));
 sg13g2_mux2_1 _20161_ (.A0(_02001_),
    .A1(net331),
    .S(net7106),
    .X(_06581_));
 sg13g2_mux2_1 _20162_ (.A0(_02000_),
    .A1(net330),
    .S(net7108),
    .X(_06582_));
 sg13g2_mux2_1 _20163_ (.A0(_01999_),
    .A1(net329),
    .S(net7108),
    .X(_06583_));
 sg13g2_mux2_1 _20164_ (.A0(_01998_),
    .A1(net328),
    .S(net7107),
    .X(_06584_));
 sg13g2_inv_1 _20165_ (.Y(_06585_),
    .A(_00121_));
 sg13g2_mux2_1 _20166_ (.A0(_01997_),
    .A1(net326),
    .S(net7107),
    .X(_06586_));
 sg13g2_mux2_1 _20167_ (.A0(_01996_),
    .A1(net325),
    .S(net7106),
    .X(_06587_));
 sg13g2_mux2_1 _20168_ (.A0(_01995_),
    .A1(net324),
    .S(net7106),
    .X(_06588_));
 sg13g2_mux2_1 _20169_ (.A0(_01994_),
    .A1(net323),
    .S(_06568_),
    .X(_06589_));
 sg13g2_mux2_1 _20170_ (.A0(_01993_),
    .A1(net322),
    .S(net7106),
    .X(_06590_));
 sg13g2_mux2_1 _20171_ (.A0(_01992_),
    .A1(net321),
    .S(net7107),
    .X(_06591_));
 sg13g2_inv_1 _20172_ (.Y(_06592_),
    .A(_00119_));
 sg13g2_mux2_1 _20173_ (.A0(_01991_),
    .A1(net320),
    .S(net7106),
    .X(_06593_));
 sg13g2_mux2_1 _20174_ (.A0(_01990_),
    .A1(net319),
    .S(net7107),
    .X(_06594_));
 sg13g2_mux2_1 _20175_ (.A0(_01989_),
    .A1(net318),
    .S(net7107),
    .X(_06595_));
 sg13g2_mux2_1 _20176_ (.A0(_01988_),
    .A1(net317),
    .S(net7106),
    .X(_06596_));
 sg13g2_inv_1 _20177_ (.Y(_06597_),
    .A(_00118_));
 sg13g2_nor2_1 _20178_ (.A(\id_stage_i.controller_i.instr_fetch_err_i ),
    .B(_02232_),
    .Y(_06598_));
 sg13g2_nand2_1 _20179_ (.Y(_06599_),
    .A(net7665),
    .B(_06598_));
 sg13g2_nor2_1 _20180_ (.A(net7981),
    .B(_06599_),
    .Y(_06600_));
 sg13g2_o21ai_1 _20181_ (.B1(_08894_),
    .Y(_06601_),
    .A1(net7920),
    .A2(_07708_));
 sg13g2_a21oi_1 _20182_ (.A1(_07812_),
    .A2(_06601_),
    .Y(_06602_),
    .B1(_07619_));
 sg13g2_nor3_1 _20183_ (.A(net7676),
    .B(net7608),
    .C(net7607),
    .Y(_06603_));
 sg13g2_o21ai_1 _20184_ (.B1(_08645_),
    .Y(_06604_),
    .A1(_07890_),
    .A2(_06603_));
 sg13g2_nor3_1 _20185_ (.A(_07570_),
    .B(net7608),
    .C(_07844_),
    .Y(_06605_));
 sg13g2_o21ai_1 _20186_ (.B1(net7925),
    .Y(_06606_),
    .A1(net7674),
    .A2(_01890_));
 sg13g2_inv_1 _20187_ (.Y(_06607_),
    .A(_00116_));
 sg13g2_a21oi_1 _20188_ (.A1(_07680_),
    .A2(_06606_),
    .Y(_06608_),
    .B1(_08696_));
 sg13g2_nor4_1 _20189_ (.A(\id_stage_i.decoder_i.illegal_c_insn_i ),
    .B(_07562_),
    .C(_06605_),
    .D(_06608_),
    .Y(_06609_));
 sg13g2_nor2_1 _20190_ (.A(net7673),
    .B(_03635_),
    .Y(_06610_));
 sg13g2_o21ai_1 _20191_ (.B1(_08533_),
    .Y(_06611_),
    .A1(_07930_),
    .A2(_06610_));
 sg13g2_nand2_1 _20192_ (.Y(_06612_),
    .A(_03634_),
    .B(_06611_));
 sg13g2_a21o_1 _20193_ (.A2(_07665_),
    .A1(_07649_),
    .B1(_07973_),
    .X(_06613_));
 sg13g2_o21ai_1 _20194_ (.B1(_06609_),
    .Y(_06614_),
    .A1(_07701_),
    .A2(_06613_));
 sg13g2_inv_1 _20195_ (.Y(_06615_),
    .A(_00114_));
 sg13g2_a21oi_1 _20196_ (.A1(_07806_),
    .A2(_06602_),
    .Y(_06616_),
    .B1(_06614_));
 sg13g2_nand3_1 _20197_ (.B(_06612_),
    .C(_06616_),
    .A(_06604_),
    .Y(_06617_));
 sg13g2_nand3b_1 _20198_ (.B(_08973_),
    .C(net7473),
    .Y(_06618_),
    .A_N(net7839));
 sg13g2_nor2_1 _20199_ (.A(_01917_),
    .B(_01887_),
    .Y(_06619_));
 sg13g2_or2_1 _20200_ (.X(_06620_),
    .B(net7932),
    .A(net7666));
 sg13g2_nor2_1 _20201_ (.A(_01915_),
    .B(_01888_),
    .Y(_06621_));
 sg13g2_nand2_1 _20202_ (.Y(_06622_),
    .A(_08510_),
    .B(_09373_));
 sg13g2_nand2_1 _20203_ (.Y(_06623_),
    .A(_06619_),
    .B(_06621_));
 sg13g2_nor4_1 _20204_ (.A(_01916_),
    .B(_01891_),
    .C(_06618_),
    .D(_06623_),
    .Y(_06624_));
 sg13g2_nor2b_1 _20205_ (.A(net7685),
    .B_N(_07834_),
    .Y(_06625_));
 sg13g2_and3_1 _20206_ (.X(_06626_),
    .A(net7517),
    .B(_08305_),
    .C(_06625_));
 sg13g2_nand2_1 _20207_ (.Y(_06627_),
    .A(net7681),
    .B(net7531));
 sg13g2_inv_1 _20208_ (.Y(_06628_),
    .A(_00112_));
 sg13g2_nand3b_1 _20209_ (.B(net7699),
    .C(net7597),
    .Y(_06629_),
    .A_N(net7680));
 sg13g2_nand3b_1 _20210_ (.B(_08313_),
    .C(_01907_),
    .Y(_06630_),
    .A_N(net7699));
 sg13g2_nor3_1 _20211_ (.A(net7677),
    .B(net7684),
    .C(net7685),
    .Y(_06631_));
 sg13g2_nand2_1 _20212_ (.Y(_06632_),
    .A(_07807_),
    .B(_06631_));
 sg13g2_nor2b_1 _20213_ (.A(net7683),
    .B_N(net7682),
    .Y(_06633_));
 sg13g2_nor2_1 _20214_ (.A(net7677),
    .B(_08711_),
    .Y(_06634_));
 sg13g2_nand4_1 _20215_ (.B(net7685),
    .C(_06633_),
    .A(net7684),
    .Y(_06635_),
    .D(_06634_));
 sg13g2_nand3_1 _20216_ (.B(net7681),
    .C(_10449_),
    .A(_01907_),
    .Y(_06636_));
 sg13g2_or2_1 _20217_ (.X(_06637_),
    .B(_06636_),
    .A(_06635_));
 sg13g2_a221oi_1 _20218_ (.B2(_06637_),
    .C1(_06627_),
    .B1(_06632_),
    .A1(_06629_),
    .Y(_06638_),
    .A2(_06630_));
 sg13g2_o21ai_1 _20219_ (.B1(_06624_),
    .Y(_06639_),
    .A1(_06626_),
    .A2(_06638_));
 sg13g2_and2_1 _20220_ (.A(_07655_),
    .B(_06639_),
    .X(_06640_));
 sg13g2_a21oi_1 _20221_ (.A1(_03638_),
    .A2(_06640_),
    .Y(_06641_),
    .B1(_06617_));
 sg13g2_nor2b_1 _20222_ (.A(_08696_),
    .B_N(_06641_),
    .Y(_06642_));
 sg13g2_and2_1 _20223_ (.A(_06600_),
    .B(_06642_),
    .X(_06643_));
 sg13g2_inv_1 _20224_ (.Y(_06644_),
    .A(_06643_));
 sg13g2_nor2_1 _20225_ (.A(net7659),
    .B(_06644_),
    .Y(_06645_));
 sg13g2_nor2_1 _20226_ (.A(net7660),
    .B(_06645_),
    .Y(_06646_));
 sg13g2_nor2b_1 _20227_ (.A(net7657),
    .B_N(net315),
    .Y(_06647_));
 sg13g2_nor2b_1 _20228_ (.A(_06646_),
    .B_N(_06647_),
    .Y(_06648_));
 sg13g2_mux2_1 _20229_ (.A0(_01987_),
    .A1(net6727),
    .S(_06648_),
    .X(_06649_));
 sg13g2_mux2_1 _20230_ (.A0(net7650),
    .A1(net6746),
    .S(_06648_),
    .X(_06650_));
 sg13g2_a22oi_1 _20231_ (.Y(_06651_),
    .B1(_06645_),
    .B2(_05858_),
    .A2(_06565_),
    .A1(net348));
 sg13g2_nor2_1 _20232_ (.A(net7660),
    .B(_06651_),
    .Y(_06652_));
 sg13g2_nand3_1 _20233_ (.B(_06565_),
    .C(_06652_),
    .A(net314),
    .Y(_06653_));
 sg13g2_o21ai_1 _20234_ (.B1(_06653_),
    .Y(_06654_),
    .A1(_05828_),
    .A2(_06652_));
 sg13g2_a21oi_1 _20235_ (.A1(net7659),
    .A2(_06647_),
    .Y(_06655_),
    .B1(_06564_));
 sg13g2_nor3_1 _20236_ (.A(net348),
    .B(net7660),
    .C(_06655_),
    .Y(_06656_));
 sg13g2_inv_1 _20237_ (.Y(_06657_),
    .A(_06658_));
 sg13g2_nand2b_1 _20238_ (.Y(_06658_),
    .B(_09282_),
    .A_N(_08696_));
 sg13g2_or2_1 _20239_ (.X(_06659_),
    .B(\alu_adder_result_ex[1] ),
    .A(\alu_adder_result_ex[0] ));
 sg13g2_nand2_1 _20240_ (.Y(_06660_),
    .A(_06658_),
    .B(_06659_));
 sg13g2_nand3_1 _20241_ (.B(net6747),
    .C(net6726),
    .A(_01889_),
    .Y(_06661_));
 sg13g2_nand2_1 _20242_ (.Y(_06662_),
    .A(_06660_),
    .B(_06661_));
 sg13g2_a21oi_1 _20243_ (.A1(_06643_),
    .A2(_06662_),
    .Y(_06663_),
    .B1(net7660));
 sg13g2_o21ai_1 _20244_ (.B1(net315),
    .Y(_06664_),
    .A1(net7658),
    .A2(_06663_));
 sg13g2_nor2_1 _20245_ (.A(net7660),
    .B(_06662_),
    .Y(_06665_));
 sg13g2_a21o_1 _20246_ (.A2(_06665_),
    .A1(_06643_),
    .B1(net7658),
    .X(_06666_));
 sg13g2_o21ai_1 _20247_ (.B1(_06664_),
    .Y(_06667_),
    .A1(net315),
    .A2(_06666_));
 sg13g2_nor2_1 _20248_ (.A(net7657),
    .B(_06667_),
    .Y(_06668_));
 sg13g2_or2_1 _20249_ (.X(_06669_),
    .B(net7657),
    .A(net315));
 sg13g2_nand2_1 _20250_ (.Y(_06670_),
    .A(net348),
    .B(net7658));
 sg13g2_a21oi_1 _20251_ (.A1(_06646_),
    .A2(_06670_),
    .Y(_06671_),
    .B1(_06669_));
 sg13g2_nand3b_1 _20252_ (.B(net7658),
    .C(_06566_),
    .Y(_06672_),
    .A_N(net315));
 sg13g2_o21ai_1 _20253_ (.B1(_06672_),
    .Y(_06673_),
    .A1(net7658),
    .A2(_06665_));
 sg13g2_o21ai_1 _20254_ (.B1(net7658),
    .Y(_06674_),
    .A1(net315),
    .A2(_06566_));
 sg13g2_or2_1 _20255_ (.X(_06675_),
    .B(_06643_),
    .A(net7660));
 sg13g2_nand2_1 _20256_ (.Y(_06676_),
    .A(net315),
    .B(_06675_));
 sg13g2_a21oi_1 _20257_ (.A1(_06674_),
    .A2(_06676_),
    .Y(_06677_),
    .B1(net7657));
 sg13g2_nand2_1 _20258_ (.Y(_06678_),
    .A(_06673_),
    .B(_06677_));
 sg13g2_o21ai_1 _20259_ (.B1(_06678_),
    .Y(_06679_),
    .A1(_05957_),
    .A2(_06677_));
 sg13g2_and2_1 _20260_ (.A(net7673),
    .B(_06642_),
    .X(net507));
 sg13g2_mux2_1 _20261_ (.A0(\load_store_unit_i.data_we_q ),
    .A1(net507),
    .S(_06648_),
    .X(_06680_));
 sg13g2_nor2_1 _20262_ (.A(_07701_),
    .B(_08696_),
    .Y(_06681_));
 sg13g2_mux2_1 _20263_ (.A0(_01982_),
    .A1(_06681_),
    .S(_06648_),
    .X(_06682_));
 sg13g2_nor2_1 _20264_ (.A(_01889_),
    .B(_06658_),
    .Y(_06683_));
 sg13g2_nand2_1 _20265_ (.Y(_06684_),
    .A(_09324_),
    .B(_06657_));
 sg13g2_mux2_1 _20266_ (.A0(_01981_),
    .A1(_06683_),
    .S(_06648_),
    .X(_06685_));
 sg13g2_nand2_1 _20267_ (.Y(_06686_),
    .A(_06648_),
    .B(_06657_));
 sg13g2_o21ai_1 _20268_ (.B1(_06686_),
    .Y(_06687_),
    .A1(net7628),
    .A2(_06648_));
 sg13g2_nor4_1 _20269_ (.A(net7675),
    .B(_01891_),
    .C(_07575_),
    .D(_07872_),
    .Y(_06688_));
 sg13g2_mux2_1 _20270_ (.A0(\load_store_unit_i.data_sign_ext_q ),
    .A1(_06688_),
    .S(_06648_),
    .X(_06689_));
 sg13g2_nor2_1 _20271_ (.A(net314),
    .B(_05858_),
    .Y(_06690_));
 sg13g2_a22oi_1 _20272_ (.Y(_06691_),
    .B1(_06690_),
    .B2(_06566_),
    .A2(_06675_),
    .A1(_06647_));
 sg13g2_nand2b_1 _20273_ (.Y(_06692_),
    .B(net7660),
    .A_N(\load_store_unit_i.lsu_err_q ));
 sg13g2_nand2b_1 _20274_ (.Y(_06693_),
    .B(net348),
    .A_N(net314));
 sg13g2_o21ai_1 _20275_ (.B1(_06692_),
    .Y(_06694_),
    .A1(net7660),
    .A2(_06693_));
 sg13g2_nand3_1 _20276_ (.B(_06647_),
    .C(_06694_),
    .A(net7659),
    .Y(_06695_));
 sg13g2_o21ai_1 _20277_ (.B1(_06695_),
    .Y(_06696_),
    .A1(net7659),
    .A2(_06691_));
 sg13g2_mux2_1 _20278_ (.A0(_01980_),
    .A1(net6624),
    .S(net6736),
    .X(_06697_));
 sg13g2_mux2_1 _20279_ (.A0(_01979_),
    .A1(net6626),
    .S(net6737),
    .X(_06698_));
 sg13g2_mux2_1 _20280_ (.A0(_01978_),
    .A1(net467),
    .S(net6737),
    .X(_06699_));
 sg13g2_mux2_1 _20281_ (.A0(_01977_),
    .A1(net6628),
    .S(net6737),
    .X(_06700_));
 sg13g2_mux2_1 _20282_ (.A0(_01976_),
    .A1(net6637),
    .S(net6737),
    .X(_06701_));
 sg13g2_mux2_1 _20283_ (.A0(_01975_),
    .A1(net464),
    .S(net6736),
    .X(_06702_));
 sg13g2_mux2_1 _20284_ (.A0(_01974_),
    .A1(net6639),
    .S(_06696_),
    .X(_06703_));
 sg13g2_mux2_1 _20285_ (.A0(_01973_),
    .A1(net6567),
    .S(net6737),
    .X(_06704_));
 sg13g2_mux2_1 _20286_ (.A0(_01972_),
    .A1(net6570),
    .S(net6737),
    .X(_06705_));
 sg13g2_mux2_1 _20287_ (.A0(_01971_),
    .A1(net6640),
    .S(net6736),
    .X(_06706_));
 sg13g2_mux2_1 _20288_ (.A0(_01970_),
    .A1(net6571),
    .S(net6738),
    .X(_06707_));
 sg13g2_mux2_1 _20289_ (.A0(_01969_),
    .A1(net6573),
    .S(net6739),
    .X(_06708_));
 sg13g2_mux2_1 _20290_ (.A0(_01968_),
    .A1(net6575),
    .S(net6739),
    .X(_06709_));
 sg13g2_mux2_1 _20291_ (.A0(_01967_),
    .A1(net6576),
    .S(net6738),
    .X(_06710_));
 sg13g2_mux2_1 _20292_ (.A0(_01966_),
    .A1(net6579),
    .S(net6738),
    .X(_06711_));
 sg13g2_mux2_1 _20293_ (.A0(_01965_),
    .A1(net6582),
    .S(net6738),
    .X(_06712_));
 sg13g2_mux2_1 _20294_ (.A0(_01964_),
    .A1(net6603),
    .S(net6738),
    .X(_06713_));
 sg13g2_mux2_1 _20295_ (.A0(_01963_),
    .A1(net6605),
    .S(net6738),
    .X(_06714_));
 sg13g2_mux2_1 _20296_ (.A0(_01962_),
    .A1(net6584),
    .S(net6738),
    .X(_06715_));
 sg13g2_mux2_1 _20297_ (.A0(_01961_),
    .A1(net6586),
    .S(net6738),
    .X(_06716_));
 sg13g2_mux2_1 _20298_ (.A0(_01960_),
    .A1(net6727),
    .S(_06696_),
    .X(_06717_));
 sg13g2_mux2_1 _20299_ (.A0(_01959_),
    .A1(net6607),
    .S(net6739),
    .X(_06718_));
 sg13g2_mux2_1 _20300_ (.A0(_01958_),
    .A1(net6608),
    .S(net6739),
    .X(_06719_));
 sg13g2_mux2_1 _20301_ (.A0(_01957_),
    .A1(net6609),
    .S(net6737),
    .X(_06720_));
 sg13g2_mux2_1 _20302_ (.A0(_01956_),
    .A1(net6610),
    .S(net6737),
    .X(_06721_));
 sg13g2_mux2_1 _20303_ (.A0(_01955_),
    .A1(net6613),
    .S(net6736),
    .X(_06722_));
 sg13g2_mux2_1 _20304_ (.A0(_01954_),
    .A1(net6615),
    .S(_06696_),
    .X(_06723_));
 sg13g2_mux2_1 _20305_ (.A0(_01953_),
    .A1(net443),
    .S(net6736),
    .X(_06724_));
 sg13g2_mux2_1 _20306_ (.A0(_01952_),
    .A1(net6601),
    .S(net6736),
    .X(_06725_));
 sg13g2_mux2_1 _20307_ (.A0(_01951_),
    .A1(net6621),
    .S(net6736),
    .X(_06726_));
 sg13g2_mux2_1 _20308_ (.A0(_01950_),
    .A1(net6622),
    .S(net6736),
    .X(_06727_));
 sg13g2_mux2_1 _20309_ (.A0(_01949_),
    .A1(net6746),
    .S(_06696_),
    .X(_06728_));
 sg13g2_nor4_1 _20310_ (.A(net6639),
    .B(net465),
    .C(net467),
    .D(net469),
    .Y(_06729_));
 sg13g2_nor2_1 _20311_ (.A(net6640),
    .B(_06659_),
    .Y(_06730_));
 sg13g2_nor4_1 _20312_ (.A(net464),
    .B(net466),
    .C(net6621),
    .D(net6609),
    .Y(_06731_));
 sg13g2_or2_1 _20313_ (.X(_06732_),
    .B(net443),
    .A(net442));
 sg13g2_nor4_1 _20314_ (.A(net444),
    .B(net6613),
    .C(net6607),
    .D(_06732_),
    .Y(_06733_));
 sg13g2_nand4_1 _20315_ (.B(_06730_),
    .C(_06731_),
    .A(_06729_),
    .Y(_06734_),
    .D(_06733_));
 sg13g2_nor2_1 _20316_ (.A(net468),
    .B(net6622),
    .Y(_06735_));
 sg13g2_nor3_1 _20317_ (.A(net6580),
    .B(net6575),
    .C(net6571),
    .Y(_06736_));
 sg13g2_nor4_1 _20318_ (.A(net446),
    .B(net6608),
    .C(net6584),
    .D(net6604),
    .Y(_06737_));
 sg13g2_nand3_1 _20319_ (.B(_06736_),
    .C(_06737_),
    .A(_06735_),
    .Y(_06738_));
 sg13g2_or4_1 _20320_ (.A(net6583),
    .B(net6577),
    .C(net6573),
    .D(net6570),
    .X(_06739_));
 sg13g2_or3_1 _20321_ (.A(net6586),
    .B(net6605),
    .C(net6567),
    .X(_06740_));
 sg13g2_nor4_2 _20322_ (.A(_06734_),
    .B(_06738_),
    .C(_06739_),
    .Y(_06741_),
    .D(_06740_));
 sg13g2_nor3_1 _20323_ (.A(_07605_),
    .B(_08028_),
    .C(_06741_),
    .Y(_06742_));
 sg13g2_nor2_1 _20324_ (.A(net7046),
    .B(net7104),
    .Y(_06743_));
 sg13g2_xnor2_1 _20325_ (.Y(_06744_),
    .A(_08153_),
    .B(_06743_));
 sg13g2_nand2_1 _20326_ (.Y(_06745_),
    .A(_07844_),
    .B(_08028_));
 sg13g2_o21ai_1 _20327_ (.B1(net7438),
    .Y(_06746_),
    .A1(_06744_),
    .A2(_06745_));
 sg13g2_and3_1 _20328_ (.X(_06747_),
    .A(_08010_),
    .B(_06741_),
    .C(_06746_));
 sg13g2_nand2_1 _20329_ (.Y(_06748_),
    .A(net7046),
    .B(_08158_));
 sg13g2_nor2_1 _20330_ (.A(net7046),
    .B(_08158_),
    .Y(_06749_));
 sg13g2_inv_1 _20331_ (.Y(_06750_),
    .A(_06749_));
 sg13g2_nand3_1 _20332_ (.B(_07844_),
    .C(_06749_),
    .A(net7438),
    .Y(_06751_));
 sg13g2_a21oi_1 _20333_ (.A1(_06748_),
    .A2(_06751_),
    .Y(_06752_),
    .B1(net7104));
 sg13g2_nand2b_1 _20334_ (.Y(_06753_),
    .B(_03811_),
    .A_N(_03611_));
 sg13g2_nand2_1 _20335_ (.Y(_06754_),
    .A(_03611_),
    .B(_03812_));
 sg13g2_mux2_1 _20336_ (.A0(_06754_),
    .A1(_06753_),
    .S(_06752_),
    .X(_06755_));
 sg13g2_nand2_1 _20337_ (.Y(_06756_),
    .A(_06753_),
    .B(_06754_));
 sg13g2_o21ai_1 _20338_ (.B1(_06755_),
    .Y(_06757_),
    .A1(net6567),
    .A2(_06756_));
 sg13g2_xor2_1 _20339_ (.B(net7104),
    .A(net7046),
    .X(_06758_));
 sg13g2_nand3_1 _20340_ (.B(_08158_),
    .C(net7104),
    .A(net7046),
    .Y(_06759_));
 sg13g2_nand3_1 _20341_ (.B(_08158_),
    .C(_06758_),
    .A(_07844_),
    .Y(_06760_));
 sg13g2_mux2_1 _20342_ (.A0(_06759_),
    .A1(_06760_),
    .S(_06757_),
    .X(_06761_));
 sg13g2_o21ai_1 _20343_ (.B1(_07844_),
    .Y(_06762_),
    .A1(net7104),
    .A2(_06750_));
 sg13g2_nand2b_1 _20344_ (.Y(_06763_),
    .B(_06762_),
    .A_N(_06757_));
 sg13g2_a21oi_1 _20345_ (.A1(_06761_),
    .A2(_06763_),
    .Y(_06764_),
    .B1(_07605_));
 sg13g2_nor2_1 _20346_ (.A(_08010_),
    .B(_06757_),
    .Y(_06765_));
 sg13g2_nor4_2 _20347_ (.A(_06742_),
    .B(_06747_),
    .C(_06764_),
    .Y(_06766_),
    .D(_06765_));
 sg13g2_nor2b_1 _20348_ (.A(_06599_),
    .B_N(_06641_),
    .Y(_06767_));
 sg13g2_nand2b_1 _20349_ (.Y(_06768_),
    .B(_06641_),
    .A_N(_06599_));
 sg13g2_nand3_1 _20350_ (.B(_07595_),
    .C(_06767_),
    .A(_02201_),
    .Y(_06769_));
 sg13g2_nand2_1 _20351_ (.Y(_06770_),
    .A(_07792_),
    .B(_03638_));
 sg13g2_nor2_1 _20352_ (.A(_08444_),
    .B(_06770_),
    .Y(_06771_));
 sg13g2_a21oi_1 _20353_ (.A1(_10165_),
    .A2(_06641_),
    .Y(_06772_),
    .B1(_08444_));
 sg13g2_and3_1 _20354_ (.X(_06773_),
    .A(net7665),
    .B(net7607),
    .C(_03638_));
 sg13g2_nand3_1 _20355_ (.B(net7607),
    .C(_03638_),
    .A(net7665),
    .Y(_06774_));
 sg13g2_nor2_1 _20356_ (.A(_06637_),
    .B(_06774_),
    .Y(_06775_));
 sg13g2_nand2_1 _20357_ (.Y(_06776_),
    .A(_02226_),
    .B(net7105));
 sg13g2_nor2_1 _20358_ (.A(_00243_),
    .B(_00242_),
    .Y(_06777_));
 sg13g2_nor3_1 _20359_ (.A(_06632_),
    .B(_06636_),
    .C(_06774_),
    .Y(_06778_));
 sg13g2_nor4_1 _20360_ (.A(_06627_),
    .B(_06629_),
    .C(_06632_),
    .D(_06774_),
    .Y(_06779_));
 sg13g2_a21oi_1 _20361_ (.A1(\cs_registers_i.csr_mstatus_tw_o ),
    .A2(_06779_),
    .Y(_06780_),
    .B1(net7313));
 sg13g2_o21ai_1 _20362_ (.B1(_06776_),
    .Y(_06781_),
    .A1(_06777_),
    .A2(_06780_));
 sg13g2_and2_1 _20363_ (.A(_06626_),
    .B(_06773_),
    .X(_06782_));
 sg13g2_nor3_1 _20364_ (.A(_06772_),
    .B(_06781_),
    .C(_06782_),
    .Y(_06783_));
 sg13g2_nor2_1 _20365_ (.A(net6901),
    .B(net6952),
    .Y(_06784_));
 sg13g2_nand2_1 _20366_ (.Y(_06785_),
    .A(_10789_),
    .B(_11684_));
 sg13g2_nor3_1 _20367_ (.A(_06617_),
    .B(_06640_),
    .C(_06770_),
    .Y(_06786_));
 sg13g2_inv_1 _20368_ (.Y(_06787_),
    .A(_06786_));
 sg13g2_inv_1 _20369_ (.Y(_06788_),
    .A(_06789_));
 sg13g2_nand2_1 _20370_ (.Y(_06789_),
    .A(_15514_),
    .B(net6932));
 sg13g2_nor2_1 _20371_ (.A(_08874_),
    .B(net6903),
    .Y(_06790_));
 sg13g2_nand2_1 _20372_ (.Y(_06791_),
    .A(net6977),
    .B(_09944_));
 sg13g2_nand2_1 _20373_ (.Y(_06792_),
    .A(net6931),
    .B(_06790_));
 sg13g2_nand2_1 _20374_ (.Y(_06793_),
    .A(net6901),
    .B(net6953));
 sg13g2_o21ai_1 _20375_ (.B1(_06789_),
    .Y(_06794_),
    .A1(_06792_),
    .A2(_06793_));
 sg13g2_a22oi_1 _20376_ (.Y(_06795_),
    .B1(_06794_),
    .B2(net6951),
    .A2(_06788_),
    .A1(_06784_));
 sg13g2_or3_1 _20377_ (.A(net6948),
    .B(net6899),
    .C(_06795_),
    .X(_06796_));
 sg13g2_nand2_1 _20378_ (.Y(_06797_),
    .A(_08641_),
    .B(_08845_));
 sg13g2_nand3_1 _20379_ (.B(_08639_),
    .C(net7077),
    .A(net7103),
    .Y(_06798_));
 sg13g2_a21o_1 _20380_ (.A2(_06798_),
    .A1(_06797_),
    .B1(_09428_),
    .X(_06799_));
 sg13g2_nand2b_1 _20381_ (.Y(_06800_),
    .B(_10789_),
    .A_N(_06799_));
 sg13g2_nor2_1 _20382_ (.A(net6953),
    .B(_06800_),
    .Y(_06801_));
 sg13g2_nor2_1 _20383_ (.A(net6888),
    .B(_06801_),
    .Y(_06802_));
 sg13g2_inv_1 _20384_ (.Y(_06803_),
    .A(_06802_));
 sg13g2_o21ai_1 _20385_ (.B1(net7292),
    .Y(_06804_),
    .A1(net7274),
    .A2(net7272));
 sg13g2_o21ai_1 _20386_ (.B1(net7039),
    .Y(_06805_),
    .A1(net7682),
    .A2(net7683));
 sg13g2_nand2_1 _20387_ (.Y(_06806_),
    .A(_06804_),
    .B(_06805_));
 sg13g2_nand3_1 _20388_ (.B(_06804_),
    .C(_06805_),
    .A(_12822_),
    .Y(_06807_));
 sg13g2_nand2_1 _20389_ (.Y(_06808_),
    .A(net6931),
    .B(_06807_));
 sg13g2_nor2_1 _20390_ (.A(_09944_),
    .B(net6952),
    .Y(_06809_));
 sg13g2_nand2_1 _20391_ (.Y(_06810_),
    .A(net6903),
    .B(_11684_));
 sg13g2_nand2_1 _20392_ (.Y(_06811_),
    .A(_13840_),
    .B(net6932));
 sg13g2_nand2_1 _20393_ (.Y(_06812_),
    .A(net6899),
    .B(_15516_));
 sg13g2_inv_1 _20394_ (.Y(_06813_),
    .A(_06814_));
 sg13g2_nand2b_1 _20395_ (.Y(_06814_),
    .B(_06786_),
    .A_N(_10787_));
 sg13g2_nand2b_1 _20396_ (.Y(_06815_),
    .B(net6948),
    .A_N(_06807_));
 sg13g2_nor2_1 _20397_ (.A(_06814_),
    .B(_06815_),
    .Y(_06816_));
 sg13g2_nand2_1 _20398_ (.Y(_06817_),
    .A(_12822_),
    .B(net6899));
 sg13g2_or3_1 _20399_ (.A(_15514_),
    .B(net6887),
    .C(_06817_),
    .X(_06818_));
 sg13g2_nor3_1 _20400_ (.A(net6976),
    .B(net6901),
    .C(_06818_),
    .Y(_06819_));
 sg13g2_or2_1 _20401_ (.X(_06820_),
    .B(_06819_),
    .A(_06816_));
 sg13g2_a22oi_1 _20402_ (.Y(_06821_),
    .B1(_06809_),
    .B2(_06820_),
    .A2(_06808_),
    .A1(_06803_));
 sg13g2_nand2_1 _20403_ (.Y(_06822_),
    .A(_06784_),
    .B(_06790_));
 sg13g2_nand3_1 _20404_ (.B(net6903),
    .C(net6900),
    .A(net6976),
    .Y(_06823_));
 sg13g2_xnor2_1 _20405_ (.Y(_06824_),
    .A(net6903),
    .B(_10789_));
 sg13g2_o21ai_1 _20406_ (.B1(_06823_),
    .Y(_06825_),
    .A1(net6976),
    .A2(_06824_));
 sg13g2_nor3_1 _20407_ (.A(net6903),
    .B(_06785_),
    .C(_06818_),
    .Y(_06826_));
 sg13g2_nor4_1 _20408_ (.A(_09944_),
    .B(net6952),
    .C(_06807_),
    .D(net6887),
    .Y(_06827_));
 sg13g2_o21ai_1 _20409_ (.B1(net6975),
    .Y(_06828_),
    .A1(_06826_),
    .A2(_06827_));
 sg13g2_nor3_1 _20410_ (.A(_15514_),
    .B(_06811_),
    .C(_06817_),
    .Y(_06829_));
 sg13g2_nand3b_1 _20411_ (.B(_06825_),
    .C(_11684_),
    .Y(_06830_),
    .A_N(_06818_));
 sg13g2_nand4_1 _20412_ (.B(_06821_),
    .C(_06828_),
    .A(_06796_),
    .Y(_06831_),
    .D(_06830_));
 sg13g2_a22oi_1 _20413_ (.Y(_06832_),
    .B1(_02031_),
    .B2(net7270),
    .A2(net7039),
    .A1(_01907_));
 sg13g2_nor2_1 _20414_ (.A(net7681),
    .B(_02031_),
    .Y(_06833_));
 sg13g2_or3_1 _20415_ (.A(_06787_),
    .B(_06832_),
    .C(_06833_),
    .X(_06834_));
 sg13g2_nor2_1 _20416_ (.A(net7031),
    .B(_06834_),
    .Y(_06835_));
 sg13g2_nand2_1 _20417_ (.Y(_06836_),
    .A(net7033),
    .B(_06835_));
 sg13g2_nor2b_1 _20418_ (.A(_06836_),
    .B_N(_06831_),
    .Y(_06837_));
 sg13g2_a21oi_1 _20419_ (.A1(net6900),
    .A2(net6952),
    .Y(_06838_),
    .B1(_09944_));
 sg13g2_nor2_1 _20420_ (.A(net6975),
    .B(net6903),
    .Y(_06839_));
 sg13g2_a221oi_1 _20421_ (.B2(net6901),
    .C1(_06815_),
    .B1(_06839_),
    .A1(net6975),
    .Y(_06840_),
    .A2(_06838_));
 sg13g2_or3_1 _20422_ (.A(_12822_),
    .B(_06806_),
    .C(net6887),
    .X(_06841_));
 sg13g2_nand3_1 _20423_ (.B(_06804_),
    .C(_06805_),
    .A(net6951),
    .Y(_06842_));
 sg13g2_nand2_1 _20424_ (.Y(_06843_),
    .A(net6930),
    .B(_06841_));
 sg13g2_nand3_1 _20425_ (.B(net6930),
    .C(_06790_),
    .A(_11684_),
    .Y(_06844_));
 sg13g2_a221oi_1 _20426_ (.B2(_06844_),
    .C1(_06840_),
    .B1(_06843_),
    .A1(_06816_),
    .Y(_06845_),
    .A2(_06839_));
 sg13g2_nor4_1 _20427_ (.A(net6903),
    .B(net6952),
    .C(net6887),
    .D(_06842_),
    .Y(_06846_));
 sg13g2_a21oi_1 _20428_ (.A1(net6903),
    .A2(_06816_),
    .Y(_06847_),
    .B1(_06846_));
 sg13g2_o21ai_1 _20429_ (.B1(_06845_),
    .Y(_06848_),
    .A1(_08874_),
    .A2(_06847_));
 sg13g2_nand3b_1 _20430_ (.B(net7033),
    .C(net7031),
    .Y(_06849_),
    .A_N(_06834_));
 sg13g2_nor2b_1 _20431_ (.A(_06849_),
    .B_N(_06848_),
    .Y(_06850_));
 sg13g2_o21ai_1 _20432_ (.B1(net6952),
    .Y(_06851_),
    .A1(_08874_),
    .A2(_10789_));
 sg13g2_o21ai_1 _20433_ (.B1(_06800_),
    .Y(_06852_),
    .A1(_10789_),
    .A2(net6952));
 sg13g2_a21oi_1 _20434_ (.A1(_09944_),
    .A2(_06851_),
    .Y(_06853_),
    .B1(_06852_));
 sg13g2_nand3_1 _20435_ (.B(_06790_),
    .C(_06813_),
    .A(net6952),
    .Y(_06854_));
 sg13g2_a21oi_1 _20436_ (.A1(net6950),
    .A2(_06854_),
    .Y(_06855_),
    .B1(_06853_));
 sg13g2_a21o_1 _20437_ (.A2(_06800_),
    .A1(net6953),
    .B1(net6950),
    .X(_06856_));
 sg13g2_nor2_1 _20438_ (.A(_06791_),
    .B(_06793_),
    .Y(_06857_));
 sg13g2_nor2_1 _20439_ (.A(net6887),
    .B(_06857_),
    .Y(_06858_));
 sg13g2_a221oi_1 _20440_ (.B2(_06858_),
    .C1(net6888),
    .B1(_06856_),
    .A1(net6948),
    .Y(_06859_),
    .A2(_06855_));
 sg13g2_nand3_1 _20441_ (.B(_13407_),
    .C(_06633_),
    .A(_08616_),
    .Y(_06860_));
 sg13g2_o21ai_1 _20442_ (.B1(_06860_),
    .Y(_06861_),
    .A1(_08616_),
    .A2(_15462_));
 sg13g2_nand2_1 _20443_ (.Y(_06862_),
    .A(net7432),
    .B(_06861_));
 sg13g2_nand3_1 _20444_ (.B(net6932),
    .C(_06861_),
    .A(net7432),
    .Y(_06863_));
 sg13g2_nor3_1 _20445_ (.A(_06849_),
    .B(_06859_),
    .C(_06863_),
    .Y(_06864_));
 sg13g2_inv_1 _20446_ (.Y(_06865_),
    .A(_06864_));
 sg13g2_nor2_1 _20447_ (.A(_06850_),
    .B(_06864_),
    .Y(_06866_));
 sg13g2_nand2b_1 _20448_ (.Y(_06867_),
    .B(_06866_),
    .A_N(_06837_));
 sg13g2_o21ai_1 _20449_ (.B1(net6931),
    .Y(_06868_),
    .A1(_06785_),
    .A2(_06790_));
 sg13g2_nand3_1 _20450_ (.B(_13838_),
    .C(_06861_),
    .A(net7432),
    .Y(_06869_));
 sg13g2_nand2_1 _20451_ (.Y(_06870_),
    .A(_02172_),
    .B(_06835_));
 sg13g2_or3_1 _20452_ (.A(net6949),
    .B(_06869_),
    .C(_06870_),
    .X(_06871_));
 sg13g2_or3_1 _20453_ (.A(net6948),
    .B(_06806_),
    .C(_06836_),
    .X(_06872_));
 sg13g2_o21ai_1 _20454_ (.B1(_06871_),
    .Y(_06873_),
    .A1(net6949),
    .A2(_06872_));
 sg13g2_nor2_1 _20455_ (.A(_06785_),
    .B(_06870_),
    .Y(_06874_));
 sg13g2_and4_1 _20456_ (.A(_09945_),
    .B(net6948),
    .C(net6899),
    .D(_06788_),
    .X(_06875_));
 sg13g2_nor4_1 _20457_ (.A(net6949),
    .B(net6948),
    .C(_06791_),
    .D(_06863_),
    .Y(_06876_));
 sg13g2_a21oi_1 _20458_ (.A1(net6949),
    .A2(_06875_),
    .Y(_06877_),
    .B1(_06876_));
 sg13g2_nor3_1 _20459_ (.A(_06785_),
    .B(_06870_),
    .C(_06877_),
    .Y(_06878_));
 sg13g2_a21o_1 _20460_ (.A2(_06873_),
    .A1(_06868_),
    .B1(_06878_),
    .X(_06879_));
 sg13g2_a221oi_1 _20461_ (.B2(net6950),
    .C1(_06872_),
    .B1(_06857_),
    .A1(_06784_),
    .Y(_06880_),
    .A2(_06791_));
 sg13g2_nor3_1 _20462_ (.A(net6975),
    .B(net6900),
    .C(_06810_),
    .Y(_06881_));
 sg13g2_inv_1 _20463_ (.Y(_06882_),
    .A(_06881_));
 sg13g2_nand2_1 _20464_ (.Y(_06883_),
    .A(net7031),
    .B(net6931));
 sg13g2_nor2_1 _20465_ (.A(net7033),
    .B(_06883_),
    .Y(_06884_));
 sg13g2_nand3_1 _20466_ (.B(net7031),
    .C(net6932),
    .A(_02172_),
    .Y(_06885_));
 sg13g2_nor4_1 _20467_ (.A(_06834_),
    .B(_06841_),
    .C(_06882_),
    .D(_06885_),
    .Y(_06886_));
 sg13g2_nor4_1 _20468_ (.A(_06867_),
    .B(_06879_),
    .C(_06880_),
    .D(net6780),
    .Y(_06887_));
 sg13g2_nor2_1 _20469_ (.A(_06784_),
    .B(net6888),
    .Y(_06888_));
 sg13g2_nor2_1 _20470_ (.A(\cs_registers_i.debug_mode_i ),
    .B(_06888_),
    .Y(_06889_));
 sg13g2_nand2b_1 _20471_ (.Y(_06890_),
    .B(_06889_),
    .A_N(_06871_));
 sg13g2_nand2b_1 _20472_ (.Y(_06891_),
    .B(_00242_),
    .A_N(_02032_));
 sg13g2_a21o_1 _20473_ (.A2(_06891_),
    .A1(_06152_),
    .B1(_02105_),
    .X(_06892_));
 sg13g2_o21ai_1 _20474_ (.B1(_06892_),
    .Y(_06893_),
    .A1(_06152_),
    .A2(_06891_));
 sg13g2_nand2_1 _20475_ (.Y(_06894_),
    .A(net6930),
    .B(_06893_));
 sg13g2_nor2_1 _20476_ (.A(\id_stage_i.controller_i.store_err_q ),
    .B(\id_stage_i.controller_i.load_err_q ),
    .Y(_06895_));
 sg13g2_nor3_1 _20477_ (.A(\id_stage_i.controller_i.store_err_q ),
    .B(\id_stage_i.controller_i.load_err_q ),
    .C(\id_stage_i.controller_i.exc_req_q ),
    .Y(_06896_));
 sg13g2_nand2b_1 _20478_ (.Y(_06897_),
    .B(_06895_),
    .A_N(\id_stage_i.controller_i.exc_req_q ));
 sg13g2_and2_1 _20479_ (.A(\cs_registers_i.debug_ebreaku_o ),
    .B(_00243_),
    .X(_06898_));
 sg13g2_a22oi_1 _20480_ (.Y(_06899_),
    .B1(_06898_),
    .B2(_00242_),
    .A2(_06777_),
    .A1(\cs_registers_i.debug_ebreakm_o ));
 sg13g2_and2_1 _20481_ (.A(_02226_),
    .B(_06899_),
    .X(_06900_));
 sg13g2_nor2_1 _20482_ (.A(_08444_),
    .B(_10165_),
    .Y(_06901_));
 sg13g2_nand2_1 _20483_ (.Y(_06902_),
    .A(net7665),
    .B(\id_stage_i.controller_i.instr_fetch_err_i ));
 sg13g2_nor2_1 _20484_ (.A(\id_stage_i.controller_i.illegal_insn_q ),
    .B(_06901_),
    .Y(_06903_));
 sg13g2_nand3_1 _20485_ (.B(_06773_),
    .C(_06903_),
    .A(_06625_),
    .Y(_06904_));
 sg13g2_or4_1 _20486_ (.A(_10465_),
    .B(_06896_),
    .C(_06900_),
    .D(_06904_),
    .X(_06905_));
 sg13g2_nand4_1 _20487_ (.B(_06625_),
    .C(_06773_),
    .A(_10463_),
    .Y(_06906_),
    .D(_06903_));
 sg13g2_and2_1 _20488_ (.A(_01603_),
    .B(_06905_),
    .X(_06907_));
 sg13g2_nor2_1 _20489_ (.A(net349),
    .B(\cs_registers_i.debug_single_step_o ),
    .Y(_06908_));
 sg13g2_nor2b_1 _20490_ (.A(_06908_),
    .B_N(_01600_),
    .Y(_06909_));
 sg13g2_or2_1 _20491_ (.X(_06910_),
    .B(_01602_),
    .A(_01606_));
 sg13g2_nor4_1 _20492_ (.A(_01605_),
    .B(_06907_),
    .C(_06909_),
    .D(_06910_),
    .Y(_06911_));
 sg13g2_nor2_1 _20493_ (.A(net7477),
    .B(_06618_),
    .Y(_06912_));
 sg13g2_nor3_1 _20494_ (.A(_07655_),
    .B(_06599_),
    .C(_06912_),
    .Y(_06913_));
 sg13g2_and3_1 _20495_ (.X(_06914_),
    .A(net6932),
    .B(_06911_),
    .C(_06913_));
 sg13g2_nand2_1 _20496_ (.Y(_06915_),
    .A(_06884_),
    .B(_06914_));
 sg13g2_nand3_1 _20497_ (.B(_06894_),
    .C(_06915_),
    .A(_06890_),
    .Y(_06916_));
 sg13g2_inv_1 _20498_ (.Y(_06917_),
    .A(_06918_));
 sg13g2_nand2b_1 _20499_ (.Y(_06918_),
    .B(net7033),
    .A_N(_06834_));
 sg13g2_and3_1 _20500_ (.X(_06919_),
    .A(net7031),
    .B(_06848_),
    .C(_06917_));
 sg13g2_nor4_1 _20501_ (.A(_06859_),
    .B(_06862_),
    .C(_06883_),
    .D(_06918_),
    .Y(_06920_));
 sg13g2_nor2_1 _20502_ (.A(net6711),
    .B(_06920_),
    .Y(_06921_));
 sg13g2_or2_1 _20503_ (.X(_06922_),
    .B(_06869_),
    .A(net6949));
 sg13g2_or2_1 _20504_ (.X(_06923_),
    .B(_06922_),
    .A(_06870_));
 sg13g2_nor2_1 _20505_ (.A(net6948),
    .B(_06836_),
    .Y(_06924_));
 sg13g2_nand3_1 _20506_ (.B(net7033),
    .C(_06835_),
    .A(_13838_),
    .Y(_06925_));
 sg13g2_o21ai_1 _20507_ (.B1(_06923_),
    .Y(_06926_),
    .A1(_06842_),
    .A2(_06925_));
 sg13g2_nand2_1 _20508_ (.Y(_06927_),
    .A(_06868_),
    .B(_06926_));
 sg13g2_a221oi_1 _20509_ (.B2(net6950),
    .C1(_06806_),
    .B1(_06857_),
    .A1(_06784_),
    .Y(_06928_),
    .A2(_06791_));
 sg13g2_or4_1 _20510_ (.A(_09944_),
    .B(_13838_),
    .C(_06789_),
    .D(_06817_),
    .X(_06929_));
 sg13g2_o21ai_1 _20511_ (.B1(_06929_),
    .Y(_06930_),
    .A1(_06792_),
    .A2(_06922_));
 sg13g2_or4_1 _20512_ (.A(net6975),
    .B(net6900),
    .C(net6887),
    .D(_06834_),
    .X(_06931_));
 sg13g2_nor4_1 _20513_ (.A(_06810_),
    .B(_06842_),
    .C(_06885_),
    .D(_06931_),
    .Y(_06932_));
 sg13g2_a221oi_1 _20514_ (.B2(_06874_),
    .C1(_06932_),
    .B1(_06930_),
    .A1(_06924_),
    .Y(_06933_),
    .A2(_06928_));
 sg13g2_nand3_1 _20515_ (.B(_06927_),
    .C(_06933_),
    .A(_06921_),
    .Y(_06934_));
 sg13g2_nor2_1 _20516_ (.A(_06837_),
    .B(_06934_),
    .Y(_06935_));
 sg13g2_nor3_1 _20517_ (.A(\cs_registers_i.debug_mode_i ),
    .B(_06888_),
    .C(_06923_),
    .Y(_06936_));
 sg13g2_nand3_1 _20518_ (.B(_06911_),
    .C(_06913_),
    .A(_06786_),
    .Y(_06937_));
 sg13g2_o21ai_1 _20519_ (.B1(_06894_),
    .Y(_06938_),
    .A1(_06885_),
    .A2(_06937_));
 sg13g2_or2_1 _20520_ (.X(_06939_),
    .B(_06938_),
    .A(_06936_));
 sg13g2_nor4_1 _20521_ (.A(_06859_),
    .B(_06862_),
    .C(_06883_),
    .D(_06918_),
    .Y(_06940_));
 sg13g2_or2_1 _20522_ (.X(_06941_),
    .B(_06940_),
    .A(_06919_));
 sg13g2_nor3_1 _20523_ (.A(_02172_),
    .B(net7031),
    .C(_06834_),
    .Y(_06942_));
 sg13g2_or4_1 _20524_ (.A(net6975),
    .B(net6900),
    .C(_06810_),
    .D(net6887),
    .X(_06943_));
 sg13g2_nor4_1 _20525_ (.A(_06834_),
    .B(_06842_),
    .C(_06885_),
    .D(_06943_),
    .Y(_06944_));
 sg13g2_inv_1 _20526_ (.Y(_06945_),
    .A(_06946_));
 sg13g2_nand2_1 _20527_ (.Y(_06946_),
    .A(_13838_),
    .B(_06942_));
 sg13g2_a21oi_1 _20528_ (.A1(_06928_),
    .A2(_06945_),
    .Y(_06947_),
    .B1(net6824));
 sg13g2_or3_1 _20529_ (.A(net7033),
    .B(net7031),
    .C(_06834_),
    .X(_06948_));
 sg13g2_or4_1 _20530_ (.A(_09944_),
    .B(_13838_),
    .C(_06789_),
    .D(_06817_),
    .X(_06949_));
 sg13g2_o21ai_1 _20531_ (.B1(_06949_),
    .Y(_06950_),
    .A1(_06792_),
    .A2(_06922_));
 sg13g2_nand2b_1 _20532_ (.Y(_06951_),
    .B(_06950_),
    .A_N(_06948_));
 sg13g2_o21ai_1 _20533_ (.B1(_06947_),
    .Y(_06952_),
    .A1(_06785_),
    .A2(_06951_));
 sg13g2_inv_1 _20534_ (.Y(_06953_),
    .A(_06954_));
 sg13g2_or2_1 _20535_ (.X(_06954_),
    .B(_06948_),
    .A(_06922_));
 sg13g2_o21ai_1 _20536_ (.B1(_06954_),
    .Y(_06955_),
    .A1(_06842_),
    .A2(_06946_));
 sg13g2_a221oi_1 _20537_ (.B2(_06868_),
    .C1(_06952_),
    .B1(_06955_),
    .A1(_06831_),
    .Y(_06956_),
    .A2(_06942_));
 sg13g2_nand2b_1 _20538_ (.Y(_06957_),
    .B(_06956_),
    .A_N(_06941_));
 sg13g2_o21ai_1 _20539_ (.B1(_06771_),
    .Y(_06958_),
    .A1(_06935_),
    .A2(_06939_));
 sg13g2_nor3_1 _20540_ (.A(net7657),
    .B(net7659),
    .C(_01983_),
    .Y(_06959_));
 sg13g2_inv_1 _20541_ (.Y(_06960_),
    .A(_06961_));
 sg13g2_nand2_1 _20542_ (.Y(_06961_),
    .A(net348),
    .B(_06959_));
 sg13g2_nor2_1 _20543_ (.A(net314),
    .B(\load_store_unit_i.lsu_err_q ),
    .Y(_06962_));
 sg13g2_nor2_1 _20544_ (.A(_06961_),
    .B(_06962_),
    .Y(_06963_));
 sg13g2_or2_1 _20545_ (.X(_06964_),
    .B(_06962_),
    .A(_06961_));
 sg13g2_or2_1 _20546_ (.X(_06965_),
    .B(_06778_),
    .A(_06775_));
 sg13g2_nor2_1 _20547_ (.A(_06779_),
    .B(_06965_),
    .Y(_06966_));
 sg13g2_and3_1 _20548_ (.X(_06967_),
    .A(net7927),
    .B(_03638_),
    .C(_06618_));
 sg13g2_nand3_1 _20549_ (.B(_03638_),
    .C(_06618_),
    .A(net7927),
    .Y(_06968_));
 sg13g2_nor2_1 _20550_ (.A(_09324_),
    .B(_06968_),
    .Y(_06969_));
 sg13g2_nand2_1 _20551_ (.Y(_06970_),
    .A(net7930),
    .B(_06967_));
 sg13g2_nor3_1 _20552_ (.A(net7699),
    .B(_06635_),
    .C(_06970_),
    .Y(_06971_));
 sg13g2_nor4_1 _20553_ (.A(net7734),
    .B(net7748),
    .C(_06632_),
    .D(_06969_),
    .Y(_06972_));
 sg13g2_nor2_1 _20554_ (.A(_06971_),
    .B(_06972_),
    .Y(_06973_));
 sg13g2_nand2_1 _20555_ (.Y(_06974_),
    .A(net7665),
    .B(net7680));
 sg13g2_nor4_1 _20556_ (.A(_06627_),
    .B(_06937_),
    .C(_06973_),
    .D(_06974_),
    .Y(_06975_));
 sg13g2_nor4_1 _20557_ (.A(_06779_),
    .B(_06963_),
    .C(_06965_),
    .D(_06975_),
    .Y(_06976_));
 sg13g2_a21oi_1 _20558_ (.A1(net7665),
    .A2(\cs_registers_i.debug_single_step_o ),
    .Y(_06977_),
    .B1(net349));
 sg13g2_nor2_1 _20559_ (.A(net7984),
    .B(_06977_),
    .Y(_06978_));
 sg13g2_or2_1 _20560_ (.X(_06979_),
    .B(_06977_),
    .A(net7984));
 sg13g2_a21oi_1 _20561_ (.A1(net436),
    .A2(_00389_),
    .Y(_06980_),
    .B1(net434));
 sg13g2_a22oi_1 _20562_ (.Y(_06981_),
    .B1(_00396_),
    .B2(net430),
    .A2(_00397_),
    .A1(net431));
 sg13g2_a22oi_1 _20563_ (.Y(_06982_),
    .B1(_00394_),
    .B2(net428),
    .A2(_00395_),
    .A1(net429));
 sg13g2_inv_1 _20564_ (.Y(_06983_),
    .A(_06982_));
 sg13g2_and2_1 _20565_ (.A(_06981_),
    .B(_06982_),
    .X(_06984_));
 sg13g2_nand2_1 _20566_ (.Y(_06985_),
    .A(net426),
    .B(_00392_));
 sg13g2_nand2_1 _20567_ (.Y(_06986_),
    .A(net427),
    .B(_00393_));
 sg13g2_and2_1 _20568_ (.A(_06985_),
    .B(_06986_),
    .X(_06987_));
 sg13g2_a22oi_1 _20569_ (.Y(_06988_),
    .B1(_00382_),
    .B2(net419),
    .A2(_00391_),
    .A1(net425));
 sg13g2_nand3_1 _20570_ (.B(_06987_),
    .C(_06988_),
    .A(_06984_),
    .Y(_06989_));
 sg13g2_a22oi_1 _20571_ (.Y(_06990_),
    .B1(_00398_),
    .B2(net432),
    .A2(_00399_),
    .A1(net433));
 sg13g2_nand2_1 _20572_ (.Y(_06991_),
    .A(net420),
    .B(_00383_));
 sg13g2_a22oi_1 _20573_ (.Y(_06992_),
    .B1(_00383_),
    .B2(net420),
    .A2(_00384_),
    .A1(net421));
 sg13g2_nand2_1 _20574_ (.Y(_06993_),
    .A(_06990_),
    .B(_06992_));
 sg13g2_inv_1 _20575_ (.Y(_06994_),
    .A(_06995_));
 sg13g2_nand2_1 _20576_ (.Y(_06995_),
    .A(net424),
    .B(_00387_));
 sg13g2_a22oi_1 _20577_ (.Y(_06996_),
    .B1(_00385_),
    .B2(net422),
    .A2(_00386_),
    .A1(net423));
 sg13g2_nand2_1 _20578_ (.Y(_06997_),
    .A(_06995_),
    .B(_06996_));
 sg13g2_nor3_1 _20579_ (.A(_06989_),
    .B(_06993_),
    .C(_06997_),
    .Y(_06998_));
 sg13g2_nand2_1 _20580_ (.Y(_06999_),
    .A(net418),
    .B(_00388_));
 sg13g2_a22oi_1 _20581_ (.Y(_07000_),
    .B1(_00388_),
    .B2(net418),
    .A2(_00390_),
    .A1(net435));
 sg13g2_and2_1 _20582_ (.A(_06998_),
    .B(_07000_),
    .X(_07001_));
 sg13g2_nand2_1 _20583_ (.Y(_07002_),
    .A(_06980_),
    .B(_07001_));
 sg13g2_o21ai_1 _20584_ (.B1(_07002_),
    .Y(_07003_),
    .A1(net434),
    .A2(\cs_registers_i.csr_mstatus_mie_o ));
 sg13g2_nor3_1 _20585_ (.A(\cs_registers_i.nmi_mode_i ),
    .B(\cs_registers_i.debug_mode_i ),
    .C(_07003_),
    .Y(_07004_));
 sg13g2_nor2_1 _20586_ (.A(_06978_),
    .B(_07004_),
    .Y(_07005_));
 sg13g2_nand2_1 _20587_ (.Y(_07006_),
    .A(net417),
    .B(net7937));
 sg13g2_nor2_1 _20588_ (.A(_01673_),
    .B(_07006_),
    .Y(_07007_));
 sg13g2_a21oi_1 _20589_ (.A1(_01835_),
    .A2(_07007_),
    .Y(_07008_),
    .B1(_01836_));
 sg13g2_a21oi_1 _20590_ (.A1(_01747_),
    .A2(_01746_),
    .Y(_07009_),
    .B1(_01705_));
 sg13g2_a21oi_1 _20591_ (.A1(net392),
    .A2(net393),
    .Y(_07010_),
    .B1(net383));
 sg13g2_nor2b_1 _20592_ (.A(net7966),
    .B_N(_07010_),
    .Y(_07011_));
 sg13g2_a21oi_1 _20593_ (.A1(net7966),
    .A2(_07009_),
    .Y(_07012_),
    .B1(_07011_));
 sg13g2_nand2_1 _20594_ (.Y(_07013_),
    .A(net7976),
    .B(_07012_));
 sg13g2_nor2_1 _20595_ (.A(_01835_),
    .B(_07007_),
    .Y(_07014_));
 sg13g2_mux2_1 _20596_ (.A0(_07008_),
    .A1(_07014_),
    .S(_07013_),
    .X(_07015_));
 sg13g2_nand3_1 _20597_ (.B(_06958_),
    .C(_06976_),
    .A(_06783_),
    .Y(_07016_));
 sg13g2_nor2_1 _20598_ (.A(_02232_),
    .B(_07016_),
    .Y(_07017_));
 sg13g2_o21ai_1 _20599_ (.B1(_02245_),
    .Y(_07018_),
    .A1(_02232_),
    .A2(_07016_));
 sg13g2_nor2b_1 _20600_ (.A(_07005_),
    .B_N(_07018_),
    .Y(_07019_));
 sg13g2_or2_1 _20601_ (.X(_07020_),
    .B(_07019_),
    .A(_07015_));
 sg13g2_and2_1 _20602_ (.A(\id_stage_i.controller_i.controller_run_o ),
    .B(_07016_),
    .X(_07021_));
 sg13g2_nor2_1 _20603_ (.A(net7985),
    .B(_06910_),
    .Y(_07022_));
 sg13g2_inv_1 _20604_ (.Y(_07023_),
    .A(_07022_));
 sg13g2_a21o_1 _20605_ (.A2(_08669_),
    .A1(net7608),
    .B1(_08648_),
    .X(_07024_));
 sg13g2_o21ai_1 _20606_ (.B1(net7981),
    .Y(_07025_),
    .A1(_07595_),
    .A2(net7377));
 sg13g2_inv_1 _20607_ (.Y(_07026_),
    .A(\alu_adder_result_ex[0] ));
 sg13g2_a21oi_1 _20608_ (.A1(_07024_),
    .A2(_07025_),
    .Y(_07027_),
    .B1(_06599_));
 sg13g2_nor2_1 _20609_ (.A(_05195_),
    .B(_07792_),
    .Y(_07028_));
 sg13g2_nor3_1 _20610_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_valid ),
    .B(net8016),
    .C(_07028_),
    .Y(_07029_));
 sg13g2_and2_1 _20611_ (.A(_08239_),
    .B(_07029_),
    .X(_07030_));
 sg13g2_nand2_1 _20612_ (.Y(_07031_),
    .A(_08239_),
    .B(_07029_));
 sg13g2_nand3_1 _20613_ (.B(_06598_),
    .C(_07030_),
    .A(_02201_),
    .Y(_07032_));
 sg13g2_a21oi_1 _20614_ (.A1(_08696_),
    .A2(_07032_),
    .Y(_07033_),
    .B1(_08444_));
 sg13g2_o21ai_1 _20615_ (.B1(_06641_),
    .Y(_07034_),
    .A1(_07027_),
    .A2(_07033_));
 sg13g2_nand2_1 _20616_ (.Y(_07035_),
    .A(_08696_),
    .B(_07031_));
 sg13g2_and2_1 _20617_ (.A(_07027_),
    .B(_07030_),
    .X(_07036_));
 sg13g2_o21ai_1 _20618_ (.B1(_07035_),
    .Y(_07037_),
    .A1(_06961_),
    .A2(_07036_));
 sg13g2_a21o_1 _20619_ (.A2(_07037_),
    .A1(net7981),
    .B1(_07034_),
    .X(_07038_));
 sg13g2_nor2_1 _20620_ (.A(_07599_),
    .B(net6056),
    .Y(_07039_));
 sg13g2_nor4_1 _20621_ (.A(net7981),
    .B(_07599_),
    .C(net6056),
    .D(_06768_),
    .Y(_07040_));
 sg13g2_inv_1 _20622_ (.Y(_07041_),
    .A(net5968));
 sg13g2_o21ai_1 _20623_ (.B1(_07038_),
    .Y(_07042_),
    .A1(_06766_),
    .A2(_06769_));
 sg13g2_nor3_1 _20624_ (.A(_07021_),
    .B(_07023_),
    .C(net5968),
    .Y(_07043_));
 sg13g2_nor4_2 _20625_ (.A(_07042_),
    .B(_07021_),
    .C(_07023_),
    .Y(_07044_),
    .D(_07020_));
 sg13g2_inv_1 _20626_ (.Y(_07045_),
    .A(_07044_));
 sg13g2_mux2_1 _20627_ (.A0(_01948_),
    .A1(_01738_),
    .S(net5935),
    .X(_07046_));
 sg13g2_mux2_1 _20628_ (.A0(_01947_),
    .A1(_01737_),
    .S(net5934),
    .X(_07047_));
 sg13g2_nand2_1 _20629_ (.Y(_07048_),
    .A(net5939),
    .B(_01736_));
 sg13g2_o21ai_1 _20630_ (.B1(_07048_),
    .Y(_07049_),
    .A1(_07450_),
    .A2(net5934));
 sg13g2_mux2_1 _20631_ (.A0(_01945_),
    .A1(_01735_),
    .S(net5939),
    .X(_07050_));
 sg13g2_mux2_1 _20632_ (.A0(_01944_),
    .A1(_01734_),
    .S(net5937),
    .X(_07051_));
 sg13g2_mux2_1 _20633_ (.A0(_01943_),
    .A1(_01733_),
    .S(net5941),
    .X(_07052_));
 sg13g2_nand2_1 _20634_ (.Y(_07053_),
    .A(net5941),
    .B(_01732_));
 sg13g2_o21ai_1 _20635_ (.B1(_07053_),
    .Y(_07054_),
    .A1(_07622_),
    .A2(net5941));
 sg13g2_mux2_1 _20636_ (.A0(_01941_),
    .A1(_01731_),
    .S(net5938),
    .X(_07055_));
 sg13g2_mux2_1 _20637_ (.A0(_01940_),
    .A1(_01730_),
    .S(net5938),
    .X(_07056_));
 sg13g2_mux2_1 _20638_ (.A0(_01939_),
    .A1(_01729_),
    .S(net5941),
    .X(_07057_));
 sg13g2_mux2_1 _20639_ (.A0(_01938_),
    .A1(_01728_),
    .S(net5938),
    .X(_07058_));
 sg13g2_mux2_1 _20640_ (.A0(_01937_),
    .A1(_01727_),
    .S(net5938),
    .X(_07059_));
 sg13g2_mux2_1 _20641_ (.A0(_01936_),
    .A1(_01726_),
    .S(net5936),
    .X(_07060_));
 sg13g2_mux2_1 _20642_ (.A0(_01935_),
    .A1(_01725_),
    .S(net5936),
    .X(_07061_));
 sg13g2_mux2_1 _20643_ (.A0(_01934_),
    .A1(_01724_),
    .S(net5936),
    .X(_07062_));
 sg13g2_mux2_1 _20644_ (.A0(_01933_),
    .A1(_01723_),
    .S(net5936),
    .X(_07063_));
 sg13g2_mux2_1 _20645_ (.A0(_01932_),
    .A1(_01722_),
    .S(net5937),
    .X(_07064_));
 sg13g2_mux2_1 _20646_ (.A0(_01931_),
    .A1(_01721_),
    .S(net5937),
    .X(_07065_));
 sg13g2_mux2_1 _20647_ (.A0(_01930_),
    .A1(_01720_),
    .S(net5937),
    .X(_07066_));
 sg13g2_mux2_1 _20648_ (.A0(_01929_),
    .A1(_01719_),
    .S(net5937),
    .X(_07067_));
 sg13g2_mux2_1 _20649_ (.A0(_01928_),
    .A1(_01718_),
    .S(net5941),
    .X(_07068_));
 sg13g2_mux2_1 _20650_ (.A0(_01927_),
    .A1(_01717_),
    .S(net5936),
    .X(_07069_));
 sg13g2_nand2_1 _20651_ (.Y(_07070_),
    .A(net5936),
    .B(_01716_));
 sg13g2_o21ai_1 _20652_ (.B1(_07070_),
    .Y(_07071_),
    .A1(_08227_),
    .A2(net5936));
 sg13g2_mux2_1 _20653_ (.A0(_01925_),
    .A1(_01715_),
    .S(net5939),
    .X(_07072_));
 sg13g2_mux2_1 _20654_ (.A0(_01924_),
    .A1(_01714_),
    .S(net5936),
    .X(_07073_));
 sg13g2_mux2_1 _20655_ (.A0(_01923_),
    .A1(_01713_),
    .S(net5935),
    .X(_07074_));
 sg13g2_mux2_1 _20656_ (.A0(_01922_),
    .A1(_01712_),
    .S(net5937),
    .X(_07075_));
 sg13g2_mux2_1 _20657_ (.A0(_01921_),
    .A1(_01711_),
    .S(net5935),
    .X(_07076_));
 sg13g2_mux2_1 _20658_ (.A0(_01920_),
    .A1(_01710_),
    .S(net5937),
    .X(_07077_));
 sg13g2_mux2_1 _20659_ (.A0(_01919_),
    .A1(_01709_),
    .S(net5935),
    .X(_07078_));
 sg13g2_nand2_1 _20660_ (.Y(_07079_),
    .A(net5934),
    .B(_01708_));
 sg13g2_o21ai_1 _20661_ (.B1(_07079_),
    .Y(_07080_),
    .A1(_08414_),
    .A2(net5934));
 sg13g2_nor3_1 _20662_ (.A(net7981),
    .B(_06599_),
    .C(_07024_),
    .Y(_07081_));
 sg13g2_a21oi_1 _20663_ (.A1(_06641_),
    .A2(_07081_),
    .Y(_07082_),
    .B1(\id_stage_i.branch_set ));
 sg13g2_nor3_1 _20664_ (.A(_02232_),
    .B(_06901_),
    .C(_07082_),
    .Y(_07083_));
 sg13g2_nor2_1 _20665_ (.A(_06897_),
    .B(_06965_),
    .Y(_07084_));
 sg13g2_nor2_1 _20666_ (.A(_02238_),
    .B(_07084_),
    .Y(_07085_));
 sg13g2_nand2_1 _20667_ (.Y(_07086_),
    .A(_06905_),
    .B(_07085_));
 sg13g2_and2_1 _20668_ (.A(\id_stage_i.controller_i.nmi_mode_d ),
    .B(_07004_),
    .X(_07087_));
 sg13g2_nand2_1 _20669_ (.Y(_07088_),
    .A(\id_stage_i.controller_i.nmi_mode_d ),
    .B(_07004_));
 sg13g2_nand2b_1 _20670_ (.Y(_07089_),
    .B(_07088_),
    .A_N(_06909_));
 sg13g2_nand2b_1 _20671_ (.Y(_07090_),
    .B(_07086_),
    .A_N(_07089_));
 sg13g2_nand2b_1 _20672_ (.Y(_07091_),
    .B(_00006_),
    .A_N(_01604_));
 sg13g2_nor4_1 _20673_ (.A(_01605_),
    .B(_07083_),
    .C(_07090_),
    .D(_07091_),
    .Y(_07092_));
 sg13g2_or4_1 _20674_ (.A(_01605_),
    .B(_07083_),
    .C(_07090_),
    .D(_07091_),
    .X(_07093_));
 sg13g2_and2_1 _20675_ (.A(net7665),
    .B(_06911_),
    .X(_07094_));
 sg13g2_o21ai_1 _20676_ (.B1(_07094_),
    .Y(_07095_),
    .A1(_07021_),
    .A2(net5968));
 sg13g2_o21ai_1 _20677_ (.B1(_07095_),
    .Y(_07096_),
    .A1(_07045_),
    .A2(_07093_));
 sg13g2_nor2_1 _20678_ (.A(net7666),
    .B(net5946),
    .Y(_07097_));
 sg13g2_mux2_1 _20679_ (.A0(net396),
    .A1(net393),
    .S(net7967),
    .X(_07098_));
 sg13g2_nor2_1 _20680_ (.A(net7957),
    .B(_07098_),
    .Y(_07099_));
 sg13g2_nand2b_1 _20681_ (.Y(_07100_),
    .B(net7968),
    .A_N(_01747_));
 sg13g2_o21ai_1 _20682_ (.B1(_07100_),
    .Y(_07101_),
    .A1(_01750_),
    .A2(net7968));
 sg13g2_a21oi_1 _20683_ (.A1(net7957),
    .A2(_07101_),
    .Y(_07102_),
    .B1(_07099_));
 sg13g2_a21o_1 _20684_ (.A2(_07101_),
    .A1(net7957),
    .B1(_07099_),
    .X(_07103_));
 sg13g2_mux2_1 _20685_ (.A0(net389),
    .A1(net406),
    .S(net7967),
    .X(_07104_));
 sg13g2_nor2_1 _20686_ (.A(net7958),
    .B(_07104_),
    .Y(_07105_));
 sg13g2_nand2b_1 _20687_ (.Y(_07106_),
    .B(net7967),
    .A_N(_01760_));
 sg13g2_o21ai_1 _20688_ (.B1(_07106_),
    .Y(_07107_),
    .A1(_01743_),
    .A2(net7967));
 sg13g2_a21oi_1 _20689_ (.A1(net7965),
    .A2(_07107_),
    .Y(_07108_),
    .B1(_07105_));
 sg13g2_a21o_1 _20690_ (.A2(_07107_),
    .A1(net7965),
    .B1(_07105_),
    .X(_07109_));
 sg13g2_mux2_1 _20691_ (.A0(net391),
    .A1(net409),
    .S(net7974),
    .X(_07110_));
 sg13g2_nor2_1 _20692_ (.A(net7963),
    .B(_07110_),
    .Y(_07111_));
 sg13g2_nand2b_1 _20693_ (.Y(_07112_),
    .B(net7970),
    .A_N(_01763_));
 sg13g2_o21ai_1 _20694_ (.B1(_07112_),
    .Y(_07113_),
    .A1(_01745_),
    .A2(net7970));
 sg13g2_a21oi_1 _20695_ (.A1(net7959),
    .A2(_07113_),
    .Y(_07114_),
    .B1(_07111_));
 sg13g2_a21o_1 _20696_ (.A2(_07113_),
    .A1(net7959),
    .B1(_07111_),
    .X(_07115_));
 sg13g2_nor2_1 _20697_ (.A(net7407),
    .B(net7403),
    .Y(_07116_));
 sg13g2_mux2_1 _20698_ (.A0(net385),
    .A1(net392),
    .S(net7968),
    .X(_07117_));
 sg13g2_nor2_1 _20699_ (.A(net7957),
    .B(_07117_),
    .Y(_07118_));
 sg13g2_nand2b_1 _20700_ (.Y(_07119_),
    .B(net7976),
    .A_N(_01746_));
 sg13g2_o21ai_1 _20701_ (.B1(_07119_),
    .Y(_07120_),
    .A1(_01739_),
    .A2(net7976));
 sg13g2_a21oi_1 _20702_ (.A1(net7966),
    .A2(_07120_),
    .Y(_07121_),
    .B1(_07118_));
 sg13g2_a21o_1 _20703_ (.A2(_07120_),
    .A1(net7966),
    .B1(_07118_),
    .X(_07122_));
 sg13g2_mux4_1 _20704_ (.S0(net7972),
    .A0(net411),
    .A1(net397),
    .A2(_01783_),
    .A3(_01751_),
    .S1(net7961),
    .X(_07123_));
 sg13g2_mux2_1 _20705_ (.A0(net390),
    .A1(net408),
    .S(net7975),
    .X(_07124_));
 sg13g2_nor2_1 _20706_ (.A(net7964),
    .B(_07124_),
    .Y(_07125_));
 sg13g2_nand2b_1 _20707_ (.Y(_07126_),
    .B(net7975),
    .A_N(_01762_));
 sg13g2_o21ai_1 _20708_ (.B1(_07126_),
    .Y(_07127_),
    .A1(_01744_),
    .A2(net7969));
 sg13g2_a21oi_1 _20709_ (.A1(net7959),
    .A2(_07127_),
    .Y(_07128_),
    .B1(_07125_));
 sg13g2_a21o_1 _20710_ (.A2(_07127_),
    .A1(net7959),
    .B1(_07125_),
    .X(_07129_));
 sg13g2_nor2_1 _20711_ (.A(net7400),
    .B(_07129_),
    .Y(_07130_));
 sg13g2_nand2_1 _20712_ (.Y(_07131_),
    .A(net7401),
    .B(_07128_));
 sg13g2_mux4_1 _20713_ (.S0(net7973),
    .A0(net413),
    .A1(net399),
    .A2(_01805_),
    .A3(_01753_),
    .S1(net7963),
    .X(_07132_));
 sg13g2_nor2_1 _20714_ (.A(net7408),
    .B(_07121_),
    .Y(_07133_));
 sg13g2_nand2_1 _20715_ (.Y(_07134_),
    .A(net7404),
    .B(_07122_));
 sg13g2_nand2_1 _20716_ (.Y(_07135_),
    .A(net7400),
    .B(_07123_));
 sg13g2_a22oi_1 _20717_ (.Y(_07136_),
    .B1(net7308),
    .B2(net7620),
    .A2(net7621),
    .A1(net7399));
 sg13g2_nand3_1 _20718_ (.B(net7621),
    .C(net7308),
    .A(net7395),
    .Y(_07137_));
 sg13g2_o21ai_1 _20719_ (.B1(_07137_),
    .Y(_07138_),
    .A1(net7306),
    .A2(_07136_));
 sg13g2_nor2_1 _20720_ (.A(net7409),
    .B(net7397),
    .Y(_07139_));
 sg13g2_mux4_1 _20721_ (.S0(net7972),
    .A0(net407),
    .A1(net394),
    .A2(_01761_),
    .A3(_01748_),
    .S1(net7961),
    .X(_07140_));
 sg13g2_mux4_1 _20722_ (.S0(net7973),
    .A0(net412),
    .A1(net398),
    .A2(_01794_),
    .A3(_01752_),
    .S1(net7963),
    .X(_07141_));
 sg13g2_inv_1 _20723_ (.Y(_07142_),
    .A(net7618));
 sg13g2_or2_1 _20724_ (.X(_07143_),
    .B(_07141_),
    .A(_07132_));
 sg13g2_mux4_1 _20725_ (.S0(net7969),
    .A0(net410),
    .A1(net395),
    .A2(_01772_),
    .A3(_01749_),
    .S1(net7960),
    .X(_07144_));
 sg13g2_nor3_1 _20726_ (.A(_07123_),
    .B(_07143_),
    .C(_07144_),
    .Y(_07145_));
 sg13g2_nor2b_1 _20727_ (.A(_07140_),
    .B_N(_07145_),
    .Y(_07146_));
 sg13g2_nor2_1 _20728_ (.A(_07108_),
    .B(net7394),
    .Y(_07147_));
 sg13g2_nand2_1 _20729_ (.Y(_07148_),
    .A(_07109_),
    .B(net7391));
 sg13g2_nor2_1 _20730_ (.A(net7399),
    .B(_07148_),
    .Y(_07149_));
 sg13g2_nand2_1 _20731_ (.Y(_07150_),
    .A(net7402),
    .B(_07147_));
 sg13g2_and2_1 _20732_ (.A(_07146_),
    .B(_07149_),
    .X(_07151_));
 sg13g2_inv_1 _20733_ (.Y(_07152_),
    .A(net6568));
 sg13g2_and2_1 _20734_ (.A(_07139_),
    .B(_07151_),
    .X(_07153_));
 sg13g2_mux4_1 _20735_ (.S0(net7967),
    .A0(net416),
    .A1(net402),
    .A2(_01834_),
    .A3(_01756_),
    .S1(net7958),
    .X(_07154_));
 sg13g2_nand2_1 _20736_ (.Y(_07155_),
    .A(net7397),
    .B(_07128_));
 sg13g2_nor2_1 _20737_ (.A(_07114_),
    .B(_07129_),
    .Y(_07156_));
 sg13g2_nor2_1 _20738_ (.A(net7401),
    .B(_07122_),
    .Y(_07157_));
 sg13g2_nand2_1 _20739_ (.Y(_07158_),
    .A(net7395),
    .B(_07156_));
 sg13g2_nor2_1 _20740_ (.A(net7404),
    .B(net7396),
    .Y(_07159_));
 sg13g2_nor2_1 _20741_ (.A(net7399),
    .B(net7394),
    .Y(_07160_));
 sg13g2_o21ai_1 _20742_ (.B1(_07147_),
    .Y(_07161_),
    .A1(net7401),
    .A2(net7395));
 sg13g2_nand2_1 _20743_ (.Y(_07162_),
    .A(_07158_),
    .B(_07161_));
 sg13g2_nor3_1 _20744_ (.A(net7413),
    .B(_07159_),
    .C(_07162_),
    .Y(_07163_));
 sg13g2_nor2_1 _20745_ (.A(_07153_),
    .B(_07163_),
    .Y(_07164_));
 sg13g2_a22oi_1 _20746_ (.Y(_07165_),
    .B1(net7616),
    .B2(_07164_),
    .A2(_07138_),
    .A1(net7409));
 sg13g2_a21oi_1 _20747_ (.A1(net5947),
    .A2(_07165_),
    .Y(_07166_),
    .B1(_07097_));
 sg13g2_nor2_1 _20748_ (.A(net7671),
    .B(net5946),
    .Y(_07167_));
 sg13g2_mux4_1 _20749_ (.S0(net7971),
    .A0(net415),
    .A1(net401),
    .A2(_01827_),
    .A3(_01755_),
    .S1(net7962),
    .X(_07168_));
 sg13g2_nor2_1 _20750_ (.A(net7408),
    .B(net7399),
    .Y(_07169_));
 sg13g2_o21ai_1 _20751_ (.B1(_07169_),
    .Y(_07170_),
    .A1(net7393),
    .A2(_07146_));
 sg13g2_nand2_1 _20752_ (.Y(_07171_),
    .A(_07139_),
    .B(_07170_));
 sg13g2_nand2_1 _20753_ (.Y(_07172_),
    .A(net7412),
    .B(net7395));
 sg13g2_nor2_1 _20754_ (.A(_07102_),
    .B(_07121_),
    .Y(_07173_));
 sg13g2_o21ai_1 _20755_ (.B1(_07109_),
    .Y(_07174_),
    .A1(_07115_),
    .A2(_07128_));
 sg13g2_and2_1 _20756_ (.A(_07173_),
    .B(_07174_),
    .X(_07175_));
 sg13g2_nand2_1 _20757_ (.Y(_07176_),
    .A(_07173_),
    .B(_07174_));
 sg13g2_nand2_1 _20758_ (.Y(_07177_),
    .A(_07172_),
    .B(_07176_));
 sg13g2_nor2_1 _20759_ (.A(_07102_),
    .B(_07122_),
    .Y(_07178_));
 sg13g2_nand2_1 _20760_ (.Y(_07179_),
    .A(_07103_),
    .B(net7397));
 sg13g2_nor2_1 _20761_ (.A(net7405),
    .B(net7394),
    .Y(_07180_));
 sg13g2_or2_1 _20762_ (.X(_07181_),
    .B(_07180_),
    .A(_07130_));
 sg13g2_or2_1 _20763_ (.X(_07182_),
    .B(_07181_),
    .A(net7302));
 sg13g2_nand4_1 _20764_ (.B(_07172_),
    .C(_07176_),
    .A(_07171_),
    .Y(_07183_),
    .D(_07182_));
 sg13g2_and2_1 _20765_ (.A(_07116_),
    .B(_07173_),
    .X(_07184_));
 sg13g2_a21o_1 _20766_ (.A2(net7305),
    .A1(net7308),
    .B1(_07184_),
    .X(_07185_));
 sg13g2_a22oi_1 _20767_ (.Y(_07186_),
    .B1(_07185_),
    .B2(net7617),
    .A2(_07183_),
    .A1(net7614));
 sg13g2_a21oi_1 _20768_ (.A1(net5946),
    .A2(_07186_),
    .Y(_07187_),
    .B1(_07167_));
 sg13g2_mux4_1 _20769_ (.S0(net7971),
    .A0(net414),
    .A1(net400),
    .A2(_01816_),
    .A3(_01754_),
    .S1(net7962),
    .X(_07188_));
 sg13g2_mux2_1 _20770_ (.A0(net7399),
    .A1(net7613),
    .S(net7405),
    .X(_07189_));
 sg13g2_mux2_1 _20771_ (.A0(net388),
    .A1(net405),
    .S(net7975),
    .X(_07190_));
 sg13g2_nor2_1 _20772_ (.A(net7960),
    .B(_07190_),
    .Y(_07191_));
 sg13g2_nand2b_1 _20773_ (.Y(_07192_),
    .B(net7969),
    .A_N(_01759_));
 sg13g2_o21ai_1 _20774_ (.B1(_07192_),
    .Y(_07193_),
    .A1(_01742_),
    .A2(net7969));
 sg13g2_a21oi_1 _20775_ (.A1(net7959),
    .A2(_07193_),
    .Y(_07194_),
    .B1(_07191_));
 sg13g2_a21o_1 _20776_ (.A2(_07193_),
    .A1(net7959),
    .B1(_07191_),
    .X(_07195_));
 sg13g2_a221oi_1 _20777_ (.B2(net7308),
    .C1(net7413),
    .B1(net7389),
    .A1(net7391),
    .Y(_07196_),
    .A2(_07189_));
 sg13g2_a21oi_1 _20778_ (.A1(_07156_),
    .A2(net7305),
    .Y(_07197_),
    .B1(_07175_));
 sg13g2_nand2b_1 _20779_ (.Y(_07198_),
    .B(net7613),
    .A_N(_07197_));
 sg13g2_o21ai_1 _20780_ (.B1(_07198_),
    .Y(_07199_),
    .A1(_07122_),
    .A2(_07196_));
 sg13g2_mux4_1 _20781_ (.S0(net7974),
    .A0(net386),
    .A1(net403),
    .A2(_01740_),
    .A3(_01757_),
    .S1(net7964),
    .X(_07200_));
 sg13g2_inv_1 _20782_ (.Y(_07201_),
    .A(_07200_));
 sg13g2_mux4_1 _20783_ (.S0(net7970),
    .A0(net387),
    .A1(net404),
    .A2(_01741_),
    .A3(_01758_),
    .S1(net7960),
    .X(_07202_));
 sg13g2_or2_1 _20784_ (.X(_07203_),
    .B(_07202_),
    .A(_07200_));
 sg13g2_nor3_1 _20785_ (.A(_07154_),
    .B(_07188_),
    .C(_07203_),
    .Y(_07204_));
 sg13g2_nor2b_1 _20786_ (.A(net7615),
    .B_N(_07204_),
    .Y(_07205_));
 sg13g2_nor2_1 _20787_ (.A(net7387),
    .B(_07205_),
    .Y(_07206_));
 sg13g2_a221oi_1 _20788_ (.B2(_07153_),
    .C1(_07199_),
    .B1(_07206_),
    .A1(net7619),
    .Y(_07207_),
    .A2(_07184_));
 sg13g2_a21oi_1 _20789_ (.A1(net7412),
    .A2(_07121_),
    .Y(_07208_),
    .B1(_07207_));
 sg13g2_nor2_1 _20790_ (.A(net7613),
    .B(_07208_),
    .Y(_07209_));
 sg13g2_a21oi_1 _20791_ (.A1(_07171_),
    .A2(_07207_),
    .Y(_07210_),
    .B1(_07209_));
 sg13g2_nand2_1 _20792_ (.Y(_07211_),
    .A(net5950),
    .B(_07210_));
 sg13g2_o21ai_1 _20793_ (.B1(_07211_),
    .Y(_07212_),
    .A1(_08510_),
    .A2(net5950));
 sg13g2_nor2_1 _20794_ (.A(_01914_),
    .B(net5945),
    .Y(_07213_));
 sg13g2_inv_1 _20795_ (.Y(_07214_),
    .A(_07215_));
 sg13g2_o21ai_1 _20796_ (.B1(_07176_),
    .Y(_07215_),
    .A1(_07103_),
    .A2(_07133_));
 sg13g2_nand2_1 _20797_ (.Y(_07216_),
    .A(_07200_),
    .B(_07202_));
 sg13g2_nor2_1 _20798_ (.A(_07195_),
    .B(_07216_),
    .Y(_07217_));
 sg13g2_or2_1 _20799_ (.X(_07218_),
    .B(_07216_),
    .A(_07195_));
 sg13g2_nor2_1 _20800_ (.A(_07150_),
    .B(_07218_),
    .Y(_07219_));
 sg13g2_a21o_1 _20801_ (.A2(_07219_),
    .A1(net7305),
    .B1(_07215_),
    .X(_07220_));
 sg13g2_a221oi_1 _20802_ (.B2(net7620),
    .C1(_07153_),
    .B1(_07220_),
    .A1(net7303),
    .Y(_07221_),
    .A2(_07181_));
 sg13g2_a21oi_1 _20803_ (.A1(net5944),
    .A2(_07221_),
    .Y(_07222_),
    .B1(_07213_));
 sg13g2_a21oi_1 _20804_ (.A1(net7408),
    .A2(_07142_),
    .Y(_07223_),
    .B1(_07116_));
 sg13g2_nor2_1 _20805_ (.A(net7398),
    .B(_07223_),
    .Y(_07224_));
 sg13g2_nor2_1 _20806_ (.A(net7398),
    .B(net7618),
    .Y(_07225_));
 sg13g2_nand2_1 _20807_ (.Y(_07226_),
    .A(_07108_),
    .B(_07156_));
 sg13g2_and2_1 _20808_ (.A(_07168_),
    .B(_07204_),
    .X(_07227_));
 sg13g2_nor2_1 _20809_ (.A(_07226_),
    .B(_07227_),
    .Y(_07228_));
 sg13g2_nor2_1 _20810_ (.A(net7618),
    .B(_07195_),
    .Y(_07229_));
 sg13g2_nor3_1 _20811_ (.A(_07150_),
    .B(_07216_),
    .C(_07229_),
    .Y(_07230_));
 sg13g2_nor3_1 _20812_ (.A(_07181_),
    .B(_07228_),
    .C(_07230_),
    .Y(_07231_));
 sg13g2_a22oi_1 _20813_ (.Y(_07232_),
    .B1(_07231_),
    .B2(net7398),
    .A2(_07225_),
    .A1(net7390));
 sg13g2_nor2_1 _20814_ (.A(net7411),
    .B(_07232_),
    .Y(_07233_));
 sg13g2_nor2_1 _20815_ (.A(net7618),
    .B(_07172_),
    .Y(_07234_));
 sg13g2_nor4_1 _20816_ (.A(net5922),
    .B(_07224_),
    .C(_07233_),
    .D(_07234_),
    .Y(_07235_));
 sg13g2_a21o_1 _20817_ (.A2(net5922),
    .A1(net7673),
    .B1(_07235_),
    .X(_07236_));
 sg13g2_a21oi_1 _20818_ (.A1(_07148_),
    .A2(_07158_),
    .Y(_07237_),
    .B1(net7413));
 sg13g2_o21ai_1 _20819_ (.B1(net7621),
    .Y(_07238_),
    .A1(_07159_),
    .A2(_07237_));
 sg13g2_o21ai_1 _20820_ (.B1(_07103_),
    .Y(_07239_),
    .A1(_07148_),
    .A2(_07217_));
 sg13g2_o21ai_1 _20821_ (.B1(_07155_),
    .Y(_07240_),
    .A1(net7413),
    .A2(_07148_));
 sg13g2_a22oi_1 _20822_ (.Y(_07241_),
    .B1(_07240_),
    .B2(net7399),
    .A2(_07239_),
    .A1(net7395));
 sg13g2_nand2_1 _20823_ (.Y(_07242_),
    .A(net7388),
    .B(_07205_));
 sg13g2_nand3_1 _20824_ (.B(_07146_),
    .C(_07242_),
    .A(net7401),
    .Y(_07243_));
 sg13g2_nand3_1 _20825_ (.B(_07147_),
    .C(_07243_),
    .A(net7411),
    .Y(_07244_));
 sg13g2_nand3_1 _20826_ (.B(_07241_),
    .C(_07244_),
    .A(_07238_),
    .Y(_07245_));
 sg13g2_o21ai_1 _20827_ (.B1(_07245_),
    .Y(_07246_),
    .A1(net7621),
    .A2(_07172_));
 sg13g2_nand2_1 _20828_ (.Y(_07247_),
    .A(_01912_),
    .B(net5922));
 sg13g2_o21ai_1 _20829_ (.B1(_07247_),
    .Y(_07248_),
    .A1(net5922),
    .A2(_07246_));
 sg13g2_nor2_1 _20830_ (.A(_01911_),
    .B(net5945),
    .Y(_07249_));
 sg13g2_a22oi_1 _20831_ (.Y(_07250_),
    .B1(_07220_),
    .B2(net7617),
    .A2(net7301),
    .A1(net7303));
 sg13g2_a21oi_1 _20832_ (.A1(net5944),
    .A2(_07250_),
    .Y(_07251_),
    .B1(_07249_));
 sg13g2_nor2_1 _20833_ (.A(net7677),
    .B(net5945),
    .Y(_07252_));
 sg13g2_mux2_1 _20834_ (.A0(net391),
    .A1(_01780_),
    .S(net7951),
    .X(_07253_));
 sg13g2_nor2b_1 _20835_ (.A(net7964),
    .B_N(net409),
    .Y(_07254_));
 sg13g2_a21oi_1 _20836_ (.A1(net7964),
    .A2(_01763_),
    .Y(_07255_),
    .B1(_07254_));
 sg13g2_nand2_1 _20837_ (.Y(_07256_),
    .A(net7970),
    .B(_07253_));
 sg13g2_o21ai_1 _20838_ (.B1(_07256_),
    .Y(_07257_),
    .A1(net7970),
    .A2(_07255_));
 sg13g2_o21ai_1 _20839_ (.B1(_07202_),
    .Y(_07258_),
    .A1(_07201_),
    .A2(_07257_));
 sg13g2_nand2_1 _20840_ (.Y(_07259_),
    .A(net7304),
    .B(net7388));
 sg13g2_a21oi_1 _20841_ (.A1(_07149_),
    .A2(_07258_),
    .Y(_07260_),
    .B1(_07259_));
 sg13g2_a21oi_1 _20842_ (.A1(_07215_),
    .A2(_07257_),
    .Y(_07261_),
    .B1(_07260_));
 sg13g2_a21oi_1 _20843_ (.A1(net5945),
    .A2(_07261_),
    .Y(_07262_),
    .B1(_07252_));
 sg13g2_nor2_1 _20844_ (.A(net7678),
    .B(net5942),
    .Y(_07263_));
 sg13g2_mux2_1 _20845_ (.A0(net390),
    .A1(_01779_),
    .S(net7955),
    .X(_07264_));
 sg13g2_nor2b_1 _20846_ (.A(net7965),
    .B_N(net408),
    .Y(_07265_));
 sg13g2_a21oi_1 _20847_ (.A1(net7965),
    .A2(_01762_),
    .Y(_07266_),
    .B1(_07265_));
 sg13g2_nand2_1 _20848_ (.Y(_07267_),
    .A(net7967),
    .B(_07264_));
 sg13g2_o21ai_1 _20849_ (.B1(_07267_),
    .Y(_07268_),
    .A1(net7967),
    .A2(_07266_));
 sg13g2_a21oi_1 _20850_ (.A1(_07143_),
    .A2(_07202_),
    .Y(_07269_),
    .B1(net7439));
 sg13g2_nor2_1 _20851_ (.A(_07194_),
    .B(_07269_),
    .Y(_07270_));
 sg13g2_o21ai_1 _20852_ (.B1(_07203_),
    .Y(_07271_),
    .A1(_07218_),
    .A2(_07268_));
 sg13g2_o21ai_1 _20853_ (.B1(_07169_),
    .Y(_07272_),
    .A1(_07270_),
    .A2(_07271_));
 sg13g2_o21ai_1 _20854_ (.B1(_07272_),
    .Y(_07273_),
    .A1(net7405),
    .A2(net7615));
 sg13g2_o21ai_1 _20855_ (.B1(net7390),
    .Y(_07274_),
    .A1(net7407),
    .A2(net7403));
 sg13g2_a221oi_1 _20856_ (.B2(net7386),
    .C1(net7302),
    .B1(_07274_),
    .A1(net7390),
    .Y(_07275_),
    .A2(_07273_));
 sg13g2_a21oi_1 _20857_ (.A1(_07215_),
    .A2(_07268_),
    .Y(_07276_),
    .B1(_07275_));
 sg13g2_a21oi_1 _20858_ (.A1(net5942),
    .A2(_07276_),
    .Y(_07277_),
    .B1(_07263_));
 sg13g2_nor2_1 _20859_ (.A(_01908_),
    .B(net5945),
    .Y(_07278_));
 sg13g2_nand2_1 _20860_ (.Y(_07279_),
    .A(_07139_),
    .B(_07147_));
 sg13g2_o21ai_1 _20861_ (.B1(net7305),
    .Y(_07280_),
    .A1(_07180_),
    .A2(net7050));
 sg13g2_o21ai_1 _20862_ (.B1(_07280_),
    .Y(_07281_),
    .A1(_07243_),
    .A2(_07279_));
 sg13g2_a21oi_1 _20863_ (.A1(net7619),
    .A2(_07220_),
    .Y(_07282_),
    .B1(_07281_));
 sg13g2_a21oi_1 _20864_ (.A1(net5945),
    .A2(_07282_),
    .Y(_07283_),
    .B1(_07278_));
 sg13g2_nor2_1 _20865_ (.A(net7680),
    .B(net5943),
    .Y(_07284_));
 sg13g2_and2_1 _20866_ (.A(net7390),
    .B(_07184_),
    .X(_07285_));
 sg13g2_nor2b_1 _20867_ (.A(net7948),
    .B_N(net389),
    .Y(_07286_));
 sg13g2_a21oi_1 _20868_ (.A1(net7948),
    .A2(_01778_),
    .Y(_07287_),
    .B1(_07286_));
 sg13g2_mux2_1 _20869_ (.A0(net406),
    .A1(_01760_),
    .S(net7958),
    .X(_07288_));
 sg13g2_nand2_1 _20870_ (.Y(_07289_),
    .A(_15152_),
    .B(_07288_));
 sg13g2_o21ai_1 _20871_ (.B1(_07289_),
    .Y(_07290_),
    .A1(_15152_),
    .A2(_07287_));
 sg13g2_nand2_1 _20872_ (.Y(_07291_),
    .A(_07149_),
    .B(_07202_));
 sg13g2_nor2_1 _20873_ (.A(_07201_),
    .B(_07290_),
    .Y(_07292_));
 sg13g2_nor2_1 _20874_ (.A(_07291_),
    .B(_07292_),
    .Y(_07293_));
 sg13g2_o21ai_1 _20875_ (.B1(net7388),
    .Y(_07294_),
    .A1(_07274_),
    .A2(_07293_));
 sg13g2_nand2_1 _20876_ (.Y(_07295_),
    .A(net7301),
    .B(_07200_));
 sg13g2_a21oi_1 _20877_ (.A1(_07294_),
    .A2(_07295_),
    .Y(_07296_),
    .B1(net7302));
 sg13g2_a221oi_1 _20878_ (.B2(_07215_),
    .C1(_07296_),
    .B1(_07290_),
    .A1(_07200_),
    .Y(_07297_),
    .A2(_07285_));
 sg13g2_a21oi_1 _20879_ (.A1(net5945),
    .A2(_07297_),
    .Y(_07298_),
    .B1(_07284_));
 sg13g2_nor2_1 _20880_ (.A(net7681),
    .B(net5943),
    .Y(_07299_));
 sg13g2_nor2b_1 _20881_ (.A(net7950),
    .B_N(net388),
    .Y(_07300_));
 sg13g2_a21oi_1 _20882_ (.A1(net7950),
    .A2(_01777_),
    .Y(_07301_),
    .B1(_07300_));
 sg13g2_nand2_1 _20883_ (.Y(_07302_),
    .A(net7969),
    .B(_07301_));
 sg13g2_mux2_1 _20884_ (.A0(net405),
    .A1(_01759_),
    .S(net7960),
    .X(_07303_));
 sg13g2_o21ai_1 _20885_ (.B1(_07302_),
    .Y(_07304_),
    .A1(net7969),
    .A2(_07303_));
 sg13g2_nor2_1 _20886_ (.A(_07214_),
    .B(_07304_),
    .Y(_07305_));
 sg13g2_a22oi_1 _20887_ (.Y(_07306_),
    .B1(net7388),
    .B2(_07130_),
    .A2(net7301),
    .A1(net7616));
 sg13g2_o21ai_1 _20888_ (.B1(net7388),
    .Y(_07307_),
    .A1(_07116_),
    .A2(_07228_));
 sg13g2_nor2b_1 _20889_ (.A(_07226_),
    .B_N(_07227_),
    .Y(_07308_));
 sg13g2_nor2_1 _20890_ (.A(net7386),
    .B(_07291_),
    .Y(_07309_));
 sg13g2_nand2_1 _20891_ (.Y(_07310_),
    .A(_07200_),
    .B(_07304_));
 sg13g2_a22oi_1 _20892_ (.Y(_07311_),
    .B1(_07309_),
    .B2(_07310_),
    .A2(_07308_),
    .A1(_07123_));
 sg13g2_nand3_1 _20893_ (.B(_07307_),
    .C(_07311_),
    .A(_07306_),
    .Y(_07312_));
 sg13g2_a221oi_1 _20894_ (.B2(net7304),
    .C1(_07305_),
    .B1(_07312_),
    .A1(net7616),
    .Y(_07313_),
    .A2(_07285_));
 sg13g2_a21oi_1 _20895_ (.A1(net5943),
    .A2(_07313_),
    .Y(_07314_),
    .B1(_07299_));
 sg13g2_nor2_1 _20896_ (.A(_01905_),
    .B(net5943),
    .Y(_07315_));
 sg13g2_a22oi_1 _20897_ (.Y(_07316_),
    .B1(net7388),
    .B2(_07116_),
    .A2(_07181_),
    .A1(_07132_));
 sg13g2_mux2_1 _20898_ (.A0(net387),
    .A1(_01776_),
    .S(net7955),
    .X(_07317_));
 sg13g2_nor2b_1 _20899_ (.A(net7964),
    .B_N(net404),
    .Y(_07318_));
 sg13g2_a21oi_1 _20900_ (.A1(net7960),
    .A2(_01758_),
    .Y(_07319_),
    .B1(_07318_));
 sg13g2_nand2_1 _20901_ (.Y(_07320_),
    .A(net7970),
    .B(_07317_));
 sg13g2_o21ai_1 _20902_ (.B1(_07320_),
    .Y(_07321_),
    .A1(net7970),
    .A2(_07319_));
 sg13g2_o21ai_1 _20903_ (.B1(_07309_),
    .Y(_07322_),
    .A1(_07201_),
    .A2(_07321_));
 sg13g2_nand2_1 _20904_ (.Y(_07323_),
    .A(net7389),
    .B(net7050));
 sg13g2_nand2_1 _20905_ (.Y(_07324_),
    .A(net7617),
    .B(_07308_));
 sg13g2_nand4_1 _20906_ (.B(_07322_),
    .C(_07323_),
    .A(_07316_),
    .Y(_07325_),
    .D(_07324_));
 sg13g2_nand2_1 _20907_ (.Y(_07326_),
    .A(net7403),
    .B(net7615));
 sg13g2_nand2_1 _20908_ (.Y(_07327_),
    .A(net7400),
    .B(net7617));
 sg13g2_o21ai_1 _20909_ (.B1(_07326_),
    .Y(_07328_),
    .A1(net7406),
    .A2(_07327_));
 sg13g2_nand3_1 _20910_ (.B(net7392),
    .C(_07328_),
    .A(_07102_),
    .Y(_07329_));
 sg13g2_nor2_1 _20911_ (.A(net7411),
    .B(net7401),
    .Y(_07330_));
 sg13g2_nand3_1 _20912_ (.B(net7615),
    .C(_07330_),
    .A(net7390),
    .Y(_07331_));
 sg13g2_a21oi_1 _20913_ (.A1(_07329_),
    .A2(_07331_),
    .Y(_07332_),
    .B1(net7306));
 sg13g2_a221oi_1 _20914_ (.B2(net7304),
    .C1(_07332_),
    .B1(_07325_),
    .A1(_07215_),
    .Y(_07333_),
    .A2(_07321_));
 sg13g2_a21oi_1 _20915_ (.A1(net5943),
    .A2(_07333_),
    .Y(_07334_),
    .B1(_07315_));
 sg13g2_nor2_1 _20916_ (.A(net7683),
    .B(net5953),
    .Y(_07335_));
 sg13g2_nor2b_1 _20917_ (.A(net7954),
    .B_N(net386),
    .Y(_07336_));
 sg13g2_a21oi_1 _20918_ (.A1(net7954),
    .A2(_01775_),
    .Y(_07337_),
    .B1(_07336_));
 sg13g2_nand2_1 _20919_ (.Y(_07338_),
    .A(net7974),
    .B(_07337_));
 sg13g2_mux2_1 _20920_ (.A0(net403),
    .A1(_01757_),
    .S(net7961),
    .X(_07339_));
 sg13g2_o21ai_1 _20921_ (.B1(_07338_),
    .Y(_07340_),
    .A1(net7974),
    .A2(_07339_));
 sg13g2_mux2_1 _20922_ (.A0(net7619),
    .A1(net7613),
    .S(net7403),
    .X(_07341_));
 sg13g2_nand3_1 _20923_ (.B(net7307),
    .C(_07341_),
    .A(net7393),
    .Y(_07342_));
 sg13g2_o21ai_1 _20924_ (.B1(_07342_),
    .Y(_07343_),
    .A1(net7307),
    .A2(_07340_));
 sg13g2_nor2_1 _20925_ (.A(net7407),
    .B(net7391),
    .Y(_07344_));
 sg13g2_nor2_1 _20926_ (.A(net7403),
    .B(net7392),
    .Y(_07345_));
 sg13g2_nand2b_1 _20927_ (.Y(_07346_),
    .B(_07345_),
    .A_N(net7613));
 sg13g2_o21ai_1 _20928_ (.B1(_07346_),
    .Y(_07347_),
    .A1(net7390),
    .A2(_07141_));
 sg13g2_a22oi_1 _20929_ (.Y(_07348_),
    .B1(_07347_),
    .B2(_07109_),
    .A2(_07340_),
    .A1(_07174_));
 sg13g2_nand2_1 _20930_ (.Y(_07349_),
    .A(_07200_),
    .B(_07340_));
 sg13g2_a22oi_1 _20931_ (.Y(_07350_),
    .B1(_07309_),
    .B2(_07349_),
    .A2(net7613),
    .A1(net7301));
 sg13g2_o21ai_1 _20932_ (.B1(net7618),
    .Y(_07351_),
    .A1(_07130_),
    .A2(_07308_));
 sg13g2_nand4_1 _20933_ (.B(_07307_),
    .C(_07350_),
    .A(net7398),
    .Y(_07352_),
    .D(_07351_));
 sg13g2_o21ai_1 _20934_ (.B1(_07352_),
    .Y(_07353_),
    .A1(net7398),
    .A2(_07348_));
 sg13g2_nor2_1 _20935_ (.A(net7411),
    .B(_07353_),
    .Y(_07354_));
 sg13g2_a21oi_1 _20936_ (.A1(net7411),
    .A2(_07343_),
    .Y(_07355_),
    .B1(_07354_));
 sg13g2_a21oi_1 _20937_ (.A1(net5952),
    .A2(_07355_),
    .Y(_07356_),
    .B1(_07335_));
 sg13g2_nor2_1 _20938_ (.A(net7684),
    .B(net5942),
    .Y(_07357_));
 sg13g2_nor2b_1 _20939_ (.A(net7948),
    .B_N(net416),
    .Y(_07358_));
 sg13g2_a21oi_1 _20940_ (.A1(net7948),
    .A2(_01774_),
    .Y(_07359_),
    .B1(_07358_));
 sg13g2_mux2_1 _20941_ (.A0(net402),
    .A1(_01756_),
    .S(net7958),
    .X(_07360_));
 sg13g2_nand2_1 _20942_ (.Y(_07361_),
    .A(_15152_),
    .B(_07360_));
 sg13g2_o21ai_1 _20943_ (.B1(_07361_),
    .Y(_07362_),
    .A1(_15152_),
    .A2(_07359_));
 sg13g2_nor2_1 _20944_ (.A(net7393),
    .B(_07330_),
    .Y(_07363_));
 sg13g2_nor3_1 _20945_ (.A(net7306),
    .B(net7386),
    .C(_07363_),
    .Y(_07364_));
 sg13g2_o21ai_1 _20946_ (.B1(_07309_),
    .Y(_07365_),
    .A1(_07201_),
    .A2(_07362_));
 sg13g2_o21ai_1 _20947_ (.B1(net7619),
    .Y(_07366_),
    .A1(_07181_),
    .A2(_07308_));
 sg13g2_nand3_1 _20948_ (.B(_07365_),
    .C(_07366_),
    .A(_07307_),
    .Y(_07367_));
 sg13g2_a221oi_1 _20949_ (.B2(net7304),
    .C1(_07364_),
    .B1(_07367_),
    .A1(_07215_),
    .Y(_07368_),
    .A2(_07362_));
 sg13g2_a21oi_1 _20950_ (.A1(net5942),
    .A2(_07368_),
    .Y(_07369_),
    .B1(_07357_));
 sg13g2_mux2_1 _20951_ (.A0(net415),
    .A1(_01773_),
    .S(net7952),
    .X(_07370_));
 sg13g2_nor2b_1 _20952_ (.A(net7962),
    .B_N(net401),
    .Y(_07371_));
 sg13g2_a21oi_1 _20953_ (.A1(net7962),
    .A2(_01755_),
    .Y(_07372_),
    .B1(_07371_));
 sg13g2_nand2_1 _20954_ (.Y(_07373_),
    .A(net7971),
    .B(_07370_));
 sg13g2_o21ai_1 _20955_ (.B1(_07373_),
    .Y(_07374_),
    .A1(net7971),
    .A2(_07372_));
 sg13g2_and2_1 _20956_ (.A(net7405),
    .B(net7620),
    .X(_07375_));
 sg13g2_a22oi_1 _20957_ (.Y(_07376_),
    .B1(_07216_),
    .B2(_07375_),
    .A2(net7611),
    .A1(net7406));
 sg13g2_o21ai_1 _20958_ (.B1(_07323_),
    .Y(_07377_),
    .A1(net7392),
    .A2(_07376_));
 sg13g2_or2_1 _20959_ (.X(_07378_),
    .B(_07308_),
    .A(_07116_));
 sg13g2_a221oi_1 _20960_ (.B2(net7620),
    .C1(_07377_),
    .B1(_07378_),
    .A1(_07219_),
    .Y(_07379_),
    .A2(_07374_));
 sg13g2_and3_1 _20961_ (.X(_07380_),
    .A(net7410),
    .B(net7620),
    .C(net7307));
 sg13g2_a221oi_1 _20962_ (.B2(_07374_),
    .C1(_07380_),
    .B1(net7051),
    .A1(_07184_),
    .Y(_07381_),
    .A2(net7611));
 sg13g2_o21ai_1 _20963_ (.B1(_07381_),
    .Y(_07382_),
    .A1(_07179_),
    .A2(_07379_));
 sg13g2_mux2_1 _20964_ (.A0(_01902_),
    .A1(_07382_),
    .S(net5948),
    .X(_07383_));
 sg13g2_nor2_1 _20965_ (.A(net7693),
    .B(net5947),
    .Y(_07384_));
 sg13g2_nand2_1 _20966_ (.Y(_07385_),
    .A(net7412),
    .B(net7307));
 sg13g2_o21ai_1 _20967_ (.B1(net7397),
    .Y(_07386_),
    .A1(_07116_),
    .A2(_07180_));
 sg13g2_o21ai_1 _20968_ (.B1(_07385_),
    .Y(_07387_),
    .A1(net7412),
    .A2(_07386_));
 sg13g2_mux2_1 _20969_ (.A0(net414),
    .A1(_01771_),
    .S(net7952),
    .X(_07388_));
 sg13g2_nor2b_1 _20970_ (.A(net7962),
    .B_N(net400),
    .Y(_07389_));
 sg13g2_a21oi_1 _20971_ (.A1(net7962),
    .A2(_01754_),
    .Y(_07390_),
    .B1(_07389_));
 sg13g2_nand2_1 _20972_ (.Y(_07391_),
    .A(net7971),
    .B(_07388_));
 sg13g2_o21ai_1 _20973_ (.B1(_07391_),
    .Y(_07392_),
    .A1(net7971),
    .A2(_07390_));
 sg13g2_nand2_1 _20974_ (.Y(_07393_),
    .A(net7400),
    .B(net7439));
 sg13g2_a22oi_1 _20975_ (.Y(_07394_),
    .B1(_07393_),
    .B2(net7392),
    .A2(_07345_),
    .A1(_07141_));
 sg13g2_nor3_1 _20976_ (.A(_07102_),
    .B(net7306),
    .C(_07394_),
    .Y(_07395_));
 sg13g2_a21o_1 _20977_ (.A2(_07392_),
    .A1(net7051),
    .B1(_07395_),
    .X(_07396_));
 sg13g2_nor3_1 _20978_ (.A(_07195_),
    .B(_07216_),
    .C(_07392_),
    .Y(_07397_));
 sg13g2_a21o_1 _20979_ (.A2(_07216_),
    .A1(_07142_),
    .B1(_07397_),
    .X(_07398_));
 sg13g2_o21ai_1 _20980_ (.B1(_07323_),
    .Y(_07399_),
    .A1(_07150_),
    .A2(_07398_));
 sg13g2_a221oi_1 _20981_ (.B2(net7304),
    .C1(_07396_),
    .B1(_07399_),
    .A1(net7618),
    .Y(_07400_),
    .A2(_07387_));
 sg13g2_a21oi_1 _20982_ (.A1(net5949),
    .A2(_07400_),
    .Y(_07401_),
    .B1(_07384_));
 sg13g2_nor2_1 _20983_ (.A(net7702),
    .B(net5948),
    .Y(_07402_));
 sg13g2_mux2_1 _20984_ (.A0(net413),
    .A1(_01770_),
    .S(net7953),
    .X(_07403_));
 sg13g2_nor2b_1 _20985_ (.A(net7962),
    .B_N(net399),
    .Y(_07404_));
 sg13g2_a21oi_1 _20986_ (.A1(net7962),
    .A2(_01753_),
    .Y(_07405_),
    .B1(_07404_));
 sg13g2_nand2_1 _20987_ (.Y(_07406_),
    .A(net7971),
    .B(_07403_));
 sg13g2_o21ai_1 _20988_ (.B1(_07406_),
    .Y(_07407_),
    .A1(net7971),
    .A2(_07405_));
 sg13g2_and2_1 _20989_ (.A(net7402),
    .B(_07123_),
    .X(_07408_));
 sg13g2_a22oi_1 _20990_ (.Y(_07409_),
    .B1(_07408_),
    .B2(net7392),
    .A2(net7620),
    .A1(net7400));
 sg13g2_nor3_1 _20991_ (.A(net7410),
    .B(_07134_),
    .C(_07409_),
    .Y(_07410_));
 sg13g2_a22oi_1 _20992_ (.Y(_07411_),
    .B1(_07159_),
    .B2(_07407_),
    .A2(net7621),
    .A1(net7404));
 sg13g2_nor2_1 _20993_ (.A(_07103_),
    .B(_07411_),
    .Y(_07412_));
 sg13g2_a21oi_1 _20994_ (.A1(net7404),
    .A2(_07217_),
    .Y(_07413_),
    .B1(net7392));
 sg13g2_nand3_1 _20995_ (.B(_07217_),
    .C(_07407_),
    .A(_07160_),
    .Y(_07414_));
 sg13g2_a21oi_1 _20996_ (.A1(_07135_),
    .A2(_07414_),
    .Y(_07415_),
    .B1(net7406));
 sg13g2_a21oi_1 _20997_ (.A1(net7621),
    .A2(_07413_),
    .Y(_07416_),
    .B1(_07415_));
 sg13g2_a21oi_1 _20998_ (.A1(_07323_),
    .A2(_07416_),
    .Y(_07417_),
    .B1(_07122_));
 sg13g2_nor3_1 _20999_ (.A(_07410_),
    .B(_07412_),
    .C(_07417_),
    .Y(_07418_));
 sg13g2_inv_1 _21000_ (.Y(_07419_),
    .A(_07418_));
 sg13g2_a22oi_1 _21001_ (.Y(_07420_),
    .B1(_07419_),
    .B2(_07172_),
    .A2(_07407_),
    .A1(_07177_));
 sg13g2_a21oi_1 _21002_ (.A1(net5948),
    .A2(_07420_),
    .Y(_07421_),
    .B1(_07402_));
 sg13g2_mux2_1 _21003_ (.A0(net412),
    .A1(_01769_),
    .S(net7953),
    .X(_07422_));
 sg13g2_nor2b_1 _21004_ (.A(net7963),
    .B_N(net398),
    .Y(_07423_));
 sg13g2_a21oi_1 _21005_ (.A1(net7963),
    .A2(_01752_),
    .Y(_07424_),
    .B1(_07423_));
 sg13g2_nand2_1 _21006_ (.Y(_07425_),
    .A(net7973),
    .B(_07422_));
 sg13g2_o21ai_1 _21007_ (.B1(_07425_),
    .Y(_07426_),
    .A1(net7972),
    .A2(_07424_));
 sg13g2_nand2_1 _21008_ (.Y(_07427_),
    .A(net7410),
    .B(net7390));
 sg13g2_nand2_1 _21009_ (.Y(_07428_),
    .A(net7307),
    .B(net7617));
 sg13g2_a21oi_1 _21010_ (.A1(_07131_),
    .A2(_07427_),
    .Y(_07429_),
    .B1(_07428_));
 sg13g2_a21oi_1 _21011_ (.A1(net7051),
    .A2(_07426_),
    .Y(_07430_),
    .B1(_07429_));
 sg13g2_nor2_1 _21012_ (.A(net7392),
    .B(_07218_),
    .Y(_07431_));
 sg13g2_nand3_1 _21013_ (.B(_07426_),
    .C(_07431_),
    .A(net7403),
    .Y(_07432_));
 sg13g2_a21oi_1 _21014_ (.A1(_07327_),
    .A2(_07432_),
    .Y(_07433_),
    .B1(net7406));
 sg13g2_a221oi_1 _21015_ (.B2(net7617),
    .C1(_07433_),
    .B1(_07413_),
    .A1(_07194_),
    .Y(_07434_),
    .A2(net7050));
 sg13g2_o21ai_1 _21016_ (.B1(_07430_),
    .Y(_07435_),
    .A1(_07179_),
    .A2(_07434_));
 sg13g2_nand2_1 _21017_ (.Y(_07436_),
    .A(net5949),
    .B(_07435_));
 sg13g2_o21ai_1 _21018_ (.B1(_07436_),
    .Y(_07437_),
    .A1(net7519),
    .A2(net5947));
 sg13g2_nor2_1 _21019_ (.A(net7403),
    .B(_07140_),
    .Y(_07438_));
 sg13g2_nand2_1 _21020_ (.Y(_07439_),
    .A(_07130_),
    .B(_07140_));
 sg13g2_o21ai_1 _21021_ (.B1(_07439_),
    .Y(_07440_),
    .A1(_07427_),
    .A2(_07438_));
 sg13g2_nand2_1 _21022_ (.Y(_07441_),
    .A(_07122_),
    .B(_07440_));
 sg13g2_nand3_1 _21023_ (.B(_07178_),
    .C(_07345_),
    .A(net7619),
    .Y(_07442_));
 sg13g2_a21oi_1 _21024_ (.A1(_07441_),
    .A2(_07442_),
    .Y(_07443_),
    .B1(net7407));
 sg13g2_nand3_1 _21025_ (.B(_07205_),
    .C(_07443_),
    .A(_07145_),
    .Y(_07444_));
 sg13g2_a21oi_1 _21026_ (.A1(_07280_),
    .A2(_07444_),
    .Y(_07445_),
    .B1(net7387));
 sg13g2_nand2_1 _21027_ (.Y(_07446_),
    .A(net7405),
    .B(_07140_));
 sg13g2_a21oi_1 _21028_ (.A1(_07160_),
    .A2(_07218_),
    .Y(_07447_),
    .B1(_07156_));
 sg13g2_nor2_1 _21029_ (.A(_07446_),
    .B(_07447_),
    .Y(_07448_));
 sg13g2_mux2_1 _21030_ (.A0(net411),
    .A1(_01768_),
    .S(net7954),
    .X(_07449_));
 sg13g2_inv_1 _21031_ (.Y(_07450_),
    .A(_01946_));
 sg13g2_nor2b_1 _21032_ (.A(net7961),
    .B_N(net397),
    .Y(_07451_));
 sg13g2_a21oi_1 _21033_ (.A1(net7961),
    .A2(_01751_),
    .Y(_07452_),
    .B1(_07451_));
 sg13g2_nand2_1 _21034_ (.Y(_07453_),
    .A(net7974),
    .B(_07449_));
 sg13g2_o21ai_1 _21035_ (.B1(_07453_),
    .Y(_07454_),
    .A1(net7974),
    .A2(_07452_));
 sg13g2_a21oi_1 _21036_ (.A1(_07219_),
    .A2(_07454_),
    .Y(_07455_),
    .B1(_07448_));
 sg13g2_a22oi_1 _21037_ (.Y(_07456_),
    .B1(_07454_),
    .B2(net7051),
    .A2(_07443_),
    .A1(_07140_));
 sg13g2_o21ai_1 _21038_ (.B1(_07456_),
    .Y(_07457_),
    .A1(_07179_),
    .A2(_07455_));
 sg13g2_o21ai_1 _21039_ (.B1(net5949),
    .Y(_07458_),
    .A1(_07445_),
    .A2(_07457_));
 sg13g2_o21ai_1 _21040_ (.B1(_07458_),
    .Y(_07459_),
    .A1(_09041_),
    .A2(net5950));
 sg13g2_a21oi_1 _21041_ (.A1(net7303),
    .A2(_07219_),
    .Y(_07460_),
    .B1(_07175_));
 sg13g2_mux2_1 _21042_ (.A0(_01897_),
    .A1(_07460_),
    .S(net5943),
    .X(_07461_));
 sg13g2_nand2b_1 _21043_ (.Y(_07462_),
    .B(net7402),
    .A_N(_07146_));
 sg13g2_a22oi_1 _21044_ (.Y(_07463_),
    .B1(_07462_),
    .B2(_07139_),
    .A2(_07157_),
    .A1(net7409));
 sg13g2_nand2_1 _21045_ (.Y(_07464_),
    .A(_07147_),
    .B(net7611));
 sg13g2_mux2_1 _21046_ (.A0(net410),
    .A1(_01767_),
    .S(net7951),
    .X(_07465_));
 sg13g2_nor2b_1 _21047_ (.A(net7960),
    .B_N(net395),
    .Y(_07466_));
 sg13g2_a21oi_1 _21048_ (.A1(net7960),
    .A2(_01749_),
    .Y(_07467_),
    .B1(_07466_));
 sg13g2_nand2_1 _21049_ (.Y(_07468_),
    .A(net7969),
    .B(_07465_));
 sg13g2_o21ai_1 _21050_ (.B1(_07468_),
    .Y(_07469_),
    .A1(net7969),
    .A2(_07467_));
 sg13g2_nand3_1 _21051_ (.B(_07149_),
    .C(net7611),
    .A(_07139_),
    .Y(_07470_));
 sg13g2_nand2_1 _21052_ (.Y(_07471_),
    .A(_07280_),
    .B(_07470_));
 sg13g2_a22oi_1 _21053_ (.Y(_07472_),
    .B1(_07471_),
    .B2(net7389),
    .A2(_07469_),
    .A1(_07220_));
 sg13g2_o21ai_1 _21054_ (.B1(_07472_),
    .Y(_07473_),
    .A1(_07463_),
    .A2(_07464_));
 sg13g2_mux2_1 _21055_ (.A0(_01896_),
    .A1(_07473_),
    .S(net5947),
    .X(_07474_));
 sg13g2_nor2_1 _21056_ (.A(_01895_),
    .B(net5947),
    .Y(_07475_));
 sg13g2_mux2_1 _21057_ (.A0(net407),
    .A1(_01766_),
    .S(net7953),
    .X(_07476_));
 sg13g2_nor2b_1 _21058_ (.A(net7961),
    .B_N(net394),
    .Y(_07477_));
 sg13g2_a21oi_1 _21059_ (.A1(net7961),
    .A2(_01748_),
    .Y(_07478_),
    .B1(_07477_));
 sg13g2_nand2_1 _21060_ (.Y(_07479_),
    .A(net7972),
    .B(_07476_));
 sg13g2_o21ai_1 _21061_ (.B1(_07479_),
    .Y(_07480_),
    .A1(net7972),
    .A2(_07478_));
 sg13g2_o21ai_1 _21062_ (.B1(net7404),
    .Y(_07481_),
    .A1(_07218_),
    .A2(_07480_));
 sg13g2_a21o_1 _21063_ (.A2(_07481_),
    .A1(net7391),
    .B1(net7400),
    .X(_07482_));
 sg13g2_nand2_1 _21064_ (.Y(_07483_),
    .A(net7407),
    .B(_07194_));
 sg13g2_nor2_1 _21065_ (.A(net7393),
    .B(net7386),
    .Y(_07484_));
 sg13g2_nand2_1 _21066_ (.Y(_07485_),
    .A(_07180_),
    .B(net7389));
 sg13g2_nand2_1 _21067_ (.Y(_07486_),
    .A(_07323_),
    .B(_07485_));
 sg13g2_nand3_1 _21068_ (.B(net7391),
    .C(net7612),
    .A(_07116_),
    .Y(_07487_));
 sg13g2_nand4_1 _21069_ (.B(_07482_),
    .C(_07485_),
    .A(_07323_),
    .Y(_07488_),
    .D(_07487_));
 sg13g2_a21o_1 _21070_ (.A2(_07480_),
    .A1(net7402),
    .B1(_07344_),
    .X(_07489_));
 sg13g2_a22oi_1 _21071_ (.Y(_07490_),
    .B1(_07489_),
    .B2(_07103_),
    .A2(_07480_),
    .A1(net7406));
 sg13g2_nand3_1 _21072_ (.B(net7396),
    .C(_07480_),
    .A(net7410),
    .Y(_07491_));
 sg13g2_o21ai_1 _21073_ (.B1(_07491_),
    .Y(_07492_),
    .A1(net7396),
    .A2(_07490_));
 sg13g2_nand2b_1 _21074_ (.Y(_07493_),
    .B(net7387),
    .A_N(_07462_));
 sg13g2_nor4_1 _21075_ (.A(_07103_),
    .B(net7306),
    .C(_07148_),
    .D(net7439),
    .Y(_07494_));
 sg13g2_a221oi_1 _21076_ (.B2(_07494_),
    .C1(_07492_),
    .B1(_07493_),
    .A1(net7304),
    .Y(_07495_),
    .A2(_07488_));
 sg13g2_a21oi_1 _21077_ (.A1(net5947),
    .A2(_07495_),
    .Y(_07496_),
    .B1(_07475_));
 sg13g2_nand3_1 _21078_ (.B(net7391),
    .C(_07493_),
    .A(_07102_),
    .Y(_07497_));
 sg13g2_o21ai_1 _21079_ (.B1(_07497_),
    .Y(_07498_),
    .A1(net7410),
    .A2(net7390));
 sg13g2_and2_1 _21080_ (.A(net7307),
    .B(net7616),
    .X(_07499_));
 sg13g2_mux2_1 _21081_ (.A0(net396),
    .A1(_01765_),
    .S(net7948),
    .X(_07500_));
 sg13g2_nor2b_1 _21082_ (.A(net7957),
    .B_N(net393),
    .Y(_07501_));
 sg13g2_a21oi_1 _21083_ (.A1(net7957),
    .A2(_01747_),
    .Y(_07502_),
    .B1(_07501_));
 sg13g2_nand2_1 _21084_ (.Y(_07503_),
    .A(net7968),
    .B(_07500_));
 sg13g2_o21ai_1 _21085_ (.B1(_07503_),
    .Y(_07504_),
    .A1(net7967),
    .A2(_07502_));
 sg13g2_a22oi_1 _21086_ (.Y(_07505_),
    .B1(_07504_),
    .B2(net7051),
    .A2(_07499_),
    .A1(_07498_));
 sg13g2_a22oi_1 _21087_ (.Y(_07506_),
    .B1(_07431_),
    .B2(_07504_),
    .A2(_07218_),
    .A1(net7616));
 sg13g2_nand2_1 _21088_ (.Y(_07507_),
    .A(net7616),
    .B(_07345_));
 sg13g2_o21ai_1 _21089_ (.B1(_07507_),
    .Y(_07508_),
    .A1(net7400),
    .A2(_07506_));
 sg13g2_a221oi_1 _21090_ (.B2(_07109_),
    .C1(_07486_),
    .B1(_07508_),
    .A1(net7308),
    .Y(_07509_),
    .A2(net7616));
 sg13g2_o21ai_1 _21091_ (.B1(_07505_),
    .Y(_07510_),
    .A1(_07179_),
    .A2(_07509_));
 sg13g2_mux2_1 _21092_ (.A0(net7809),
    .A1(_07510_),
    .S(net5948),
    .X(_07511_));
 sg13g2_nor2_1 _21093_ (.A(net7819),
    .B(net5948),
    .Y(_07512_));
 sg13g2_nor2b_1 _21094_ (.A(net7949),
    .B_N(net385),
    .Y(_07513_));
 sg13g2_a21oi_1 _21095_ (.A1(net7949),
    .A2(_01764_),
    .Y(_07514_),
    .B1(_07513_));
 sg13g2_mux2_1 _21096_ (.A0(net392),
    .A1(_01746_),
    .S(net7957),
    .X(_07515_));
 sg13g2_nand2_1 _21097_ (.Y(_07516_),
    .A(_15152_),
    .B(_07515_));
 sg13g2_o21ai_1 _21098_ (.B1(_07516_),
    .Y(_07517_),
    .A1(_15152_),
    .A2(_07514_));
 sg13g2_a21oi_1 _21099_ (.A1(net7614),
    .A2(_07493_),
    .Y(_07518_),
    .B1(_07128_));
 sg13g2_nor2_1 _21100_ (.A(net7306),
    .B(_07518_),
    .Y(_07519_));
 sg13g2_a21oi_1 _21101_ (.A1(net7306),
    .A2(_07517_),
    .Y(_07520_),
    .B1(_07519_));
 sg13g2_nor2_1 _21102_ (.A(net7409),
    .B(_07520_),
    .Y(_07521_));
 sg13g2_nand2b_1 _21103_ (.Y(_07522_),
    .B(_07174_),
    .A_N(_07517_));
 sg13g2_nand2b_1 _21104_ (.Y(_07523_),
    .B(_07344_),
    .A_N(net7614));
 sg13g2_a21oi_1 _21105_ (.A1(_07522_),
    .A2(_07523_),
    .Y(_07524_),
    .B1(net7396));
 sg13g2_nor2_1 _21106_ (.A(_07132_),
    .B(_07227_),
    .Y(_07525_));
 sg13g2_nand2_1 _21107_ (.Y(_07526_),
    .A(_07116_),
    .B(net7615));
 sg13g2_a21oi_1 _21108_ (.A1(_07483_),
    .A2(_07526_),
    .Y(_07527_),
    .B1(net7392));
 sg13g2_a21oi_1 _21109_ (.A1(_07130_),
    .A2(net7615),
    .Y(_07528_),
    .B1(_07527_));
 sg13g2_o21ai_1 _21110_ (.B1(_07528_),
    .Y(_07529_),
    .A1(_07226_),
    .A2(_07525_));
 sg13g2_mux2_1 _21111_ (.A0(net7615),
    .A1(_07517_),
    .S(_07217_),
    .X(_07530_));
 sg13g2_a21oi_1 _21112_ (.A1(_07149_),
    .A2(_07530_),
    .Y(_07531_),
    .B1(_07529_));
 sg13g2_a21oi_1 _21113_ (.A1(net7396),
    .A2(_07531_),
    .Y(_07532_),
    .B1(_07524_));
 sg13g2_a21oi_1 _21114_ (.A1(net7409),
    .A2(_07532_),
    .Y(_07533_),
    .B1(_07521_));
 sg13g2_a21oi_1 _21115_ (.A1(net5948),
    .A2(_07533_),
    .Y(_07534_),
    .B1(_07512_));
 sg13g2_nor2_1 _21116_ (.A(net7900),
    .B(net5948),
    .Y(_07535_));
 sg13g2_xnor2_1 _21117_ (.Y(_07536_),
    .A(net7397),
    .B(_07128_));
 sg13g2_nand3_1 _21118_ (.B(_07139_),
    .C(_07493_),
    .A(net7391),
    .Y(_07537_));
 sg13g2_o21ai_1 _21119_ (.B1(_07537_),
    .Y(_07538_),
    .A1(net7413),
    .A2(_07536_));
 sg13g2_a22oi_1 _21120_ (.Y(_07539_),
    .B1(_07538_),
    .B2(net7404),
    .A2(net7305),
    .A1(net7308));
 sg13g2_inv_1 _21121_ (.Y(_07540_),
    .A(_07539_));
 sg13g2_nand3b_1 _21122_ (.B(_07485_),
    .C(net7396),
    .Y(_07541_),
    .A_N(_07219_));
 sg13g2_a21oi_1 _21123_ (.A1(_07141_),
    .A2(net7050),
    .Y(_07542_),
    .B1(_07541_));
 sg13g2_o21ai_1 _21124_ (.B1(_07103_),
    .Y(_07543_),
    .A1(net7396),
    .A2(_07160_));
 sg13g2_nor2_1 _21125_ (.A(_07542_),
    .B(_07543_),
    .Y(_07544_));
 sg13g2_nand2b_1 _21126_ (.Y(_07545_),
    .B(_07172_),
    .A_N(_07159_));
 sg13g2_a221oi_1 _21127_ (.B2(net7401),
    .C1(_07544_),
    .B1(_07545_),
    .A1(net7613),
    .Y(_07546_),
    .A2(_07540_));
 sg13g2_a21oi_1 _21128_ (.A1(net5948),
    .A2(_07546_),
    .Y(_07547_),
    .B1(_07535_));
 sg13g2_a21oi_1 _21129_ (.A1(_07143_),
    .A2(_07195_),
    .Y(_07548_),
    .B1(_07216_));
 sg13g2_nor3_1 _21130_ (.A(_07150_),
    .B(net7302),
    .C(_07548_),
    .Y(_07549_));
 sg13g2_nand2_1 _21131_ (.Y(_07550_),
    .A(net7621),
    .B(net7050));
 sg13g2_nand3_1 _21132_ (.B(_07485_),
    .C(_07550_),
    .A(net7305),
    .Y(_07551_));
 sg13g2_a21oi_1 _21133_ (.A1(net7306),
    .A2(_07551_),
    .Y(_07552_),
    .B1(_07549_));
 sg13g2_a21oi_1 _21134_ (.A1(net7391),
    .A2(net7302),
    .Y(_07553_),
    .B1(_07552_));
 sg13g2_mux2_1 _21135_ (.A0(_01891_),
    .A1(_07553_),
    .S(net5942),
    .X(_07554_));
 sg13g2_nor2b_1 _21136_ (.A(net7981),
    .B_N(\id_stage_i.controller_i.instr_valid_i ),
    .Y(_07555_));
 sg13g2_a21oi_1 _21137_ (.A1(_07122_),
    .A2(net7393),
    .Y(_07556_),
    .B1(net7303));
 sg13g2_nand2b_1 _21138_ (.Y(_07557_),
    .B(\id_stage_i.controller_i.instr_valid_i ),
    .A_N(\id_stage_i.id_fsm_q ));
 sg13g2_a21oi_1 _21139_ (.A1(_07132_),
    .A2(net7386),
    .Y(_07558_),
    .B1(net7439));
 sg13g2_and2_1 _21140_ (.A(_01897_),
    .B(_01886_),
    .X(_07559_));
 sg13g2_a21oi_1 _21141_ (.A1(_07483_),
    .A2(_07558_),
    .Y(_07560_),
    .B1(_07291_));
 sg13g2_a221oi_1 _21142_ (.B2(net7617),
    .C1(_07560_),
    .B1(_07228_),
    .A1(net7301),
    .Y(_07561_),
    .A2(net7388));
 sg13g2_nand2_1 _21143_ (.Y(_07562_),
    .A(_01897_),
    .B(_01886_));
 sg13g2_a22oi_1 _21144_ (.Y(_07563_),
    .B1(_07561_),
    .B2(net7303),
    .A2(_07556_),
    .A1(net7405));
 sg13g2_nand2_1 _21145_ (.Y(_07564_),
    .A(net5942),
    .B(_07563_));
 sg13g2_o21ai_1 _21146_ (.B1(_07564_),
    .Y(_07565_),
    .A1(_09282_),
    .A2(net5942));
 sg13g2_nor2_1 _21147_ (.A(_01889_),
    .B(net5946),
    .Y(_07566_));
 sg13g2_nor2_1 _21148_ (.A(_01911_),
    .B(_01908_),
    .Y(_07567_));
 sg13g2_a21oi_1 _21149_ (.A1(net7409),
    .A2(_07160_),
    .Y(_07568_),
    .B1(net7408));
 sg13g2_nor3_1 _21150_ (.A(_07121_),
    .B(net7387),
    .C(_07568_),
    .Y(_07569_));
 sg13g2_or2_1 _21151_ (.X(_07570_),
    .B(_01908_),
    .A(_01911_));
 sg13g2_a22oi_1 _21152_ (.Y(_07571_),
    .B1(_07345_),
    .B2(net7307),
    .A2(net7389),
    .A1(net7397));
 sg13g2_nor2_1 _21153_ (.A(net7409),
    .B(_07571_),
    .Y(_07572_));
 sg13g2_o21ai_1 _21154_ (.B1(net7408),
    .Y(_07573_),
    .A1(_07130_),
    .A2(_07484_));
 sg13g2_a21oi_1 _21155_ (.A1(net7620),
    .A2(net7618),
    .Y(_07574_),
    .B1(_07216_));
 sg13g2_nand2_1 _21156_ (.Y(_07575_),
    .A(_07559_),
    .B(net7609));
 sg13g2_o21ai_1 _21157_ (.B1(_07195_),
    .Y(_07576_),
    .A1(net7407),
    .A2(_07574_));
 sg13g2_a22oi_1 _21158_ (.Y(_07577_),
    .B1(_07576_),
    .B2(_07160_),
    .A2(_07228_),
    .A1(net7619));
 sg13g2_a21oi_1 _21159_ (.A1(_07573_),
    .A2(_07577_),
    .Y(_07578_),
    .B1(net7302));
 sg13g2_nor3_1 _21160_ (.A(_07569_),
    .B(_07572_),
    .C(_07578_),
    .Y(_07579_));
 sg13g2_a21oi_1 _21161_ (.A1(net5946),
    .A2(_07579_),
    .Y(_07580_),
    .B1(_07566_));
 sg13g2_a21oi_1 _21162_ (.A1(net7389),
    .A2(net7612),
    .Y(_07581_),
    .B1(net7399));
 sg13g2_nor2_1 _21163_ (.A(net7393),
    .B(net7302),
    .Y(_07582_));
 sg13g2_o21ai_1 _21164_ (.B1(_07582_),
    .Y(_07583_),
    .A1(net7408),
    .A2(_07581_));
 sg13g2_and3_1 _21165_ (.X(_07584_),
    .A(net7412),
    .B(_07146_),
    .C(_07160_));
 sg13g2_o21ai_1 _21166_ (.B1(net7307),
    .Y(_07585_),
    .A1(_07330_),
    .A2(_07584_));
 sg13g2_nand4_1 _21167_ (.B(net7611),
    .C(_07583_),
    .A(net5944),
    .Y(_07586_),
    .D(_07585_));
 sg13g2_and2_1 _21168_ (.A(_01914_),
    .B(_01913_),
    .X(_07587_));
 sg13g2_o21ai_1 _21169_ (.B1(_07586_),
    .Y(_07588_),
    .A1(_09373_),
    .A2(net5950));
 sg13g2_nor2_1 _21170_ (.A(_07121_),
    .B(_07151_),
    .Y(_07589_));
 sg13g2_nand2_1 _21171_ (.Y(_07590_),
    .A(net7672),
    .B(_01913_));
 sg13g2_a21oi_1 _21172_ (.A1(_07121_),
    .A2(net7612),
    .Y(_07591_),
    .B1(_07589_));
 sg13g2_nor2_1 _21173_ (.A(net7395),
    .B(_07330_),
    .Y(_07592_));
 sg13g2_nand3b_1 _21174_ (.B(_01913_),
    .C(net7672),
    .Y(_07593_),
    .A_N(net7675));
 sg13g2_a21oi_1 _21175_ (.A1(net7404),
    .A2(_07131_),
    .Y(_07594_),
    .B1(net7413));
 sg13g2_nor2_1 _21176_ (.A(_07575_),
    .B(net7608),
    .Y(_07595_));
 sg13g2_nor3_1 _21177_ (.A(_07157_),
    .B(_07592_),
    .C(_07594_),
    .Y(_07596_));
 sg13g2_nor2_1 _21178_ (.A(net7612),
    .B(_07596_),
    .Y(_07597_));
 sg13g2_a221oi_1 _21179_ (.B2(net7412),
    .C1(_07597_),
    .B1(_07591_),
    .A1(net7303),
    .Y(_07598_),
    .A2(net7301));
 sg13g2_or2_1 _21180_ (.X(_07599_),
    .B(net7608),
    .A(_07575_));
 sg13g2_mux2_1 _21181_ (.A0(net7932),
    .A1(_07598_),
    .S(net5950),
    .X(_07600_));
 sg13g2_a21oi_1 _21182_ (.A1(net7408),
    .A2(_07139_),
    .Y(_07601_),
    .B1(_07175_));
 sg13g2_nor4_1 _21183_ (.A(_07557_),
    .B(_07562_),
    .C(_07570_),
    .D(_07593_),
    .Y(_07602_));
 sg13g2_mux2_1 _21184_ (.A0(_01886_),
    .A1(_07601_),
    .S(net5943),
    .X(_07603_));
 sg13g2_mux2_1 _21185_ (.A0(_01885_),
    .A1(net7616),
    .S(net5950),
    .X(_07604_));
 sg13g2_nand2_1 _21186_ (.Y(_07605_),
    .A(_07555_),
    .B(_07595_));
 sg13g2_mux2_1 _21187_ (.A0(_01884_),
    .A1(net7614),
    .S(net5946),
    .X(_07606_));
 sg13g2_mux2_1 _21188_ (.A0(_01883_),
    .A1(net7613),
    .S(net5949),
    .X(_07607_));
 sg13g2_nor2b_1 _21189_ (.A(net7672),
    .B_N(net7675),
    .Y(_07608_));
 sg13g2_mux2_1 _21190_ (.A0(_01882_),
    .A1(net7620),
    .S(net5949),
    .X(_07609_));
 sg13g2_mux2_1 _21191_ (.A0(_01881_),
    .A1(net7618),
    .S(net5951),
    .X(_07610_));
 sg13g2_mux2_1 _21192_ (.A0(_01880_),
    .A1(net7621),
    .S(net5951),
    .X(_07611_));
 sg13g2_mux2_1 _21193_ (.A0(_01879_),
    .A1(net7617),
    .S(net5951),
    .X(_07612_));
 sg13g2_mux2_1 _21194_ (.A0(_01878_),
    .A1(net7619),
    .S(net5944),
    .X(_07613_));
 sg13g2_nand3_1 _21195_ (.B(net7609),
    .C(_07608_),
    .A(net7610),
    .Y(_07614_));
 sg13g2_mux2_1 _21196_ (.A0(_01877_),
    .A1(net7412),
    .S(net5944),
    .X(_07615_));
 sg13g2_and4_1 _21197_ (.A(_01913_),
    .B(_07559_),
    .C(_07567_),
    .D(_07608_),
    .X(_07616_));
 sg13g2_mux2_1 _21198_ (.A0(_01876_),
    .A1(net7401),
    .S(net5952),
    .X(_07617_));
 sg13g2_mux2_1 _21199_ (.A0(_01875_),
    .A1(net7393),
    .S(net5952),
    .X(_07618_));
 sg13g2_nand4_1 _21200_ (.B(_07559_),
    .C(_07567_),
    .A(net7674),
    .Y(_07619_),
    .D(_07608_));
 sg13g2_mux2_1 _21201_ (.A0(_01874_),
    .A1(net7408),
    .S(net5944),
    .X(_07620_));
 sg13g2_mux2_1 _21202_ (.A0(_01873_),
    .A1(net7388),
    .S(net5944),
    .X(_07621_));
 sg13g2_inv_1 _21203_ (.Y(_07622_),
    .A(_01942_));
 sg13g2_mux2_1 _21204_ (.A0(_01872_),
    .A1(net7611),
    .S(net5950),
    .X(_07623_));
 sg13g2_mux2_1 _21205_ (.A0(_01871_),
    .A1(net7612),
    .S(net5952),
    .X(_07624_));
 sg13g2_mux2_1 _21206_ (.A0(_01870_),
    .A1(net7398),
    .S(net5952),
    .X(_07625_));
 sg13g2_mux2_1 _21207_ (.A0(net7933),
    .A1(_07172_),
    .S(net5950),
    .X(_07626_));
 sg13g2_nor2b_1 _21208_ (.A(net7956),
    .B_N(net383),
    .Y(_07627_));
 sg13g2_nor2b_1 _21209_ (.A(_01836_),
    .B_N(_01835_),
    .Y(_07628_));
 sg13g2_a22oi_1 _21210_ (.Y(_07629_),
    .B1(_07628_),
    .B2(net383),
    .A2(_01706_),
    .A1(_01836_));
 sg13g2_nor4_1 _21211_ (.A(_15152_),
    .B(_01705_),
    .C(net5922),
    .D(_07629_),
    .Y(_07630_));
 sg13g2_a21o_1 _21212_ (.A2(net5922),
    .A1(\id_stage_i.controller_i.instr_fetch_err_plus2_i ),
    .B1(_07630_),
    .X(_07631_));
 sg13g2_nand2_1 _21213_ (.Y(_07632_),
    .A(_01836_),
    .B(net7976));
 sg13g2_nand3_1 _21214_ (.B(_01746_),
    .C(net7976),
    .A(_01747_),
    .Y(_07633_));
 sg13g2_nand2_1 _21215_ (.Y(_07634_),
    .A(_01835_),
    .B(_07633_));
 sg13g2_nor3_1 _21216_ (.A(_01910_),
    .B(_01907_),
    .C(_01906_),
    .Y(_07635_));
 sg13g2_a22oi_1 _21217_ (.Y(_07636_),
    .B1(_07634_),
    .B2(net383),
    .A2(_01705_),
    .A1(_01835_));
 sg13g2_a21oi_1 _21218_ (.A1(_01706_),
    .A2(_07012_),
    .Y(_07637_),
    .B1(_01705_));
 sg13g2_nor2b_1 _21219_ (.A(_07632_),
    .B_N(_07637_),
    .Y(_07638_));
 sg13g2_a21oi_1 _21220_ (.A1(_07632_),
    .A2(_07636_),
    .Y(_07639_),
    .B1(_07638_));
 sg13g2_nand2_1 _21221_ (.Y(_07640_),
    .A(net5941),
    .B(_07639_));
 sg13g2_o21ai_1 _21222_ (.B1(_07640_),
    .Y(_07641_),
    .A1(_10165_),
    .A2(net5941));
 sg13g2_a21oi_1 _21223_ (.A1(net7439),
    .A2(net7611),
    .Y(_07642_),
    .B1(_07150_));
 sg13g2_nor2_1 _21224_ (.A(net7389),
    .B(_07226_),
    .Y(_07643_));
 sg13g2_nor3_1 _21225_ (.A(_01905_),
    .B(_01904_),
    .C(_01903_),
    .Y(_07644_));
 sg13g2_a22oi_1 _21226_ (.Y(_07645_),
    .B1(_07643_),
    .B2(_07146_),
    .A2(_07642_),
    .A1(net7389));
 sg13g2_nand2b_1 _21227_ (.Y(_07646_),
    .B(net7303),
    .A_N(_07645_));
 sg13g2_a21oi_1 _21228_ (.A1(net7393),
    .A2(_07205_),
    .Y(_07647_),
    .B1(_07484_));
 sg13g2_o21ai_1 _21229_ (.B1(net7405),
    .Y(_07648_),
    .A1(net7401),
    .A2(_07647_));
 sg13g2_and2_1 _21230_ (.A(_07635_),
    .B(_07644_),
    .X(_07649_));
 sg13g2_nor4_1 _21231_ (.A(net7413),
    .B(net7396),
    .C(_07143_),
    .D(_07344_),
    .Y(_07650_));
 sg13g2_or2_1 _21232_ (.X(_07651_),
    .B(_07650_),
    .A(_07153_));
 sg13g2_and2_1 _21233_ (.A(net7386),
    .B(_07205_),
    .X(_07652_));
 sg13g2_a221oi_1 _21234_ (.B2(_07652_),
    .C1(_07175_),
    .B1(_07651_),
    .A1(net7411),
    .Y(_07653_),
    .A2(_07648_));
 sg13g2_o21ai_1 _21235_ (.B1(_07646_),
    .Y(_07654_),
    .A1(net7398),
    .A2(_07653_));
 sg13g2_nor2_1 _21236_ (.A(net7927),
    .B(net7930),
    .Y(_07655_));
 sg13g2_mux2_1 _21237_ (.A0(\id_stage_i.decoder_i.illegal_c_insn_i ),
    .A1(_07654_),
    .S(net5942),
    .X(_07656_));
 sg13g2_or2_1 _21238_ (.X(_07657_),
    .B(_01600_),
    .A(_01605_));
 sg13g2_nor2_1 _21239_ (.A(\id_stage_i.controller_i.nmi_mode_d ),
    .B(_07657_),
    .Y(_07658_));
 sg13g2_or2_1 _21240_ (.X(_07659_),
    .B(_07657_),
    .A(\id_stage_i.controller_i.nmi_mode_d ));
 sg13g2_nor2_1 _21241_ (.A(\id_stage_i.controller_i.controller_run_o ),
    .B(_07659_),
    .Y(_07660_));
 sg13g2_nand2_1 _21242_ (.Y(_07661_),
    .A(_02232_),
    .B(_07658_));
 sg13g2_nor2_1 _21243_ (.A(_01603_),
    .B(_07661_),
    .Y(_07662_));
 sg13g2_nor2_1 _21244_ (.A(_01604_),
    .B(_01601_),
    .Y(_07663_));
 sg13g2_a21oi_1 _21245_ (.A1(_07662_),
    .A2(_07663_),
    .Y(_07664_),
    .B1(_01839_));
 sg13g2_nand2_1 _21246_ (.Y(_07665_),
    .A(_01909_),
    .B(_09244_));
 sg13g2_o21ai_1 _21247_ (.B1(_01836_),
    .Y(_07666_),
    .A1(_01838_),
    .A2(_01837_));
 sg13g2_o21ai_1 _21248_ (.B1(_07664_),
    .Y(_07667_),
    .A1(net6762),
    .A2(_07666_));
 sg13g2_and2_1 _21249_ (.A(net7455),
    .B(_07667_),
    .X(_07668_));
 sg13g2_inv_1 _21250_ (.Y(net538),
    .A(_07668_));
 sg13g2_nor3_1 _21251_ (.A(net7926),
    .B(net7931),
    .C(_07665_),
    .Y(_07669_));
 sg13g2_nor2_1 _21252_ (.A(net384),
    .B(_07668_),
    .Y(_07670_));
 sg13g2_nor3_1 _21253_ (.A(_02232_),
    .B(_07085_),
    .C(_07659_),
    .Y(_07671_));
 sg13g2_nor2_1 _21254_ (.A(_02238_),
    .B(_06896_),
    .Y(_07672_));
 sg13g2_nand2_1 _21255_ (.Y(_07673_),
    .A(net7985),
    .B(_06897_));
 sg13g2_a21oi_1 _21256_ (.A1(_01603_),
    .A2(_06965_),
    .Y(_07674_),
    .B1(_07658_));
 sg13g2_nor2_1 _21257_ (.A(net7437),
    .B(_07674_),
    .Y(_07675_));
 sg13g2_nor2_1 _21258_ (.A(\id_stage_i.controller_i.controller_run_o ),
    .B(_07675_),
    .Y(_07676_));
 sg13g2_o21ai_1 _21259_ (.B1(_02232_),
    .Y(_07677_),
    .A1(net7437),
    .A2(_07674_));
 sg13g2_a21o_1 _21260_ (.A2(_07672_),
    .A1(\cs_registers_i.debug_mode_i ),
    .B1(_07657_),
    .X(_07678_));
 sg13g2_nor2_1 _21261_ (.A(_07677_),
    .B(_07678_),
    .Y(_07679_));
 sg13g2_nand2_1 _21262_ (.Y(_07680_),
    .A(_01890_),
    .B(net7929));
 sg13g2_nor2_1 _21263_ (.A(_02232_),
    .B(net7626),
    .Y(_07681_));
 sg13g2_a21oi_1 _21264_ (.A1(net7313),
    .A2(_06896_),
    .Y(_07682_),
    .B1(_07681_));
 sg13g2_inv_1 _21265_ (.Y(_07683_),
    .A(_07684_));
 sg13g2_nand2_1 _21266_ (.Y(_07684_),
    .A(net7986),
    .B(net7105));
 sg13g2_nand3_1 _21267_ (.B(_07659_),
    .C(_07684_),
    .A(\id_stage_i.controller_i.controller_run_o ),
    .Y(_07685_));
 sg13g2_o21ai_1 _21268_ (.B1(_07685_),
    .Y(_07686_),
    .A1(_02238_),
    .A2(_07682_));
 sg13g2_nand2_1 _21269_ (.Y(_07687_),
    .A(_00381_),
    .B(net6927));
 sg13g2_nor2_1 _21270_ (.A(net7313),
    .B(_07661_),
    .Y(_07688_));
 sg13g2_o21ai_1 _21271_ (.B1(_07684_),
    .Y(_07689_),
    .A1(net7313),
    .A2(_07661_));
 sg13g2_a21o_1 _21272_ (.A2(_07689_),
    .A1(net7626),
    .B1(_07662_),
    .X(_07690_));
 sg13g2_and2_1 _21273_ (.A(net7986),
    .B(_06896_),
    .X(_07691_));
 sg13g2_nand2_1 _21274_ (.Y(_07692_),
    .A(net7985),
    .B(_06896_));
 sg13g2_nand2_1 _21275_ (.Y(_07693_),
    .A(net7105),
    .B(_07691_));
 sg13g2_nor2_1 _21276_ (.A(_09282_),
    .B(net7931),
    .Y(_07694_));
 sg13g2_nor2_1 _21277_ (.A(_07661_),
    .B(_07693_),
    .Y(_07695_));
 sg13g2_nand3_1 _21278_ (.B(_07660_),
    .C(_07691_),
    .A(net7105),
    .Y(_07696_));
 sg13g2_nand2b_1 _21279_ (.Y(_07697_),
    .B(_07688_),
    .A_N(net7105));
 sg13g2_nand2_1 _21280_ (.Y(_07698_),
    .A(net7928),
    .B(_09324_));
 sg13g2_o21ai_1 _21281_ (.B1(net6923),
    .Y(_07699_),
    .A1(_00279_),
    .A2(net7047));
 sg13g2_nand2_1 _21282_ (.Y(_07700_),
    .A(_07687_),
    .B(_07699_));
 sg13g2_nand2b_1 _21283_ (.Y(_07701_),
    .B(net7929),
    .A_N(_01890_));
 sg13g2_a221oi_1 _21284_ (.B2(_00530_),
    .C1(_07700_),
    .B1(net6881),
    .A1(net469),
    .Y(_07702_),
    .A2(net6884));
 sg13g2_o21ai_1 _21285_ (.B1(_07697_),
    .Y(_07703_),
    .A1(_07684_),
    .A2(_07688_));
 sg13g2_a21oi_1 _21286_ (.A1(net7626),
    .A2(_07703_),
    .Y(_07704_),
    .B1(_07662_));
 sg13g2_nor2_1 _21287_ (.A(net313),
    .B(net6922),
    .Y(_07705_));
 sg13g2_nor2_1 _21288_ (.A(_07702_),
    .B(_07705_),
    .Y(_07706_));
 sg13g2_nand2_1 _21289_ (.Y(_07707_),
    .A(net6760),
    .B(_07706_));
 sg13g2_nand2_1 _21290_ (.Y(_07708_),
    .A(_07698_),
    .B(_07701_));
 sg13g2_o21ai_1 _21291_ (.B1(_07707_),
    .Y(_07709_),
    .A1(_15492_),
    .A2(net6761));
 sg13g2_mux2_1 _21292_ (.A0(_01869_),
    .A1(_07709_),
    .S(net7454),
    .X(net537));
 sg13g2_nor2_1 _21293_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .B(_07667_),
    .Y(_07710_));
 sg13g2_nand2b_1 _21294_ (.Y(_07711_),
    .B(_10215_),
    .A_N(_07667_));
 sg13g2_nor2_1 _21295_ (.A(net384),
    .B(_07711_),
    .Y(_07712_));
 sg13g2_mux2_1 _21296_ (.A0(_01869_),
    .A1(net537),
    .S(net6648),
    .X(_07713_));
 sg13g2_nand2_1 _21297_ (.Y(_07714_),
    .A(_01703_),
    .B(net6775));
 sg13g2_nor2_1 _21298_ (.A(net312),
    .B(_07704_),
    .Y(_07715_));
 sg13g2_nor2_1 _21299_ (.A(_00278_),
    .B(_07661_),
    .Y(_07716_));
 sg13g2_o21ai_1 _21300_ (.B1(_07697_),
    .Y(_07717_),
    .A1(_07684_),
    .A2(_07716_));
 sg13g2_a221oi_1 _21301_ (.B2(net7626),
    .C1(_07662_),
    .B1(_07717_),
    .A1(_00380_),
    .Y(_07718_),
    .A2(_07686_));
 sg13g2_inv_1 _21302_ (.Y(_07719_),
    .A(_07718_));
 sg13g2_a221oi_1 _21303_ (.B2(_00529_),
    .C1(_07719_),
    .B1(_07679_),
    .A1(net468),
    .Y(_07720_),
    .A2(net6885));
 sg13g2_nor2_1 _21304_ (.A(_07715_),
    .B(_07720_),
    .Y(_07721_));
 sg13g2_nand2_1 _21305_ (.Y(_07722_),
    .A(net6762),
    .B(_07721_));
 sg13g2_and2_1 _21306_ (.A(_07714_),
    .B(_07722_),
    .X(_07723_));
 sg13g2_nand2_1 _21307_ (.Y(_07724_),
    .A(_07714_),
    .B(_07722_));
 sg13g2_mux2_1 _21308_ (.A0(_01868_),
    .A1(_07724_),
    .S(net7454),
    .X(net536));
 sg13g2_mux2_1 _21309_ (.A0(_01868_),
    .A1(net536),
    .S(net6648),
    .X(_07725_));
 sg13g2_nand2_1 _21310_ (.Y(_07726_),
    .A(_00379_),
    .B(_07686_));
 sg13g2_o21ai_1 _21311_ (.B1(_07690_),
    .Y(_07727_),
    .A1(_00277_),
    .A2(_07696_));
 sg13g2_nand3_1 _21312_ (.B(_07726_),
    .C(_07727_),
    .A(net6768),
    .Y(_07728_));
 sg13g2_a21oi_1 _21313_ (.A1(net467),
    .A2(net6885),
    .Y(_07729_),
    .B1(_07728_));
 sg13g2_a21oi_1 _21314_ (.A1(_15523_),
    .A2(net6776),
    .Y(_07730_),
    .B1(_07729_));
 sg13g2_mux2_1 _21315_ (.A0(_01867_),
    .A1(_07730_),
    .S(net7454),
    .X(net535));
 sg13g2_mux2_1 _21316_ (.A0(_01867_),
    .A1(net535),
    .S(net6648),
    .X(_07731_));
 sg13g2_nand2_1 _21317_ (.Y(_07732_),
    .A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .B(_01866_));
 sg13g2_nor3_1 _21318_ (.A(_07657_),
    .B(net7437),
    .C(_07677_),
    .Y(_07733_));
 sg13g2_nand2_1 _21319_ (.Y(_07734_),
    .A(net434),
    .B(_02211_));
 sg13g2_a21oi_1 _21320_ (.A1(_06998_),
    .A2(_07734_),
    .Y(_07735_),
    .B1(_07088_));
 sg13g2_nand2_1 _21321_ (.Y(_07736_),
    .A(_07733_),
    .B(_07735_));
 sg13g2_a22oi_1 _21322_ (.Y(_07737_),
    .B1(_07695_),
    .B2(_00276_),
    .A2(net6929),
    .A1(_00378_));
 sg13g2_nand3_1 _21323_ (.B(_07736_),
    .C(_07737_),
    .A(net6768),
    .Y(_07738_));
 sg13g2_nand2b_1 _21324_ (.Y(_07739_),
    .B(net7930),
    .A_N(net7921));
 sg13g2_a21oi_1 _21325_ (.A1(net466),
    .A2(net6886),
    .Y(_07740_),
    .B1(_07738_));
 sg13g2_a21oi_1 _21326_ (.A1(_15529_),
    .A2(net6776),
    .Y(_07741_),
    .B1(_07740_));
 sg13g2_inv_1 _21327_ (.Y(_07742_),
    .A(_07741_));
 sg13g2_o21ai_1 _21328_ (.B1(_07732_),
    .Y(net534),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .A2(_07742_));
 sg13g2_mux2_1 _21329_ (.A0(_01866_),
    .A1(net534),
    .S(_07712_),
    .X(_07743_));
 sg13g2_and2_1 _21330_ (.A(net6762),
    .B(_07704_),
    .X(_07744_));
 sg13g2_a21o_1 _21331_ (.A2(_07739_),
    .A1(_08711_),
    .B1(_09282_),
    .X(_07745_));
 sg13g2_nand2b_1 _21332_ (.Y(_07746_),
    .B(_07734_),
    .A_N(_06997_));
 sg13g2_nor2_1 _21333_ (.A(_06989_),
    .B(_06999_),
    .Y(_07747_));
 sg13g2_nor3_1 _21334_ (.A(_06993_),
    .B(_07746_),
    .C(_07747_),
    .Y(_07748_));
 sg13g2_nor3_1 _21335_ (.A(net7734),
    .B(net7748),
    .C(_08306_),
    .Y(_07749_));
 sg13g2_nand3b_1 _21336_ (.B(net7437),
    .C(_07749_),
    .Y(_07750_),
    .A_N(_06904_));
 sg13g2_o21ai_1 _21337_ (.B1(_07750_),
    .Y(_07751_),
    .A1(_07088_),
    .A2(_07748_));
 sg13g2_a22oi_1 _21338_ (.Y(_07752_),
    .B1(_07686_),
    .B2(_00377_),
    .A2(_07671_),
    .A1(net465));
 sg13g2_o21ai_1 _21339_ (.B1(_07752_),
    .Y(_07753_),
    .A1(_06067_),
    .A2(_07696_));
 sg13g2_a21o_1 _21340_ (.A2(_07751_),
    .A1(_07733_),
    .B1(_07753_),
    .X(_07754_));
 sg13g2_and2_1 _21341_ (.A(_01700_),
    .B(net6776),
    .X(_07755_));
 sg13g2_a21o_1 _21342_ (.A2(_07754_),
    .A1(_07744_),
    .B1(_07755_),
    .X(_07756_));
 sg13g2_xnor2_1 _21343_ (.Y(_07757_),
    .A(net7921),
    .B(net7930));
 sg13g2_mux2_1 _21344_ (.A0(_01865_),
    .A1(_07756_),
    .S(net7454),
    .X(net533));
 sg13g2_mux2_1 _21345_ (.A0(_01865_),
    .A1(net533),
    .S(net6648),
    .X(_07758_));
 sg13g2_nor2_1 _21346_ (.A(_06984_),
    .B(_06993_),
    .Y(_07759_));
 sg13g2_or3_1 _21347_ (.A(_07001_),
    .B(_07746_),
    .C(_07759_),
    .X(_07760_));
 sg13g2_nor2b_1 _21348_ (.A(_06782_),
    .B_N(_06903_),
    .Y(_07761_));
 sg13g2_nor2b_1 _21349_ (.A(_06895_),
    .B_N(_07761_),
    .Y(_07762_));
 sg13g2_a22oi_1 _21350_ (.Y(_07763_),
    .B1(_07762_),
    .B2(net7985),
    .A2(_07760_),
    .A1(_07087_));
 sg13g2_nand2b_1 _21351_ (.Y(_07764_),
    .B(_07733_),
    .A_N(_07763_));
 sg13g2_a22oi_1 _21352_ (.Y(_07765_),
    .B1(_07695_),
    .B2(_00274_),
    .A2(net6929),
    .A1(_00376_));
 sg13g2_nand3_1 _21353_ (.B(_07764_),
    .C(_07765_),
    .A(net6768),
    .Y(_07766_));
 sg13g2_a21oi_1 _21354_ (.A1(net464),
    .A2(net6886),
    .Y(_07767_),
    .B1(_07766_));
 sg13g2_a21oi_1 _21355_ (.A1(_15536_),
    .A2(net6776),
    .Y(_07768_),
    .B1(_07767_));
 sg13g2_mux2_1 _21356_ (.A0(_01864_),
    .A1(_07768_),
    .S(net7454),
    .X(net532));
 sg13g2_mux2_1 _21357_ (.A0(_01864_),
    .A1(net532),
    .S(net6647),
    .X(_07769_));
 sg13g2_nand2_1 _21358_ (.Y(_07770_),
    .A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .B(_01863_));
 sg13g2_a22oi_1 _21359_ (.Y(_07771_),
    .B1(_07749_),
    .B2(_06777_),
    .A2(_06900_),
    .A1(_10463_));
 sg13g2_or2_1 _21360_ (.X(_07772_),
    .B(_07771_),
    .A(_06904_));
 sg13g2_nor2b_1 _21361_ (.A(_06782_),
    .B_N(\id_stage_i.controller_i.store_err_q ),
    .Y(_07773_));
 sg13g2_o21ai_1 _21362_ (.B1(_06902_),
    .Y(_07774_),
    .A1(\id_stage_i.controller_i.illegal_insn_q ),
    .A2(_07773_));
 sg13g2_a221oi_1 _21363_ (.B2(_07774_),
    .C1(_07673_),
    .B1(_07772_),
    .A1(_06895_),
    .Y(_07775_),
    .A2(_07761_));
 sg13g2_o21ai_1 _21364_ (.B1(_06981_),
    .Y(_07776_),
    .A1(_06983_),
    .A2(_06987_));
 sg13g2_nand2_1 _21365_ (.Y(_07777_),
    .A(_06990_),
    .B(_07776_));
 sg13g2_nand2_1 _21366_ (.Y(_07778_),
    .A(_06992_),
    .B(_07777_));
 sg13g2_nand2_1 _21367_ (.Y(_07779_),
    .A(_06996_),
    .B(_07778_));
 sg13g2_nor2_1 _21368_ (.A(_01891_),
    .B(_01890_),
    .Y(_07780_));
 sg13g2_nor2b_1 _21369_ (.A(_06998_),
    .B_N(_07734_),
    .Y(_07781_));
 sg13g2_nand3_1 _21370_ (.B(_07779_),
    .C(_07781_),
    .A(_06995_),
    .Y(_07782_));
 sg13g2_or2_1 _21371_ (.X(_07783_),
    .B(net7927),
    .A(net7921));
 sg13g2_a21oi_1 _21372_ (.A1(_07087_),
    .A2(_07782_),
    .Y(_07784_),
    .B1(_07775_));
 sg13g2_nand2b_1 _21373_ (.Y(_07785_),
    .B(_07733_),
    .A_N(_07784_));
 sg13g2_nand2_1 _21374_ (.Y(_07786_),
    .A(_06896_),
    .B(_07657_));
 sg13g2_o21ai_1 _21375_ (.B1(_07786_),
    .Y(_07787_),
    .A1(_02226_),
    .A2(_06896_));
 sg13g2_nand3_1 _21376_ (.B(_07676_),
    .C(_07787_),
    .A(net7985),
    .Y(_07788_));
 sg13g2_a22oi_1 _21377_ (.Y(_07789_),
    .B1(_07695_),
    .B2(_00273_),
    .A2(net6929),
    .A1(_00375_));
 sg13g2_nor3_1 _21378_ (.A(net7925),
    .B(_01890_),
    .C(net7931),
    .Y(_07790_));
 sg13g2_nand4_1 _21379_ (.B(_07785_),
    .C(_07788_),
    .A(net6768),
    .Y(_07791_),
    .D(_07789_));
 sg13g2_or3_1 _21380_ (.A(net7925),
    .B(net7926),
    .C(net7931),
    .X(_07792_));
 sg13g2_a21oi_1 _21381_ (.A1(net463),
    .A2(net6886),
    .Y(_07793_),
    .B1(_07791_));
 sg13g2_a21oi_1 _21382_ (.A1(_15542_),
    .A2(_07092_),
    .Y(_07794_),
    .B1(_07793_));
 sg13g2_inv_1 _21383_ (.Y(_07795_),
    .A(_07794_));
 sg13g2_o21ai_1 _21384_ (.B1(_07770_),
    .Y(net531),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .A2(_07795_));
 sg13g2_mux2_1 _21385_ (.A0(_01863_),
    .A1(net531),
    .S(_07712_),
    .X(_07796_));
 sg13g2_nand2_1 _21386_ (.Y(_07797_),
    .A(_00374_),
    .B(net6926));
 sg13g2_o21ai_1 _21387_ (.B1(net6923),
    .Y(_07798_),
    .A1(_00272_),
    .A2(net7047));
 sg13g2_nand2_1 _21388_ (.Y(_07799_),
    .A(_07797_),
    .B(_07798_));
 sg13g2_mux2_1 _21389_ (.A0(_07757_),
    .A1(_07792_),
    .S(_08711_),
    .X(_07800_));
 sg13g2_a221oi_1 _21390_ (.B2(_00528_),
    .C1(_07799_),
    .B1(net6881),
    .A1(net6567),
    .Y(_07801_),
    .A2(net6884));
 sg13g2_o21ai_1 _21391_ (.B1(net6764),
    .Y(_07802_),
    .A1(net311),
    .A2(net6922));
 sg13g2_or2_1 _21392_ (.X(_07803_),
    .B(_07802_),
    .A(_07801_));
 sg13g2_nand2_1 _21393_ (.Y(_07804_),
    .A(_01697_),
    .B(net6774));
 sg13g2_a21oi_1 _21394_ (.A1(_01697_),
    .A2(net6774),
    .Y(_07805_),
    .B1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ));
 sg13g2_nand3_1 _21395_ (.B(_07745_),
    .C(_07800_),
    .A(_07649_),
    .Y(_07806_));
 sg13g2_nor3_1 _21396_ (.A(_01909_),
    .B(net7682),
    .C(_01904_),
    .Y(_07807_));
 sg13g2_a22oi_1 _21397_ (.Y(net530),
    .B1(_07803_),
    .B2(_07805_),
    .A2(_10417_),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ));
 sg13g2_nand2_1 _21398_ (.Y(_07808_),
    .A(net6648),
    .B(net530));
 sg13g2_o21ai_1 _21399_ (.B1(_07808_),
    .Y(_07809_),
    .A1(_10417_),
    .A2(net6648));
 sg13g2_nand2_1 _21400_ (.Y(_07810_),
    .A(_00373_),
    .B(net6926));
 sg13g2_o21ai_1 _21401_ (.B1(net6923),
    .Y(_07811_),
    .A1(_00271_),
    .A2(net7047));
 sg13g2_and2_1 _21402_ (.A(_07635_),
    .B(_07807_),
    .X(_07812_));
 sg13g2_nand2_1 _21403_ (.Y(_07813_),
    .A(_07810_),
    .B(_07811_));
 sg13g2_a221oi_1 _21404_ (.B2(_00527_),
    .C1(_07813_),
    .B1(net6881),
    .A1(net6570),
    .Y(_07814_),
    .A2(net6884));
 sg13g2_nand2_1 _21405_ (.Y(_07815_),
    .A(_07635_),
    .B(_07807_));
 sg13g2_o21ai_1 _21406_ (.B1(net6764),
    .Y(_07816_),
    .A1(net310),
    .A2(net6921));
 sg13g2_nor2_1 _21407_ (.A(_07814_),
    .B(_07816_),
    .Y(_07817_));
 sg13g2_a21o_1 _21408_ (.A2(net6770),
    .A1(_01696_),
    .B1(_07817_),
    .X(_07818_));
 sg13g2_mux2_1 _21409_ (.A0(_01861_),
    .A1(_07818_),
    .S(net7452),
    .X(net529));
 sg13g2_mux2_1 _21410_ (.A0(_01861_),
    .A1(net529),
    .S(net6646),
    .X(_07819_));
 sg13g2_nor2_1 _21411_ (.A(net7455),
    .B(_01860_),
    .Y(_07820_));
 sg13g2_nand3_1 _21412_ (.B(_00391_),
    .C(_06985_),
    .A(net425),
    .Y(_07821_));
 sg13g2_a22oi_1 _21413_ (.Y(_07822_),
    .B1(_06986_),
    .B2(_07821_),
    .A2(_00394_),
    .A1(net428));
 sg13g2_a21oi_1 _21414_ (.A1(net429),
    .A2(_00395_),
    .Y(_07823_),
    .B1(_07822_));
 sg13g2_a21oi_1 _21415_ (.A1(net430),
    .A2(_00396_),
    .Y(_07824_),
    .B1(_07823_));
 sg13g2_a21oi_1 _21416_ (.A1(net431),
    .A2(_00397_),
    .Y(_07825_),
    .B1(_07824_));
 sg13g2_o21ai_1 _21417_ (.B1(_07812_),
    .Y(_07826_),
    .A1(_01903_),
    .A2(net7607));
 sg13g2_a21oi_1 _21418_ (.A1(net432),
    .A2(_00398_),
    .Y(_07827_),
    .B1(_07825_));
 sg13g2_a21o_1 _21419_ (.A2(_00399_),
    .A1(net433),
    .B1(_07827_),
    .X(_07828_));
 sg13g2_a22oi_1 _21420_ (.Y(_07829_),
    .B1(_06991_),
    .B2(_07828_),
    .A2(_00384_),
    .A1(net421));
 sg13g2_a21oi_1 _21421_ (.A1(net422),
    .A2(_00385_),
    .Y(_07830_),
    .B1(_07829_));
 sg13g2_a21oi_1 _21422_ (.A1(net423),
    .A2(_00386_),
    .Y(_07831_),
    .B1(_07830_));
 sg13g2_o21ai_1 _21423_ (.B1(_07781_),
    .Y(_07832_),
    .A1(_06994_),
    .A2(_07831_));
 sg13g2_or3_1 _21424_ (.A(\id_stage_i.controller_i.illegal_insn_q ),
    .B(_06782_),
    .C(_06895_),
    .X(_07833_));
 sg13g2_and3_1 _21425_ (.X(_07834_),
    .A(_08711_),
    .B(_07635_),
    .C(_07644_));
 sg13g2_nand3_1 _21426_ (.B(_07772_),
    .C(_07833_),
    .A(_06902_),
    .Y(_07835_));
 sg13g2_a22oi_1 _21427_ (.Y(_07836_),
    .B1(_07835_),
    .B2(net7437),
    .A2(_07832_),
    .A1(_07087_));
 sg13g2_inv_1 _21428_ (.Y(_07837_),
    .A(_07836_));
 sg13g2_nand2b_1 _21429_ (.Y(_07838_),
    .B(_07733_),
    .A_N(_07836_));
 sg13g2_a22oi_1 _21430_ (.Y(_07839_),
    .B1(_07695_),
    .B2(_00270_),
    .A2(net6929),
    .A1(_00372_));
 sg13g2_nand2_1 _21431_ (.Y(_07840_),
    .A(_07838_),
    .B(_07839_));
 sg13g2_nor2_1 _21432_ (.A(net7920),
    .B(_09282_),
    .Y(_07841_));
 sg13g2_a21o_1 _21433_ (.A2(net6886),
    .A1(net460),
    .B1(_07840_),
    .X(_07842_));
 sg13g2_nand2_1 _21434_ (.Y(_07843_),
    .A(_07744_),
    .B(_07842_));
 sg13g2_nand2b_1 _21435_ (.Y(_07844_),
    .B(net7927),
    .A_N(net7921));
 sg13g2_a22oi_1 _21436_ (.Y(_07845_),
    .B1(_07744_),
    .B2(_07842_),
    .A2(net6776),
    .A1(_01695_));
 sg13g2_a21oi_1 _21437_ (.A1(net7455),
    .A2(_07845_),
    .Y(net528),
    .B1(_07820_));
 sg13g2_mux2_1 _21438_ (.A0(_01860_),
    .A1(net528),
    .S(net6645),
    .X(_07846_));
 sg13g2_nand2_1 _21439_ (.Y(_07847_),
    .A(_00371_),
    .B(net6926));
 sg13g2_o21ai_1 _21440_ (.B1(net6923),
    .Y(_07848_),
    .A1(_00269_),
    .A2(net7047));
 sg13g2_nand2_1 _21441_ (.Y(_07849_),
    .A(_07847_),
    .B(_07848_));
 sg13g2_nor2_1 _21442_ (.A(net7930),
    .B(_07844_),
    .Y(_07850_));
 sg13g2_a221oi_1 _21443_ (.B2(_00526_),
    .C1(_07849_),
    .B1(net6881),
    .A1(net6571),
    .Y(_07851_),
    .A2(net6884));
 sg13g2_o21ai_1 _21444_ (.B1(net6764),
    .Y(_07852_),
    .A1(net309),
    .A2(net6922));
 sg13g2_nor2_1 _21445_ (.A(_07851_),
    .B(_07852_),
    .Y(_07853_));
 sg13g2_a21o_1 _21446_ (.A2(net6770),
    .A1(_01694_),
    .B1(_07853_),
    .X(_07854_));
 sg13g2_mux2_1 _21447_ (.A0(_01859_),
    .A1(_07854_),
    .S(net7452),
    .X(net527));
 sg13g2_mux2_1 _21448_ (.A0(_01859_),
    .A1(net527),
    .S(net6646),
    .X(_07855_));
 sg13g2_o21ai_1 _21449_ (.B1(_07676_),
    .Y(_07856_),
    .A1(_00525_),
    .A2(_07678_));
 sg13g2_inv_1 _21450_ (.Y(_07857_),
    .A(_07858_));
 sg13g2_o21ai_1 _21451_ (.B1(net6923),
    .Y(_07858_),
    .A1(_00268_),
    .A2(net7047));
 sg13g2_a221oi_1 _21452_ (.B2(_00370_),
    .C1(_07857_),
    .B1(net6927),
    .A1(net6573),
    .Y(_07859_),
    .A2(net6884));
 sg13g2_a21o_1 _21453_ (.A2(_07850_),
    .A1(_07834_),
    .B1(net7683),
    .X(_07860_));
 sg13g2_o21ai_1 _21454_ (.B1(net6764),
    .Y(_07861_),
    .A1(net308),
    .A2(net6921));
 sg13g2_a21oi_1 _21455_ (.A1(_07856_),
    .A2(_07859_),
    .Y(_07862_),
    .B1(_07861_));
 sg13g2_a21o_1 _21456_ (.A2(net6770),
    .A1(_01693_),
    .B1(_07862_),
    .X(_07863_));
 sg13g2_a21o_1 _21457_ (.A2(_07826_),
    .A1(_07806_),
    .B1(_07860_),
    .X(_07864_));
 sg13g2_mux2_1 _21458_ (.A0(_01858_),
    .A1(_07863_),
    .S(net7452),
    .X(net526));
 sg13g2_mux2_1 _21459_ (.A0(_01858_),
    .A1(net526),
    .S(net6646),
    .X(_07865_));
 sg13g2_o21ai_1 _21460_ (.B1(_07676_),
    .Y(_07866_),
    .A1(_00524_),
    .A2(_07678_));
 sg13g2_inv_1 _21461_ (.Y(_07867_),
    .A(_07868_));
 sg13g2_o21ai_1 _21462_ (.B1(net6925),
    .Y(_07868_),
    .A1(_00267_),
    .A2(net7049));
 sg13g2_a221oi_1 _21463_ (.B2(_00369_),
    .C1(_07867_),
    .B1(net6928),
    .A1(net6575),
    .Y(_07869_),
    .A2(net6883));
 sg13g2_nor2_1 _21464_ (.A(net7672),
    .B(_01913_),
    .Y(_07870_));
 sg13g2_o21ai_1 _21465_ (.B1(net6765),
    .Y(_07871_),
    .A1(net307),
    .A2(net6920));
 sg13g2_or2_1 _21466_ (.X(_07872_),
    .B(_01913_),
    .A(_01914_));
 sg13g2_a21o_1 _21467_ (.A2(_07869_),
    .A1(_07866_),
    .B1(_07871_),
    .X(_07873_));
 sg13g2_o21ai_1 _21468_ (.B1(_07873_),
    .Y(_07874_),
    .A1(_15556_),
    .A2(net6767));
 sg13g2_mux2_1 _21469_ (.A0(_01857_),
    .A1(_07874_),
    .S(net7452),
    .X(net525));
 sg13g2_mux2_1 _21470_ (.A0(_01857_),
    .A1(net525),
    .S(net6646),
    .X(_07875_));
 sg13g2_nand2_1 _21471_ (.Y(_07876_),
    .A(_00368_),
    .B(net6928));
 sg13g2_o21ai_1 _21472_ (.B1(net6924),
    .Y(_07877_),
    .A1(_00266_),
    .A2(net7048));
 sg13g2_nand2_1 _21473_ (.Y(_07878_),
    .A(_07876_),
    .B(_07877_));
 sg13g2_a221oi_1 _21474_ (.B2(_00523_),
    .C1(_07878_),
    .B1(net6882),
    .A1(net6577),
    .Y(_07879_),
    .A2(net6883));
 sg13g2_o21ai_1 _21475_ (.B1(net6765),
    .Y(_07880_),
    .A1(net306),
    .A2(net6920));
 sg13g2_nor2b_1 _21476_ (.A(net7675),
    .B_N(net7676),
    .Y(_07881_));
 sg13g2_nor2_1 _21477_ (.A(_07879_),
    .B(_07880_),
    .Y(_07882_));
 sg13g2_a21o_1 _21478_ (.A2(net6773),
    .A1(_01691_),
    .B1(_07882_),
    .X(_07883_));
 sg13g2_mux2_1 _21479_ (.A0(_01856_),
    .A1(_07883_),
    .S(net7453),
    .X(net524));
 sg13g2_nand2b_1 _21480_ (.Y(_07884_),
    .B(net7676),
    .A_N(net7675));
 sg13g2_mux2_1 _21481_ (.A0(_01856_),
    .A1(net524),
    .S(net6647),
    .X(_07885_));
 sg13g2_o21ai_1 _21482_ (.B1(_07676_),
    .Y(_07886_),
    .A1(_00522_),
    .A2(_07678_));
 sg13g2_inv_1 _21483_ (.Y(_07887_),
    .A(_07888_));
 sg13g2_o21ai_1 _21484_ (.B1(net6924),
    .Y(_07888_),
    .A1(_00265_),
    .A2(net7048));
 sg13g2_a221oi_1 _21485_ (.B2(_00367_),
    .C1(_07887_),
    .B1(net6926),
    .A1(net455),
    .Y(_07889_),
    .A2(net6883));
 sg13g2_nor3_1 _21486_ (.A(_07780_),
    .B(_07872_),
    .C(_07884_),
    .Y(_07890_));
 sg13g2_o21ai_1 _21487_ (.B1(net6765),
    .Y(_07891_),
    .A1(net305),
    .A2(net6920));
 sg13g2_a21oi_1 _21488_ (.A1(_07886_),
    .A2(_07889_),
    .Y(_07892_),
    .B1(_07891_));
 sg13g2_a21o_1 _21489_ (.A2(net6773),
    .A1(_01690_),
    .B1(_07892_),
    .X(_07893_));
 sg13g2_mux2_1 _21490_ (.A0(_01855_),
    .A1(_07893_),
    .S(net7452),
    .X(net523));
 sg13g2_mux2_1 _21491_ (.A0(_01855_),
    .A1(net523),
    .S(net6646),
    .X(_07894_));
 sg13g2_nand4_1 _21492_ (.B(_07783_),
    .C(_07870_),
    .A(net7679),
    .Y(_07895_),
    .D(_07881_));
 sg13g2_nand2_1 _21493_ (.Y(_07896_),
    .A(_00366_),
    .B(net6928));
 sg13g2_and2_1 _21494_ (.A(net7610),
    .B(_07895_),
    .X(_07897_));
 sg13g2_o21ai_1 _21495_ (.B1(net6925),
    .Y(_07898_),
    .A1(_00264_),
    .A2(net7049));
 sg13g2_nand2_1 _21496_ (.Y(_07899_),
    .A(_07896_),
    .B(_07898_));
 sg13g2_a221oi_1 _21497_ (.B2(_00521_),
    .C1(_07899_),
    .B1(net6882),
    .A1(net454),
    .Y(_07900_),
    .A2(net6883));
 sg13g2_o21ai_1 _21498_ (.B1(net6766),
    .Y(_07901_),
    .A1(net304),
    .A2(net6921));
 sg13g2_or2_1 _21499_ (.X(_07902_),
    .B(_07901_),
    .A(_07900_));
 sg13g2_o21ai_1 _21500_ (.B1(_07902_),
    .Y(_07903_),
    .A1(_15560_),
    .A2(net6767));
 sg13g2_mux2_1 _21501_ (.A0(_01854_),
    .A1(_07903_),
    .S(net7452),
    .X(net522));
 sg13g2_nand2b_1 _21502_ (.Y(_07904_),
    .B(_01911_),
    .A_N(net7679));
 sg13g2_mux2_1 _21503_ (.A0(_01854_),
    .A1(net522),
    .S(net6646),
    .X(_07905_));
 sg13g2_nand2_1 _21504_ (.Y(_07906_),
    .A(_00365_),
    .B(net6928));
 sg13g2_o21ai_1 _21505_ (.B1(net6925),
    .Y(_07907_),
    .A1(_00263_),
    .A2(net7049));
 sg13g2_nand2_1 _21506_ (.Y(_07908_),
    .A(_07906_),
    .B(_07907_));
 sg13g2_a221oi_1 _21507_ (.B2(_00520_),
    .C1(_07908_),
    .B1(net6882),
    .A1(net6604),
    .Y(_07909_),
    .A2(net6883));
 sg13g2_and2_1 _21508_ (.A(_01911_),
    .B(net7679),
    .X(_07910_));
 sg13g2_o21ai_1 _21509_ (.B1(net6765),
    .Y(_07911_),
    .A1(net303),
    .A2(net6920));
 sg13g2_nor2_1 _21510_ (.A(_07909_),
    .B(_07911_),
    .Y(_07912_));
 sg13g2_a21o_1 _21511_ (.A2(net6773),
    .A1(_01688_),
    .B1(_07912_),
    .X(_07913_));
 sg13g2_mux2_1 _21512_ (.A0(_01853_),
    .A1(_07913_),
    .S(net7453),
    .X(net521));
 sg13g2_mux2_1 _21513_ (.A0(_01853_),
    .A1(net521),
    .S(net6647),
    .X(_07914_));
 sg13g2_nand2_1 _21514_ (.Y(_07915_),
    .A(_00364_),
    .B(net6928));
 sg13g2_o21ai_1 _21515_ (.B1(net6925),
    .Y(_07916_),
    .A1(_00262_),
    .A2(net7049));
 sg13g2_nand2_1 _21516_ (.Y(_07917_),
    .A(_07915_),
    .B(_07916_));
 sg13g2_a22oi_1 _21517_ (.Y(_07918_),
    .B1(_07910_),
    .B2(_07870_),
    .A2(_07904_),
    .A1(_07587_));
 sg13g2_a221oi_1 _21518_ (.B2(_00519_),
    .C1(_07917_),
    .B1(net6882),
    .A1(net6606),
    .Y(_07919_),
    .A2(_07671_));
 sg13g2_o21ai_1 _21519_ (.B1(net6766),
    .Y(_07920_),
    .A1(net302),
    .A2(net6921));
 sg13g2_nor2_1 _21520_ (.A(_07919_),
    .B(_07920_),
    .Y(_07921_));
 sg13g2_a21o_1 _21521_ (.A2(net6773),
    .A1(_01687_),
    .B1(_07921_),
    .X(_07922_));
 sg13g2_mux2_1 _21522_ (.A0(_01852_),
    .A1(_07922_),
    .S(net7453),
    .X(net520));
 sg13g2_mux2_1 _21523_ (.A0(_01852_),
    .A1(net520),
    .S(net6647),
    .X(_07923_));
 sg13g2_nand2_1 _21524_ (.Y(_07924_),
    .A(_00363_),
    .B(net6928));
 sg13g2_nor2b_1 _21525_ (.A(_01912_),
    .B_N(_01908_),
    .Y(_07925_));
 sg13g2_o21ai_1 _21526_ (.B1(_07690_),
    .Y(_07926_),
    .A1(_00261_),
    .A2(net7049));
 sg13g2_nand2_1 _21527_ (.Y(_07927_),
    .A(_07924_),
    .B(_07926_));
 sg13g2_a221oi_1 _21528_ (.B2(_00518_),
    .C1(_07927_),
    .B1(net6882),
    .A1(net6584),
    .Y(_07928_),
    .A2(_07671_));
 sg13g2_o21ai_1 _21529_ (.B1(net6764),
    .Y(_07929_),
    .A1(net301),
    .A2(net6922));
 sg13g2_nor2_1 _21530_ (.A(net7676),
    .B(_07925_),
    .Y(_07930_));
 sg13g2_nor2_1 _21531_ (.A(_07928_),
    .B(_07929_),
    .Y(_07931_));
 sg13g2_a21o_1 _21532_ (.A2(net6772),
    .A1(_01686_),
    .B1(_07931_),
    .X(_07932_));
 sg13g2_mux2_1 _21533_ (.A0(_01851_),
    .A1(_07932_),
    .S(net7453),
    .X(net519));
 sg13g2_mux2_1 _21534_ (.A0(_01851_),
    .A1(net519),
    .S(net6647),
    .X(_07933_));
 sg13g2_o21ai_1 _21535_ (.B1(_07676_),
    .Y(_07934_),
    .A1(_00517_),
    .A2(_07678_));
 sg13g2_or3_1 _21536_ (.A(_01914_),
    .B(net7676),
    .C(_07925_),
    .X(_07935_));
 sg13g2_inv_1 _21537_ (.Y(_07936_),
    .A(_07937_));
 sg13g2_o21ai_1 _21538_ (.B1(_07690_),
    .Y(_07937_),
    .A1(_00260_),
    .A2(net7049));
 sg13g2_a221oi_1 _21539_ (.B2(_00362_),
    .C1(_07936_),
    .B1(net6928),
    .A1(net450),
    .Y(_07938_),
    .A2(net6883));
 sg13g2_o21ai_1 _21540_ (.B1(net6765),
    .Y(_07939_),
    .A1(net300),
    .A2(net6920));
 sg13g2_o21ai_1 _21541_ (.B1(_07935_),
    .Y(_07940_),
    .A1(net7675),
    .A2(_07918_));
 sg13g2_a21oi_1 _21542_ (.A1(_07934_),
    .A2(_07938_),
    .Y(_07941_),
    .B1(_07939_));
 sg13g2_a21o_1 _21543_ (.A2(net6772),
    .A1(_01685_),
    .B1(_07941_),
    .X(_07942_));
 sg13g2_mux2_1 _21544_ (.A0(_01850_),
    .A1(_07942_),
    .S(net7453),
    .X(net518));
 sg13g2_mux2_1 _21545_ (.A0(_01850_),
    .A1(net518),
    .S(net6647),
    .X(_07943_));
 sg13g2_nand2_1 _21546_ (.Y(_07944_),
    .A(_00360_),
    .B(net6928));
 sg13g2_o21ai_1 _21547_ (.B1(net6924),
    .Y(_07945_),
    .A1(_00258_),
    .A2(net7048));
 sg13g2_nor2_1 _21548_ (.A(net7679),
    .B(_07562_),
    .Y(_07946_));
 sg13g2_nand2_1 _21549_ (.Y(_07947_),
    .A(_07944_),
    .B(_07945_));
 sg13g2_nand3b_1 _21550_ (.B(_01897_),
    .C(_01886_),
    .Y(_07948_),
    .A_N(_01908_));
 sg13g2_a221oi_1 _21551_ (.B2(_00516_),
    .C1(_07947_),
    .B1(net6882),
    .A1(net6607),
    .Y(_07949_),
    .A2(net6883));
 sg13g2_o21ai_1 _21552_ (.B1(net6765),
    .Y(_07950_),
    .A1(net299),
    .A2(net6920));
 sg13g2_nor2_1 _21553_ (.A(_07949_),
    .B(_07950_),
    .Y(_07951_));
 sg13g2_inv_1 _21554_ (.Y(_07952_),
    .A(_07953_));
 sg13g2_a21o_1 _21555_ (.A2(net6772),
    .A1(_01684_),
    .B1(_07951_),
    .X(_07953_));
 sg13g2_mux2_1 _21556_ (.A0(_01849_),
    .A1(_07953_),
    .S(net7454),
    .X(net517));
 sg13g2_nand2b_1 _21557_ (.Y(_07954_),
    .B(_01912_),
    .A_N(_01911_));
 sg13g2_mux2_1 _21558_ (.A0(_01849_),
    .A1(net517),
    .S(net6647),
    .X(_07955_));
 sg13g2_nor2_1 _21559_ (.A(net7451),
    .B(_01848_),
    .Y(_07956_));
 sg13g2_nand2_1 _21560_ (.Y(_07957_),
    .A(_00359_),
    .B(net6926));
 sg13g2_o21ai_1 _21561_ (.B1(net6923),
    .Y(_07958_),
    .A1(_00257_),
    .A2(net7047));
 sg13g2_nand2_1 _21562_ (.Y(_07959_),
    .A(_07957_),
    .B(_07958_));
 sg13g2_a221oi_1 _21563_ (.B2(_00515_),
    .C1(_07959_),
    .B1(net6881),
    .A1(net6608),
    .Y(_07960_),
    .A2(net6884));
 sg13g2_o21ai_1 _21564_ (.B1(net6764),
    .Y(_07961_),
    .A1(net298),
    .A2(net6921));
 sg13g2_nor2_1 _21565_ (.A(_07960_),
    .B(_07961_),
    .Y(_07962_));
 sg13g2_a21oi_1 _21566_ (.A1(_01683_),
    .A2(net6772),
    .Y(_07963_),
    .B1(_07962_));
 sg13g2_a21oi_1 _21567_ (.A1(net7451),
    .A2(_07963_),
    .Y(net516),
    .B1(_07956_));
 sg13g2_nor2_1 _21568_ (.A(_07872_),
    .B(_07954_),
    .Y(_07964_));
 sg13g2_mux2_1 _21569_ (.A0(_01848_),
    .A1(net516),
    .S(net6645),
    .X(_07965_));
 sg13g2_nor2_1 _21570_ (.A(net7451),
    .B(_01847_),
    .Y(_07966_));
 sg13g2_nand2_1 _21571_ (.Y(_07967_),
    .A(_00358_),
    .B(net6926));
 sg13g2_o21ai_1 _21572_ (.B1(net6923),
    .Y(_07968_),
    .A1(_00256_),
    .A2(net7047));
 sg13g2_nand2_1 _21573_ (.Y(_07969_),
    .A(_07967_),
    .B(_07968_));
 sg13g2_nor3_1 _21574_ (.A(_07872_),
    .B(_07948_),
    .C(_07954_),
    .Y(_07970_));
 sg13g2_a221oi_1 _21575_ (.B2(_00514_),
    .C1(_07969_),
    .B1(net6881),
    .A1(net6609),
    .Y(_07971_),
    .A2(net6884));
 sg13g2_o21ai_1 _21576_ (.B1(net6765),
    .Y(_07972_),
    .A1(net297),
    .A2(net6920));
 sg13g2_inv_1 _21577_ (.Y(_07973_),
    .A(_07970_));
 sg13g2_nor2_1 _21578_ (.A(_07971_),
    .B(_07972_),
    .Y(_07974_));
 sg13g2_a21oi_1 _21579_ (.A1(_01682_),
    .A2(net6772),
    .Y(_07975_),
    .B1(_07974_));
 sg13g2_a21oi_1 _21580_ (.A1(net7451),
    .A2(_07975_),
    .Y(net515),
    .B1(_07966_));
 sg13g2_mux2_1 _21581_ (.A0(_01847_),
    .A1(net515),
    .S(net6645),
    .X(_07976_));
 sg13g2_nor2_1 _21582_ (.A(net7451),
    .B(_01846_),
    .Y(_07977_));
 sg13g2_or4_1 _21583_ (.A(_01910_),
    .B(_01907_),
    .C(net7681),
    .D(net7682),
    .X(_07978_));
 sg13g2_o21ai_1 _21584_ (.B1(_07676_),
    .Y(_07979_),
    .A1(_00513_),
    .A2(_07678_));
 sg13g2_nand2_1 _21585_ (.Y(_07980_),
    .A(_00357_),
    .B(net6926));
 sg13g2_o21ai_1 _21586_ (.B1(net6923),
    .Y(_07981_),
    .A1(_00255_),
    .A2(net7047));
 sg13g2_nand3b_1 _21587_ (.B(net7931),
    .C(net7921),
    .Y(_07982_),
    .A_N(net7928));
 sg13g2_nand3_1 _21588_ (.B(_07980_),
    .C(_07981_),
    .A(_07979_),
    .Y(_07983_));
 sg13g2_a21oi_1 _21589_ (.A1(net446),
    .A2(net6885),
    .Y(_07984_),
    .B1(_07983_));
 sg13g2_o21ai_1 _21590_ (.B1(net6763),
    .Y(_07985_),
    .A1(net296),
    .A2(net6922));
 sg13g2_nor2_1 _21591_ (.A(_07984_),
    .B(_07985_),
    .Y(_07986_));
 sg13g2_a21oi_1 _21592_ (.A1(_01681_),
    .A2(net6775),
    .Y(_07987_),
    .B1(_07986_));
 sg13g2_inv_1 _21593_ (.Y(_07988_),
    .A(_07987_));
 sg13g2_a21oi_1 _21594_ (.A1(net7451),
    .A2(_07987_),
    .Y(net514),
    .B1(_07977_));
 sg13g2_mux2_1 _21595_ (.A0(_01846_),
    .A1(net514),
    .S(net6645),
    .X(_07989_));
 sg13g2_nand2_1 _21596_ (.Y(_07990_),
    .A(_00356_),
    .B(net6929));
 sg13g2_o21ai_1 _21597_ (.B1(_07690_),
    .Y(_07991_),
    .A1(_00254_),
    .A2(net7049));
 sg13g2_nand2_1 _21598_ (.Y(_07992_),
    .A(_07990_),
    .B(_07991_));
 sg13g2_nor2b_1 _21599_ (.A(_07982_),
    .B_N(_07978_),
    .Y(_07993_));
 sg13g2_a221oi_1 _21600_ (.B2(_00512_),
    .C1(_07992_),
    .B1(net6882),
    .A1(net445),
    .Y(_07994_),
    .A2(_07671_));
 sg13g2_o21ai_1 _21601_ (.B1(net6768),
    .Y(_07995_),
    .A1(net295),
    .A2(_07704_));
 sg13g2_or2_1 _21602_ (.X(_07996_),
    .B(_07995_),
    .A(_07994_));
 sg13g2_o21ai_1 _21603_ (.B1(_07996_),
    .Y(_07997_),
    .A1(_02013_),
    .A2(net6761));
 sg13g2_mux2_1 _21604_ (.A0(_01845_),
    .A1(_07997_),
    .S(net7451),
    .X(net513));
 sg13g2_mux2_1 _21605_ (.A0(_01845_),
    .A1(net513),
    .S(net6645),
    .X(_07998_));
 sg13g2_nor2_1 _21606_ (.A(_00253_),
    .B(_07661_),
    .Y(_07999_));
 sg13g2_o21ai_1 _21607_ (.B1(_07697_),
    .Y(_08000_),
    .A1(_07684_),
    .A2(_07999_));
 sg13g2_a221oi_1 _21608_ (.B2(net7626),
    .C1(_07662_),
    .B1(_08000_),
    .A1(_00355_),
    .Y(_08001_),
    .A2(net6927));
 sg13g2_inv_1 _21609_ (.Y(_08002_),
    .A(_08001_));
 sg13g2_o21ai_1 _21610_ (.B1(_07970_),
    .Y(_08003_),
    .A1(_07841_),
    .A2(_07993_));
 sg13g2_a221oi_1 _21611_ (.B2(_00511_),
    .C1(_08002_),
    .B1(_07679_),
    .A1(net444),
    .Y(_08004_),
    .A2(net6885));
 sg13g2_o21ai_1 _21612_ (.B1(net6763),
    .Y(_08005_),
    .A1(net294),
    .A2(_07704_));
 sg13g2_or2_1 _21613_ (.X(_08006_),
    .B(_08005_),
    .A(_08004_));
 sg13g2_o21ai_1 _21614_ (.B1(_08006_),
    .Y(_08007_),
    .A1(_02016_),
    .A2(net6761));
 sg13g2_nand3_1 _21615_ (.B(_07940_),
    .C(_08003_),
    .A(_07897_),
    .Y(_08008_));
 sg13g2_mux2_1 _21616_ (.A0(_01844_),
    .A1(_08007_),
    .S(net7451),
    .X(net512));
 sg13g2_mux2_1 _21617_ (.A0(_01844_),
    .A1(net512),
    .S(net6645),
    .X(_08009_));
 sg13g2_a21oi_1 _21618_ (.A1(_07616_),
    .A2(_07864_),
    .Y(_08010_),
    .B1(_08008_));
 sg13g2_nand2_1 _21619_ (.Y(_08011_),
    .A(_00510_),
    .B(net6881));
 sg13g2_a21o_1 _21620_ (.A2(_07864_),
    .A1(_07616_),
    .B1(_08008_),
    .X(_08012_));
 sg13g2_nor3_1 _21621_ (.A(_07662_),
    .B(_07683_),
    .C(_07688_),
    .Y(_08013_));
 sg13g2_nor2_1 _21622_ (.A(net7438),
    .B(_08012_),
    .Y(_08014_));
 sg13g2_nand2_1 _21623_ (.Y(_08015_),
    .A(net7105),
    .B(_07660_));
 sg13g2_nand2_1 _21624_ (.Y(_08016_),
    .A(_07605_),
    .B(_08010_));
 sg13g2_o21ai_1 _21625_ (.B1(net7626),
    .Y(_08017_),
    .A1(_00252_),
    .A2(_08015_));
 sg13g2_a21oi_1 _21626_ (.A1(net7986),
    .A2(_08017_),
    .Y(_08018_),
    .B1(_08013_));
 sg13g2_nor2_1 _21627_ (.A(net7674),
    .B(_07993_),
    .Y(_08019_));
 sg13g2_a221oi_1 _21628_ (.B2(_00354_),
    .C1(_08018_),
    .B1(net6927),
    .A1(net6600),
    .Y(_08020_),
    .A2(net6884));
 sg13g2_o21ai_1 _21629_ (.B1(net6764),
    .Y(_08021_),
    .A1(net293),
    .A2(net6922));
 sg13g2_a21oi_1 _21630_ (.A1(_08011_),
    .A2(_08020_),
    .Y(_08022_),
    .B1(_08021_));
 sg13g2_a21o_1 _21631_ (.A2(net6774),
    .A1(_01678_),
    .B1(_08022_),
    .X(_08023_));
 sg13g2_mux2_1 _21632_ (.A0(_01843_),
    .A1(_08023_),
    .S(net7455),
    .X(net511));
 sg13g2_mux2_1 _21633_ (.A0(_01843_),
    .A1(net511),
    .S(net6645),
    .X(_08024_));
 sg13g2_nand2_1 _21634_ (.Y(_08025_),
    .A(_00509_),
    .B(net6881));
 sg13g2_nor2_1 _21635_ (.A(net7921),
    .B(_07701_),
    .Y(_08026_));
 sg13g2_o21ai_1 _21636_ (.B1(net7626),
    .Y(_08027_),
    .A1(_00251_),
    .A2(_08015_));
 sg13g2_nand2_1 _21637_ (.Y(_08028_),
    .A(net7930),
    .B(_07780_));
 sg13g2_a21oi_1 _21638_ (.A1(net7986),
    .A2(_08027_),
    .Y(_08029_),
    .B1(_08013_));
 sg13g2_a221oi_1 _21639_ (.B2(_00353_),
    .C1(_08029_),
    .B1(net6927),
    .A1(net442),
    .Y(_08030_),
    .A2(net6885));
 sg13g2_o21ai_1 _21640_ (.B1(net6764),
    .Y(_08031_),
    .A1(net292),
    .A2(net6922));
 sg13g2_o21ai_1 _21641_ (.B1(_08028_),
    .Y(_08032_),
    .A1(_09244_),
    .A2(net7930));
 sg13g2_a21oi_1 _21642_ (.A1(_08025_),
    .A2(_08030_),
    .Y(_08033_),
    .B1(_08031_));
 sg13g2_a21o_1 _21643_ (.A2(net6774),
    .A1(_01677_),
    .B1(_08033_),
    .X(_08034_));
 sg13g2_mux2_1 _21644_ (.A0(_01842_),
    .A1(_08034_),
    .S(net7455),
    .X(net510));
 sg13g2_mux2_1 _21645_ (.A0(_01842_),
    .A1(net510),
    .S(net6645),
    .X(_08035_));
 sg13g2_nor2_1 _21646_ (.A(net291),
    .B(net6921),
    .Y(_08036_));
 sg13g2_o21ai_1 _21647_ (.B1(_07676_),
    .Y(_08037_),
    .A1(_00508_),
    .A2(_07678_));
 sg13g2_o21ai_1 _21648_ (.B1(net6924),
    .Y(_08038_),
    .A1(_00250_),
    .A2(net7048));
 sg13g2_inv_1 _21649_ (.Y(_08039_),
    .A(_08038_));
 sg13g2_a221oi_1 _21650_ (.B2(_00352_),
    .C1(_08039_),
    .B1(net6927),
    .A1(net6621),
    .Y(_08040_),
    .A2(net6883));
 sg13g2_a21oi_1 _21651_ (.A1(_08037_),
    .A2(_08040_),
    .Y(_08041_),
    .B1(_08036_));
 sg13g2_inv_1 _21652_ (.Y(_08042_),
    .A(_08041_));
 sg13g2_nand2_1 _21653_ (.Y(_08043_),
    .A(net6760),
    .B(_08041_));
 sg13g2_o21ai_1 _21654_ (.B1(_08043_),
    .Y(_08044_),
    .A1(_02025_),
    .A2(net6760));
 sg13g2_mux2_1 _21655_ (.A0(_01841_),
    .A1(_08044_),
    .S(net7452),
    .X(net509));
 sg13g2_mux2_1 _21656_ (.A0(_01841_),
    .A1(net509),
    .S(net6646),
    .X(_08045_));
 sg13g2_nor2_1 _21657_ (.A(net290),
    .B(_07704_),
    .Y(_08046_));
 sg13g2_a221oi_1 _21658_ (.B2(_08032_),
    .C1(_08563_),
    .B1(_07834_),
    .A1(_07806_),
    .Y(_08047_),
    .A2(_07826_));
 sg13g2_o21ai_1 _21659_ (.B1(net7626),
    .Y(_08048_),
    .A1(_00249_),
    .A2(_08015_));
 sg13g2_a21oi_1 _21660_ (.A1(net7986),
    .A2(_08048_),
    .Y(_08049_),
    .B1(_08013_));
 sg13g2_a21o_1 _21661_ (.A2(net6927),
    .A1(_00351_),
    .B1(_08049_),
    .X(_08050_));
 sg13g2_a221oi_1 _21662_ (.B2(_00507_),
    .C1(_08050_),
    .B1(_07679_),
    .A1(net440),
    .Y(_08051_),
    .A2(net6885));
 sg13g2_or3_1 _21663_ (.A(net6773),
    .B(_08046_),
    .C(_08051_),
    .X(_08052_));
 sg13g2_o21ai_1 _21664_ (.B1(_08052_),
    .Y(_08053_),
    .A1(_02029_),
    .A2(net6760));
 sg13g2_mux2_1 _21665_ (.A0(_01840_),
    .A1(_08053_),
    .S(net7452),
    .X(net508));
 sg13g2_mux2_1 _21666_ (.A0(_01840_),
    .A1(net508),
    .S(net6646),
    .X(_08054_));
 sg13g2_and2_1 _21667_ (.A(net384),
    .B(net538),
    .X(_08055_));
 sg13g2_a21oi_1 _21668_ (.A1(net7937),
    .A2(_08055_),
    .Y(_08056_),
    .B1(_01839_));
 sg13g2_a21oi_1 _21669_ (.A1(net417),
    .A2(net7937),
    .Y(_08057_),
    .B1(_08056_));
 sg13g2_nand2b_1 _21670_ (.Y(_08058_),
    .B(net417),
    .A_N(_01839_));
 sg13g2_a21oi_1 _21671_ (.A1(net7937),
    .A2(_08058_),
    .Y(_08059_),
    .B1(_08055_));
 sg13g2_inv_1 _21672_ (.Y(_08060_),
    .A(_08059_));
 sg13g2_a21oi_1 _21673_ (.A1(net385),
    .A2(net396),
    .Y(_08061_),
    .B1(net383));
 sg13g2_a21oi_1 _21674_ (.A1(_01750_),
    .A2(_01739_),
    .Y(_08062_),
    .B1(_01705_));
 sg13g2_mux2_1 _21675_ (.A0(_08061_),
    .A1(_08062_),
    .S(_01835_),
    .X(_08063_));
 sg13g2_inv_1 _21676_ (.Y(_08064_),
    .A(_08065_));
 sg13g2_nand2_1 _21677_ (.Y(_08065_),
    .A(_15152_),
    .B(_08063_));
 sg13g2_nor2_1 _21678_ (.A(_07045_),
    .B(_08064_),
    .Y(_08066_));
 sg13g2_nand2_2 _21679_ (.Y(_08067_),
    .A(_08065_),
    .B(_07044_));
 sg13g2_nand2_1 _21680_ (.Y(_08068_),
    .A(net7956),
    .B(_07007_));
 sg13g2_a21oi_1 _21681_ (.A1(_01836_),
    .A2(_07007_),
    .Y(_08069_),
    .B1(_01837_));
 sg13g2_nor3_1 _21682_ (.A(net6761),
    .B(_08066_),
    .C(_08069_),
    .Y(_08070_));
 sg13g2_nor3_1 _21683_ (.A(_07614_),
    .B(_08019_),
    .C(_08047_),
    .Y(_08071_));
 sg13g2_a21o_1 _21684_ (.A2(_08067_),
    .A1(_07008_),
    .B1(net6761),
    .X(_08072_));
 sg13g2_a21oi_1 _21685_ (.A1(_08066_),
    .A2(_08069_),
    .Y(_08073_),
    .B1(_08072_));
 sg13g2_mux2_1 _21686_ (.A0(_07008_),
    .A1(_07014_),
    .S(_08067_),
    .X(_08074_));
 sg13g2_nor2_1 _21687_ (.A(net6761),
    .B(_08074_),
    .Y(_08075_));
 sg13g2_nand3b_1 _21688_ (.B(_07007_),
    .C(_08067_),
    .Y(_08076_),
    .A_N(_01835_));
 sg13g2_o21ai_1 _21689_ (.B1(_08076_),
    .Y(_08077_),
    .A1(_08067_),
    .A2(_07008_));
 sg13g2_a22oi_1 _21690_ (.Y(_08078_),
    .B1(_07970_),
    .B2(net7920),
    .A2(_07602_),
    .A1(_09282_));
 sg13g2_nor2_1 _21691_ (.A(_01834_),
    .B(net5812),
    .Y(_08079_));
 sg13g2_a21oi_1 _21692_ (.A1(net5812),
    .A2(_07359_),
    .Y(_08080_),
    .B1(_08079_));
 sg13g2_nor2_1 _21693_ (.A(_01837_),
    .B(_08068_),
    .Y(_08081_));
 sg13g2_mux2_1 _21694_ (.A0(_01833_),
    .A1(net409),
    .S(net7298),
    .X(_08082_));
 sg13g2_mux2_1 _21695_ (.A0(_01832_),
    .A1(net408),
    .S(net7297),
    .X(_08083_));
 sg13g2_mux2_1 _21696_ (.A0(_01831_),
    .A1(net406),
    .S(net7297),
    .X(_08084_));
 sg13g2_mux2_1 _21697_ (.A0(_01830_),
    .A1(net405),
    .S(net7297),
    .X(_08085_));
 sg13g2_mux2_1 _21698_ (.A0(_01829_),
    .A1(net404),
    .S(net7298),
    .X(_08086_));
 sg13g2_mux2_1 _21699_ (.A0(_01828_),
    .A1(net403),
    .S(net7298),
    .X(_08087_));
 sg13g2_mux2_1 _21700_ (.A0(_01827_),
    .A1(_07370_),
    .S(net5818),
    .X(_08088_));
 sg13g2_mux2_1 _21701_ (.A0(_01826_),
    .A1(net402),
    .S(net7297),
    .X(_08089_));
 sg13g2_a21oi_1 _21702_ (.A1(net7928),
    .A2(_07602_),
    .Y(_08090_),
    .B1(_09324_));
 sg13g2_mux2_1 _21703_ (.A0(_01825_),
    .A1(net401),
    .S(net7300),
    .X(_08091_));
 sg13g2_mux2_1 _21704_ (.A0(_01824_),
    .A1(net400),
    .S(net7300),
    .X(_08092_));
 sg13g2_mux2_1 _21705_ (.A0(_01823_),
    .A1(net399),
    .S(net7300),
    .X(_08093_));
 sg13g2_mux2_1 _21706_ (.A0(_01822_),
    .A1(net398),
    .S(net7300),
    .X(_08094_));
 sg13g2_mux2_1 _21707_ (.A0(_01821_),
    .A1(net397),
    .S(net7298),
    .X(_08095_));
 sg13g2_mux2_1 _21708_ (.A0(_01820_),
    .A1(net395),
    .S(net7297),
    .X(_08096_));
 sg13g2_mux2_1 _21709_ (.A0(_01819_),
    .A1(net394),
    .S(_08081_),
    .X(_08097_));
 sg13g2_mux2_1 _21710_ (.A0(_01818_),
    .A1(net393),
    .S(net7299),
    .X(_08098_));
 sg13g2_mux2_1 _21711_ (.A0(_01817_),
    .A1(net392),
    .S(net7299),
    .X(_08099_));
 sg13g2_a21o_1 _21712_ (.A2(_08078_),
    .A1(_09324_),
    .B1(_08090_),
    .X(_08100_));
 sg13g2_mux2_1 _21713_ (.A0(_01816_),
    .A1(_07388_),
    .S(net5818),
    .X(_08101_));
 sg13g2_a22oi_1 _21714_ (.Y(_08102_),
    .B1(_07970_),
    .B2(net7929),
    .A2(_07602_),
    .A1(net7928));
 sg13g2_mux2_1 _21715_ (.A0(_01815_),
    .A1(net391),
    .S(net7298),
    .X(_08103_));
 sg13g2_mux2_1 _21716_ (.A0(_01814_),
    .A1(net390),
    .S(net7297),
    .X(_08104_));
 sg13g2_mux2_1 _21717_ (.A0(_01813_),
    .A1(net389),
    .S(net7299),
    .X(_08105_));
 sg13g2_mux2_1 _21718_ (.A0(_01812_),
    .A1(net388),
    .S(net7297),
    .X(_08106_));
 sg13g2_mux2_1 _21719_ (.A0(_01811_),
    .A1(net387),
    .S(net7298),
    .X(_08107_));
 sg13g2_or2_1 _21720_ (.X(_08108_),
    .B(_08102_),
    .A(net7920));
 sg13g2_mux2_1 _21721_ (.A0(_01810_),
    .A1(net386),
    .S(net7298),
    .X(_08109_));
 sg13g2_mux2_1 _21722_ (.A0(_01809_),
    .A1(net416),
    .S(net7299),
    .X(_08110_));
 sg13g2_mux2_1 _21723_ (.A0(_01808_),
    .A1(net415),
    .S(net7300),
    .X(_08111_));
 sg13g2_mux2_1 _21724_ (.A0(_01807_),
    .A1(net414),
    .S(net7300),
    .X(_08112_));
 sg13g2_mux2_1 _21725_ (.A0(_01806_),
    .A1(net413),
    .S(net7300),
    .X(_08113_));
 sg13g2_mux2_1 _21726_ (.A0(_01805_),
    .A1(_07403_),
    .S(net5818),
    .X(_08114_));
 sg13g2_mux2_1 _21727_ (.A0(_01804_),
    .A1(net412),
    .S(net7300),
    .X(_08115_));
 sg13g2_mux2_1 _21728_ (.A0(_01803_),
    .A1(net411),
    .S(net7298),
    .X(_08116_));
 sg13g2_mux2_1 _21729_ (.A0(_01802_),
    .A1(net410),
    .S(net7299),
    .X(_08117_));
 sg13g2_mux2_1 _21730_ (.A0(_01801_),
    .A1(net407),
    .S(_08081_),
    .X(_08118_));
 sg13g2_mux2_1 _21731_ (.A0(_01800_),
    .A1(net396),
    .S(net7299),
    .X(_08119_));
 sg13g2_mux2_1 _21732_ (.A0(_01799_),
    .A1(net385),
    .S(_08081_),
    .X(_08120_));
 sg13g2_nand2_1 _21733_ (.Y(_08121_),
    .A(_07007_),
    .B(_07628_));
 sg13g2_mux2_2 _21734_ (.A0(_08069_),
    .A1(_08121_),
    .S(_08067_),
    .X(_08122_));
 sg13g2_nor2b_1 _21735_ (.A(net7947),
    .B_N(net409),
    .Y(_08123_));
 sg13g2_a21oi_1 _21736_ (.A1(net7944),
    .A2(_01833_),
    .Y(_08124_),
    .B1(_08123_));
 sg13g2_nand4_1 _21737_ (.B(_07940_),
    .C(_08100_),
    .A(_07897_),
    .Y(_08125_),
    .D(_08108_));
 sg13g2_nor2_1 _21738_ (.A(_08071_),
    .B(_08125_),
    .Y(_08126_));
 sg13g2_nand2_2 _21739_ (.Y(_08127_),
    .A(net5874),
    .B(_01798_));
 sg13g2_o21ai_1 _21740_ (.B1(_08127_),
    .Y(_08128_),
    .A1(net5875),
    .A2(_08124_));
 sg13g2_nor2b_1 _21741_ (.A(net7940),
    .B_N(net408),
    .Y(_08129_));
 sg13g2_a21oi_1 _21742_ (.A1(net7940),
    .A2(_01832_),
    .Y(_08130_),
    .B1(_08129_));
 sg13g2_nand2_1 _21743_ (.Y(_08131_),
    .A(net7438),
    .B(_07757_));
 sg13g2_nand2_2 _21744_ (.Y(_08132_),
    .A(net5871),
    .B(_01797_));
 sg13g2_nand4_1 _21745_ (.B(net7920),
    .C(_07635_),
    .A(_08711_),
    .Y(_08133_),
    .D(_07644_));
 sg13g2_o21ai_1 _21746_ (.B1(_08132_),
    .Y(_08134_),
    .A1(net5871),
    .A2(_08130_));
 sg13g2_nor2b_1 _21747_ (.A(net7941),
    .B_N(net406),
    .Y(_08135_));
 sg13g2_a21oi_1 _21748_ (.A1(net7941),
    .A2(_01831_),
    .Y(_08136_),
    .B1(_08135_));
 sg13g2_nand2_2 _21749_ (.Y(_08137_),
    .A(net5870),
    .B(_01796_));
 sg13g2_nand4_1 _21750_ (.B(net7610),
    .C(net7609),
    .A(net7929),
    .Y(_08138_),
    .D(_07608_));
 sg13g2_o21ai_1 _21751_ (.B1(_08137_),
    .Y(_08139_),
    .A1(net5870),
    .A2(_08136_));
 sg13g2_a21oi_1 _21752_ (.A1(net7674),
    .A2(_08133_),
    .Y(_08140_),
    .B1(_08138_));
 sg13g2_nor2b_1 _21753_ (.A(net7939),
    .B_N(net405),
    .Y(_08141_));
 sg13g2_a21oi_1 _21754_ (.A1(net7940),
    .A2(_01830_),
    .Y(_08142_),
    .B1(_08141_));
 sg13g2_nand2_2 _21755_ (.Y(_08143_),
    .A(net5871),
    .B(_01795_));
 sg13g2_o21ai_1 _21756_ (.B1(_08143_),
    .Y(_08144_),
    .A1(net5871),
    .A2(_08142_));
 sg13g2_o21ai_1 _21757_ (.B1(net7927),
    .Y(_08145_),
    .A1(net7438),
    .A2(_08140_));
 sg13g2_mux2_1 _21758_ (.A0(_01794_),
    .A1(_07422_),
    .S(net5816),
    .X(_08146_));
 sg13g2_nor2b_1 _21759_ (.A(net7947),
    .B_N(net404),
    .Y(_08147_));
 sg13g2_a21oi_1 _21760_ (.A1(net7947),
    .A2(_01829_),
    .Y(_08148_),
    .B1(_08147_));
 sg13g2_nand2_2 _21761_ (.Y(_08149_),
    .A(net5873),
    .B(_01793_));
 sg13g2_o21ai_1 _21762_ (.B1(_08149_),
    .Y(_08150_),
    .A1(net5873),
    .A2(_08148_));
 sg13g2_nor2b_1 _21763_ (.A(net7943),
    .B_N(net403),
    .Y(_08151_));
 sg13g2_a21oi_1 _21764_ (.A1(net7943),
    .A2(_01828_),
    .Y(_08152_),
    .B1(_08151_));
 sg13g2_and2_1 _21765_ (.A(_08131_),
    .B(_08145_),
    .X(_08153_));
 sg13g2_nand2_1 _21766_ (.Y(_08154_),
    .A(_08131_),
    .B(_08145_));
 sg13g2_nand2_2 _21767_ (.Y(_08155_),
    .A(net5876),
    .B(_01792_));
 sg13g2_o21ai_1 _21768_ (.B1(_08155_),
    .Y(_08156_),
    .A1(net5876),
    .A2(_08152_));
 sg13g2_nor2b_1 _21769_ (.A(net7941),
    .B_N(net402),
    .Y(_08157_));
 sg13g2_nand2_1 _21770_ (.Y(_08158_),
    .A(_08010_),
    .B(_08153_));
 sg13g2_a21oi_1 _21771_ (.A1(net7941),
    .A2(_01826_),
    .Y(_08159_),
    .B1(_08157_));
 sg13g2_nor4_1 _21772_ (.A(_08012_),
    .B(_08071_),
    .C(_08125_),
    .D(_08154_),
    .Y(_08160_));
 sg13g2_nand2_2 _21773_ (.Y(_08161_),
    .A(net5870),
    .B(_01791_));
 sg13g2_o21ai_1 _21774_ (.B1(_08161_),
    .Y(_08162_),
    .A1(_08122_),
    .A2(_08159_));
 sg13g2_nor2b_1 _21775_ (.A(net7946),
    .B_N(net401),
    .Y(_08163_));
 sg13g2_a21oi_1 _21776_ (.A1(net7946),
    .A2(_01825_),
    .Y(_08164_),
    .B1(_08163_));
 sg13g2_nor3_1 _21777_ (.A(net7678),
    .B(_07978_),
    .C(_07982_),
    .Y(_08165_));
 sg13g2_nand2_2 _21778_ (.Y(_08166_),
    .A(net5878),
    .B(_01790_));
 sg13g2_o21ai_1 _21779_ (.B1(_08166_),
    .Y(_08167_),
    .A1(net5877),
    .A2(_08164_));
 sg13g2_nor2b_1 _21780_ (.A(net7945),
    .B_N(net400),
    .Y(_08168_));
 sg13g2_a21oi_1 _21781_ (.A1(net7945),
    .A2(_01824_),
    .Y(_08169_),
    .B1(_08168_));
 sg13g2_o21ai_1 _21782_ (.B1(_07970_),
    .Y(_08170_),
    .A1(_07694_),
    .A2(_08165_));
 sg13g2_nand2_2 _21783_ (.Y(_08171_),
    .A(net5878),
    .B(_01789_));
 sg13g2_o21ai_1 _21784_ (.B1(_08171_),
    .Y(_08172_),
    .A1(net5878),
    .A2(_08169_));
 sg13g2_nor2b_1 _21785_ (.A(net7946),
    .B_N(net399),
    .Y(_08173_));
 sg13g2_nand3_1 _21786_ (.B(net7438),
    .C(_07739_),
    .A(net7477),
    .Y(_08174_));
 sg13g2_a21oi_1 _21787_ (.A1(net7946),
    .A2(_01823_),
    .Y(_08175_),
    .B1(_08173_));
 sg13g2_and2_1 _21788_ (.A(_07616_),
    .B(_07649_),
    .X(_08176_));
 sg13g2_nand2_2 _21789_ (.Y(_08177_),
    .A(net5877),
    .B(_01788_));
 sg13g2_o21ai_1 _21790_ (.B1(_08177_),
    .Y(_08178_),
    .A1(net5877),
    .A2(_08175_));
 sg13g2_nor2b_1 _21791_ (.A(net7942),
    .B_N(net398),
    .Y(_08179_));
 sg13g2_a21oi_1 _21792_ (.A1(net7942),
    .A2(_01822_),
    .Y(_08180_),
    .B1(_08179_));
 sg13g2_a21oi_1 _21793_ (.A1(_07698_),
    .A2(_07982_),
    .Y(_08181_),
    .B1(net7678));
 sg13g2_nand2_2 _21794_ (.Y(_08182_),
    .A(net5877),
    .B(_01787_));
 sg13g2_o21ai_1 _21795_ (.B1(_08182_),
    .Y(_08183_),
    .A1(net5877),
    .A2(_08180_));
 sg13g2_nor2b_1 _21796_ (.A(net7943),
    .B_N(net397),
    .Y(_08184_));
 sg13g2_a21oi_1 _21797_ (.A1(net7943),
    .A2(_01821_),
    .Y(_08185_),
    .B1(_08184_));
 sg13g2_o21ai_1 _21798_ (.B1(_08176_),
    .Y(_08186_),
    .A1(_07669_),
    .A2(_08181_));
 sg13g2_nand2_2 _21799_ (.Y(_08187_),
    .A(net5875),
    .B(_01786_));
 sg13g2_o21ai_1 _21800_ (.B1(_08187_),
    .Y(_08188_),
    .A1(net5876),
    .A2(_08185_));
 sg13g2_nor2b_1 _21801_ (.A(net7939),
    .B_N(net395),
    .Y(_08189_));
 sg13g2_a21oi_1 _21802_ (.A1(net7939),
    .A2(_01820_),
    .Y(_08190_),
    .B1(_08189_));
 sg13g2_nand2_2 _21803_ (.Y(_08191_),
    .A(net5872),
    .B(_01785_));
 sg13g2_o21ai_1 _21804_ (.B1(_08191_),
    .Y(_08192_),
    .A1(net5873),
    .A2(_08190_));
 sg13g2_nor2b_1 _21805_ (.A(net7942),
    .B_N(net394),
    .Y(_08193_));
 sg13g2_a21oi_1 _21806_ (.A1(net7942),
    .A2(_01819_),
    .Y(_08194_),
    .B1(_08193_));
 sg13g2_and3_1 _21807_ (.X(_08195_),
    .A(_08170_),
    .B(_08174_),
    .C(_08186_));
 sg13g2_nand2_2 _21808_ (.Y(_08196_),
    .A(net5876),
    .B(_01784_));
 sg13g2_o21ai_1 _21809_ (.B1(_08196_),
    .Y(_08197_),
    .A1(net5876),
    .A2(_08194_));
 sg13g2_nand3_1 _21810_ (.B(_07649_),
    .C(_07665_),
    .A(_07616_),
    .Y(_08198_));
 sg13g2_mux2_1 _21811_ (.A0(_01783_),
    .A1(_07449_),
    .S(net5814),
    .X(_08199_));
 sg13g2_nor2b_1 _21812_ (.A(net7938),
    .B_N(net393),
    .Y(_08200_));
 sg13g2_a21oi_1 _21813_ (.A1(net7938),
    .A2(_01818_),
    .Y(_08201_),
    .B1(_08200_));
 sg13g2_a221oi_1 _21814_ (.B2(_07973_),
    .C1(_07701_),
    .B1(_08198_),
    .A1(net7921),
    .Y(_08202_),
    .A2(_07978_));
 sg13g2_nand2_2 _21815_ (.Y(_08203_),
    .A(net5869),
    .B(_01782_));
 sg13g2_o21ai_1 _21816_ (.B1(_08203_),
    .Y(_08204_),
    .A1(net5869),
    .A2(_08201_));
 sg13g2_inv_1 _21817_ (.Y(_08205_),
    .A(net7295));
 sg13g2_nor2b_1 _21818_ (.A(net7938),
    .B_N(net392),
    .Y(_08206_));
 sg13g2_a21oi_1 _21819_ (.A1(net7938),
    .A2(_01817_),
    .Y(_08207_),
    .B1(_08206_));
 sg13g2_a21oi_1 _21820_ (.A1(net7438),
    .A2(_08026_),
    .Y(_08208_),
    .B1(_08202_));
 sg13g2_nand2_2 _21821_ (.Y(_08209_),
    .A(net5869),
    .B(_01781_));
 sg13g2_o21ai_1 _21822_ (.B1(_08209_),
    .Y(_08210_),
    .A1(net5869),
    .A2(_08207_));
 sg13g2_nor2b_1 _21823_ (.A(net7944),
    .B_N(net391),
    .Y(_08211_));
 sg13g2_a21oi_1 _21824_ (.A1(net7944),
    .A2(_01815_),
    .Y(_08212_),
    .B1(_08211_));
 sg13g2_nor2b_1 _21825_ (.A(_08195_),
    .B_N(_08208_),
    .Y(_08213_));
 sg13g2_nand2_2 _21826_ (.Y(_08214_),
    .A(net5874),
    .B(_01780_));
 sg13g2_o21ai_1 _21827_ (.B1(_08214_),
    .Y(_08215_),
    .A1(net5875),
    .A2(_08212_));
 sg13g2_nor2b_1 _21828_ (.A(net7940),
    .B_N(net390),
    .Y(_08216_));
 sg13g2_a21oi_1 _21829_ (.A1(net7940),
    .A2(_01814_),
    .Y(_08217_),
    .B1(_08216_));
 sg13g2_nand2_2 _21830_ (.Y(_08218_),
    .A(net5871),
    .B(_01779_));
 sg13g2_o21ai_1 _21831_ (.B1(_08218_),
    .Y(_08219_),
    .A1(net5871),
    .A2(_08217_));
 sg13g2_nor2b_1 _21832_ (.A(net7941),
    .B_N(net389),
    .Y(_08220_));
 sg13g2_a21oi_1 _21833_ (.A1(net7941),
    .A2(_01813_),
    .Y(_08221_),
    .B1(_08220_));
 sg13g2_and2_1 _21834_ (.A(_08160_),
    .B(_08208_),
    .X(_08222_));
 sg13g2_nand2_2 _21835_ (.Y(_08223_),
    .A(net5870),
    .B(_01778_));
 sg13g2_o21ai_1 _21836_ (.B1(_08223_),
    .Y(_08224_),
    .A1(net5870),
    .A2(_08221_));
 sg13g2_nor2b_1 _21837_ (.A(net7939),
    .B_N(net388),
    .Y(_08225_));
 sg13g2_a21oi_1 _21838_ (.A1(net7939),
    .A2(_01812_),
    .Y(_08226_),
    .B1(_08225_));
 sg13g2_inv_1 _21839_ (.Y(_08227_),
    .A(_01926_));
 sg13g2_a21oi_1 _21840_ (.A1(_08160_),
    .A2(_08213_),
    .Y(_08228_),
    .B1(_08016_));
 sg13g2_nand2_2 _21841_ (.Y(_08229_),
    .A(net5871),
    .B(_01777_));
 sg13g2_o21ai_1 _21842_ (.B1(_08229_),
    .Y(_08230_),
    .A1(net5871),
    .A2(_08226_));
 sg13g2_nor2b_1 _21843_ (.A(net7939),
    .B_N(net387),
    .Y(_08231_));
 sg13g2_a21oi_1 _21844_ (.A1(net7947),
    .A2(_01811_),
    .Y(_08232_),
    .B1(_08231_));
 sg13g2_and2_1 _21845_ (.A(net7674),
    .B(_01903_),
    .X(_08233_));
 sg13g2_nand2_2 _21846_ (.Y(_08234_),
    .A(net5873),
    .B(_01776_));
 sg13g2_o21ai_1 _21847_ (.B1(_08234_),
    .Y(_08235_),
    .A1(net5873),
    .A2(_08232_));
 sg13g2_nor2b_1 _21848_ (.A(net7943),
    .B_N(net386),
    .Y(_08236_));
 sg13g2_a21oi_1 _21849_ (.A1(net7943),
    .A2(_01810_),
    .Y(_08237_),
    .B1(_08236_));
 sg13g2_nand4_1 _21850_ (.B(net7609),
    .C(_07608_),
    .A(net7610),
    .Y(_08238_),
    .D(_08233_));
 sg13g2_nor2_1 _21851_ (.A(_07815_),
    .B(_08238_),
    .Y(_08239_));
 sg13g2_nand2_2 _21852_ (.Y(_08240_),
    .A(net5875),
    .B(_01775_));
 sg13g2_o21ai_1 _21853_ (.B1(_08240_),
    .Y(_08241_),
    .A1(net5875),
    .A2(_08237_));
 sg13g2_or2_1 _21854_ (.X(_08242_),
    .B(_08238_),
    .A(_07815_));
 sg13g2_nor2b_1 _21855_ (.A(net7941),
    .B_N(net416),
    .Y(_08243_));
 sg13g2_a21oi_1 _21856_ (.A1(net7947),
    .A2(_01809_),
    .Y(_08244_),
    .B1(_08243_));
 sg13g2_nand2_2 _21857_ (.Y(_08245_),
    .A(_08122_),
    .B(_01774_));
 sg13g2_o21ai_1 _21858_ (.B1(_08245_),
    .Y(_08246_),
    .A1(net5870),
    .A2(_08244_));
 sg13g2_nor2b_1 _21859_ (.A(net7945),
    .B_N(net415),
    .Y(_08247_));
 sg13g2_a21oi_1 _21860_ (.A1(net7945),
    .A2(_01808_),
    .Y(_08248_),
    .B1(_08247_));
 sg13g2_nor3_1 _21861_ (.A(_08894_),
    .B(_07619_),
    .C(_07815_),
    .Y(_08249_));
 sg13g2_nand3_1 _21862_ (.B(_07616_),
    .C(_07812_),
    .A(net7684),
    .Y(_08250_));
 sg13g2_and2_1 _21863_ (.A(_08228_),
    .B(net7376),
    .X(_08251_));
 sg13g2_nand2_2 _21864_ (.Y(_08252_),
    .A(net5878),
    .B(_01773_));
 sg13g2_o21ai_1 _21865_ (.B1(_08252_),
    .Y(_08253_),
    .A1(net5879),
    .A2(_08248_));
 sg13g2_inv_1 _21866_ (.Y(_08254_),
    .A(_08251_));
 sg13g2_nor2b_1 _21867_ (.A(net7715),
    .B_N(net7696),
    .Y(_08255_));
 sg13g2_mux2_1 _21868_ (.A0(_01772_),
    .A1(_07465_),
    .S(net5814),
    .X(_08256_));
 sg13g2_nor2b_1 _21869_ (.A(net7945),
    .B_N(net414),
    .Y(_08257_));
 sg13g2_a21oi_1 _21870_ (.A1(net7945),
    .A2(_01807_),
    .Y(_08258_),
    .B1(_08257_));
 sg13g2_nand2_2 _21871_ (.Y(_08259_),
    .A(net5878),
    .B(_01771_));
 sg13g2_o21ai_1 _21872_ (.B1(_08259_),
    .Y(_08260_),
    .A1(net5878),
    .A2(_08258_));
 sg13g2_nor2b_1 _21873_ (.A(net7945),
    .B_N(net413),
    .Y(_08261_));
 sg13g2_a21oi_1 _21874_ (.A1(net7945),
    .A2(_01806_),
    .Y(_08262_),
    .B1(_08261_));
 sg13g2_nand2_2 _21875_ (.Y(_08263_),
    .A(net5878),
    .B(_01770_));
 sg13g2_o21ai_1 _21876_ (.B1(_08263_),
    .Y(_08264_),
    .A1(net5879),
    .A2(_08262_));
 sg13g2_nor2b_1 _21877_ (.A(net7942),
    .B_N(net412),
    .Y(_08265_));
 sg13g2_a21oi_1 _21878_ (.A1(net7942),
    .A2(_01804_),
    .Y(_08266_),
    .B1(_08265_));
 sg13g2_nand2_2 _21879_ (.Y(_08267_),
    .A(net5877),
    .B(_01769_));
 sg13g2_o21ai_1 _21880_ (.B1(_08267_),
    .Y(_08268_),
    .A1(net5877),
    .A2(_08266_));
 sg13g2_nor2b_1 _21881_ (.A(net7944),
    .B_N(net411),
    .Y(_08269_));
 sg13g2_a21oi_1 _21882_ (.A1(net7944),
    .A2(_01803_),
    .Y(_08270_),
    .B1(_08269_));
 sg13g2_nand2_2 _21883_ (.Y(_08271_),
    .A(net5875),
    .B(_01768_));
 sg13g2_o21ai_1 _21884_ (.B1(_08271_),
    .Y(_08272_),
    .A1(net5875),
    .A2(_08270_));
 sg13g2_nor2b_1 _21885_ (.A(net7939),
    .B_N(net410),
    .Y(_08273_));
 sg13g2_a21oi_1 _21886_ (.A1(net7939),
    .A2(_01802_),
    .Y(_08274_),
    .B1(_08273_));
 sg13g2_nand2_2 _21887_ (.Y(_08275_),
    .A(net5872),
    .B(_01767_));
 sg13g2_o21ai_1 _21888_ (.B1(_08275_),
    .Y(_08276_),
    .A1(net5873),
    .A2(_08274_));
 sg13g2_nor2b_1 _21889_ (.A(net7942),
    .B_N(net407),
    .Y(_08277_));
 sg13g2_a21oi_1 _21890_ (.A1(net7942),
    .A2(_01801_),
    .Y(_08278_),
    .B1(_08277_));
 sg13g2_mux4_1 _21891_ (.S0(net7761),
    .A0(_00788_),
    .A1(_00820_),
    .A2(_00852_),
    .A3(_00887_),
    .S1(net7732),
    .X(_08279_));
 sg13g2_nand2_2 _21892_ (.Y(_08280_),
    .A(net5876),
    .B(_01766_));
 sg13g2_o21ai_1 _21893_ (.B1(_08280_),
    .Y(_08281_),
    .A1(net5876),
    .A2(_08278_));
 sg13g2_and2_1 _21894_ (.A(net7606),
    .B(_08279_),
    .X(_08282_));
 sg13g2_nor2b_1 _21895_ (.A(net7938),
    .B_N(net396),
    .Y(_08283_));
 sg13g2_a21oi_1 _21896_ (.A1(net7938),
    .A2(_01800_),
    .Y(_08284_),
    .B1(_08283_));
 sg13g2_nand2b_1 _21897_ (.Y(_08285_),
    .B(net7732),
    .A_N(_01901_));
 sg13g2_nand2_2 _21898_ (.Y(_08286_),
    .A(net5869),
    .B(_01765_));
 sg13g2_o21ai_1 _21899_ (.B1(_08286_),
    .Y(_08287_),
    .A1(_08122_),
    .A2(_08284_));
 sg13g2_nor2_1 _21900_ (.A(_09041_),
    .B(_08285_),
    .Y(_08288_));
 sg13g2_nor2b_1 _21901_ (.A(net7938),
    .B_N(net385),
    .Y(_08289_));
 sg13g2_a21oi_1 _21902_ (.A1(net7938),
    .A2(_01799_),
    .Y(_08290_),
    .B1(_08289_));
 sg13g2_nand3b_1 _21903_ (.B(net7743),
    .C(net7803),
    .Y(_08291_),
    .A_N(net7695));
 sg13g2_nand2_1 _21904_ (.Y(_08292_),
    .A(net7699),
    .B(_00756_));
 sg13g2_nand2_2 _21905_ (.Y(_08293_),
    .A(net5869),
    .B(_01764_));
 sg13g2_o21ai_1 _21906_ (.B1(_08293_),
    .Y(_08294_),
    .A1(net5869),
    .A2(_08290_));
 sg13g2_nor2_1 _21907_ (.A(_01763_),
    .B(net5815),
    .Y(_08295_));
 sg13g2_nor2b_1 _21908_ (.A(net7951),
    .B_N(net409),
    .Y(_08296_));
 sg13g2_a21oi_1 _21909_ (.A1(net7951),
    .A2(_01798_),
    .Y(_08297_),
    .B1(_08296_));
 sg13g2_nand2b_1 _21910_ (.Y(_08298_),
    .B(_01566_),
    .A_N(net7699));
 sg13g2_a21oi_1 _21911_ (.A1(net5815),
    .A2(_08297_),
    .Y(_08299_),
    .B1(_08295_));
 sg13g2_a21oi_1 _21912_ (.A1(_08292_),
    .A2(_08298_),
    .Y(_08300_),
    .B1(net7601));
 sg13g2_nor2_1 _21913_ (.A(_01762_),
    .B(net5813),
    .Y(_08301_));
 sg13g2_nor2b_1 _21914_ (.A(net7950),
    .B_N(net408),
    .Y(_08302_));
 sg13g2_a21oi_1 _21915_ (.A1(net7950),
    .A2(_01797_),
    .Y(_08303_),
    .B1(_08302_));
 sg13g2_a21oi_1 _21916_ (.A1(net5813),
    .A2(_08303_),
    .Y(_08304_),
    .B1(_08301_));
 sg13g2_nor2_1 _21917_ (.A(_01901_),
    .B(net7717),
    .Y(_08305_));
 sg13g2_or2_1 _21918_ (.X(_08306_),
    .B(net7702),
    .A(net7693));
 sg13g2_nor2b_1 _21919_ (.A(net7734),
    .B_N(_01898_),
    .Y(_08307_));
 sg13g2_mux2_1 _21920_ (.A0(_01761_),
    .A1(_07476_),
    .S(net5816),
    .X(_08308_));
 sg13g2_nor2_1 _21921_ (.A(_01760_),
    .B(net5812),
    .Y(_08309_));
 sg13g2_nor2b_1 _21922_ (.A(net7955),
    .B_N(net406),
    .Y(_08310_));
 sg13g2_a21oi_1 _21923_ (.A1(net7955),
    .A2(_01796_),
    .Y(_08311_),
    .B1(_08310_));
 sg13g2_nand3b_1 _21924_ (.B(net7762),
    .C(_00862_),
    .Y(_08312_),
    .A_N(net7733));
 sg13g2_nor2b_1 _21925_ (.A(_01898_),
    .B_N(_01899_),
    .Y(_08313_));
 sg13g2_a21oi_1 _21926_ (.A1(net5812),
    .A2(_08311_),
    .Y(_08314_),
    .B1(_08309_));
 sg13g2_nor2_1 _21927_ (.A(_01759_),
    .B(net5813),
    .Y(_08315_));
 sg13g2_nor2b_1 _21928_ (.A(net7950),
    .B_N(net405),
    .Y(_08316_));
 sg13g2_a21oi_1 _21929_ (.A1(net7950),
    .A2(_01795_),
    .Y(_08317_),
    .B1(_08316_));
 sg13g2_nand3b_1 _21930_ (.B(_01214_),
    .C(net7733),
    .Y(_08318_),
    .A_N(net7761));
 sg13g2_a21oi_1 _21931_ (.A1(net5813),
    .A2(_08317_),
    .Y(_08319_),
    .B1(_08315_));
 sg13g2_nor2_1 _21932_ (.A(_01758_),
    .B(net5814),
    .Y(_08320_));
 sg13g2_nor2b_1 _21933_ (.A(net7951),
    .B_N(net404),
    .Y(_08321_));
 sg13g2_a21oi_1 _21934_ (.A1(net7951),
    .A2(_01793_),
    .Y(_08322_),
    .B1(_08321_));
 sg13g2_a21oi_1 _21935_ (.A1(_08312_),
    .A2(_08318_),
    .Y(_08323_),
    .B1(_08306_));
 sg13g2_a21oi_1 _21936_ (.A1(net5814),
    .A2(_08322_),
    .Y(_08324_),
    .B1(_08320_));
 sg13g2_nor2_1 _21937_ (.A(_01757_),
    .B(net5815),
    .Y(_08325_));
 sg13g2_nor2b_1 _21938_ (.A(net7954),
    .B_N(net403),
    .Y(_08326_));
 sg13g2_a21oi_1 _21939_ (.A1(net7954),
    .A2(_01792_),
    .Y(_08327_),
    .B1(_08326_));
 sg13g2_nor4_1 _21940_ (.A(net7689),
    .B(_08282_),
    .C(_08300_),
    .D(_08323_),
    .Y(_08328_));
 sg13g2_a21oi_1 _21941_ (.A1(net5815),
    .A2(_08327_),
    .Y(_08329_),
    .B1(_08325_));
 sg13g2_nor2_1 _21942_ (.A(_01756_),
    .B(net5812),
    .Y(_08330_));
 sg13g2_nor2b_1 _21943_ (.A(net7948),
    .B_N(net402),
    .Y(_08331_));
 sg13g2_a21oi_1 _21944_ (.A1(net7948),
    .A2(_01791_),
    .Y(_08332_),
    .B1(_08331_));
 sg13g2_a21oi_1 _21945_ (.A1(net5812),
    .A2(_08332_),
    .Y(_08333_),
    .B1(_08330_));
 sg13g2_nor2_1 _21946_ (.A(_01755_),
    .B(net5818),
    .Y(_08334_));
 sg13g2_mux2_1 _21947_ (.A0(_00660_),
    .A1(_00692_),
    .S(net7760),
    .X(_08335_));
 sg13g2_nor2b_1 _21948_ (.A(net7952),
    .B_N(net401),
    .Y(_08336_));
 sg13g2_a21oi_1 _21949_ (.A1(net7952),
    .A2(_01790_),
    .Y(_08337_),
    .B1(_08336_));
 sg13g2_a21oi_1 _21950_ (.A1(net5817),
    .A2(_08337_),
    .Y(_08338_),
    .B1(_08334_));
 sg13g2_nor2_1 _21951_ (.A(_01754_),
    .B(net5818),
    .Y(_08339_));
 sg13g2_nor2b_1 _21952_ (.A(net7952),
    .B_N(net400),
    .Y(_08340_));
 sg13g2_a21oi_1 _21953_ (.A1(net7952),
    .A2(_01789_),
    .Y(_08341_),
    .B1(_08340_));
 sg13g2_a21oi_1 _21954_ (.A1(net5818),
    .A2(_08341_),
    .Y(_08342_),
    .B1(_08339_));
 sg13g2_nor2_1 _21955_ (.A(_01753_),
    .B(net5818),
    .Y(_08343_));
 sg13g2_nor2b_1 _21956_ (.A(net7952),
    .B_N(net399),
    .Y(_08344_));
 sg13g2_a21oi_1 _21957_ (.A1(net7952),
    .A2(_01788_),
    .Y(_08345_),
    .B1(_08344_));
 sg13g2_a21oi_1 _21958_ (.A1(net5817),
    .A2(_08345_),
    .Y(_08346_),
    .B1(_08343_));
 sg13g2_nor2_1 _21959_ (.A(_01752_),
    .B(net5816),
    .Y(_08347_));
 sg13g2_nor2b_1 _21960_ (.A(net7953),
    .B_N(net398),
    .Y(_08348_));
 sg13g2_a21oi_1 _21961_ (.A1(net7953),
    .A2(_01787_),
    .Y(_08349_),
    .B1(_08348_));
 sg13g2_a221oi_1 _21962_ (.B2(_09011_),
    .C1(net7692),
    .B1(_08335_),
    .A1(_00724_),
    .Y(_08350_),
    .A2(net7593));
 sg13g2_a21oi_1 _21963_ (.A1(net5816),
    .A2(_08349_),
    .Y(_08351_),
    .B1(_08347_));
 sg13g2_nor2_1 _21964_ (.A(_01751_),
    .B(net5816),
    .Y(_08352_));
 sg13g2_nor2b_1 _21965_ (.A(net7954),
    .B_N(net397),
    .Y(_08353_));
 sg13g2_a21oi_1 _21966_ (.A1(net7954),
    .A2(_01786_),
    .Y(_08354_),
    .B1(_08353_));
 sg13g2_a21oi_1 _21967_ (.A1(net5816),
    .A2(_08354_),
    .Y(_08355_),
    .B1(_08352_));
 sg13g2_mux2_1 _21968_ (.A0(_01750_),
    .A1(_07500_),
    .S(net5810),
    .X(_08356_));
 sg13g2_nor2_1 _21969_ (.A(_01749_),
    .B(net5813),
    .Y(_08357_));
 sg13g2_nor2b_1 _21970_ (.A(net7951),
    .B_N(net395),
    .Y(_08358_));
 sg13g2_a21oi_1 _21971_ (.A1(net7951),
    .A2(_01785_),
    .Y(_08359_),
    .B1(_08358_));
 sg13g2_a21oi_1 _21972_ (.A1(net5815),
    .A2(_08359_),
    .Y(_08360_),
    .B1(_08357_));
 sg13g2_nor2_1 _21973_ (.A(_01748_),
    .B(net5815),
    .Y(_08361_));
 sg13g2_nor2b_1 _21974_ (.A(net7953),
    .B_N(net394),
    .Y(_08362_));
 sg13g2_a21oi_1 _21975_ (.A1(net7953),
    .A2(_01784_),
    .Y(_08363_),
    .B1(_08362_));
 sg13g2_a21oi_1 _21976_ (.A1(net5815),
    .A2(_08363_),
    .Y(_08364_),
    .B1(_08361_));
 sg13g2_nor2_1 _21977_ (.A(_01747_),
    .B(net5810),
    .Y(_08365_));
 sg13g2_nor2b_1 _21978_ (.A(net7949),
    .B_N(net393),
    .Y(_08366_));
 sg13g2_a21oi_1 _21979_ (.A1(net7949),
    .A2(_01782_),
    .Y(_08367_),
    .B1(_08366_));
 sg13g2_a21oi_1 _21980_ (.A1(net5810),
    .A2(_08367_),
    .Y(_08368_),
    .B1(_08365_));
 sg13g2_nor2_1 _21981_ (.A(_01746_),
    .B(net5810),
    .Y(_08369_));
 sg13g2_nor2b_1 _21982_ (.A(net7949),
    .B_N(net392),
    .Y(_08370_));
 sg13g2_a21oi_1 _21983_ (.A1(net7949),
    .A2(_01781_),
    .Y(_08371_),
    .B1(_08370_));
 sg13g2_a21oi_1 _21984_ (.A1(net5810),
    .A2(_08371_),
    .Y(_08372_),
    .B1(_08369_));
 sg13g2_mux4_1 _21985_ (.S0(net7761),
    .A0(_00922_),
    .A1(_00957_),
    .A2(_00992_),
    .A3(_01028_),
    .S1(net7732),
    .X(_08373_));
 sg13g2_mux2_1 _21986_ (.A0(_01745_),
    .A1(_07253_),
    .S(net5814),
    .X(_08374_));
 sg13g2_mux2_1 _21987_ (.A0(_01744_),
    .A1(_07264_),
    .S(net5812),
    .X(_08375_));
 sg13g2_o21ai_1 _21988_ (.B1(net7700),
    .Y(_08376_),
    .A1(_08946_),
    .A2(_08373_));
 sg13g2_nor2_1 _21989_ (.A(_01743_),
    .B(net5811),
    .Y(_08377_));
 sg13g2_a21oi_1 _21990_ (.A1(net5811),
    .A2(_07287_),
    .Y(_08378_),
    .B1(_08377_));
 sg13g2_nor2_1 _21991_ (.A(_01742_),
    .B(net5813),
    .Y(_08379_));
 sg13g2_a21oi_1 _21992_ (.A1(net5813),
    .A2(_07301_),
    .Y(_08380_),
    .B1(_08379_));
 sg13g2_o21ai_1 _21993_ (.B1(_08328_),
    .Y(_08381_),
    .A1(_08376_),
    .A2(_08350_));
 sg13g2_mux2_1 _21994_ (.A0(_01741_),
    .A1(_07317_),
    .S(net5814),
    .X(_08382_));
 sg13g2_nor2_1 _21995_ (.A(_01740_),
    .B(net5814),
    .Y(_08383_));
 sg13g2_nor2b_1 _21996_ (.A(net7697),
    .B_N(net7691),
    .Y(_08384_));
 sg13g2_nand2b_1 _21997_ (.Y(_08385_),
    .B(_01902_),
    .A_N(net7697));
 sg13g2_a21oi_1 _21998_ (.A1(net5814),
    .A2(_07337_),
    .Y(_08386_),
    .B1(_08383_));
 sg13g2_nor2_1 _21999_ (.A(net7712),
    .B(_08385_),
    .Y(_08387_));
 sg13g2_nor2_1 _22000_ (.A(_01739_),
    .B(net5810),
    .Y(_08388_));
 sg13g2_nand2b_1 _22001_ (.Y(_08389_),
    .B(net7590),
    .A_N(net7703));
 sg13g2_a21oi_1 _22002_ (.A1(net5810),
    .A2(_07514_),
    .Y(_08390_),
    .B1(_08388_));
 sg13g2_and4_1 _22003_ (.A(_01733_),
    .B(_01732_),
    .C(_01729_),
    .D(_08065_),
    .X(_08391_));
 sg13g2_and2_1 _22004_ (.A(_01734_),
    .B(_08391_),
    .X(_08392_));
 sg13g2_and4_1 _22005_ (.A(_01737_),
    .B(_01736_),
    .C(_01735_),
    .D(_08392_),
    .X(_08393_));
 sg13g2_and2_1 _22006_ (.A(_01738_),
    .B(_08393_),
    .X(_08394_));
 sg13g2_and2_1 _22007_ (.A(net5940),
    .B(_08394_),
    .X(_08395_));
 sg13g2_nand2_1 _22008_ (.Y(_08396_),
    .A(_07045_),
    .B(net6776));
 sg13g2_nand2_1 _22009_ (.Y(_08397_),
    .A(net5940),
    .B(_08393_));
 sg13g2_xor2_1 _22010_ (.B(_08397_),
    .A(_01738_),
    .X(_08398_));
 sg13g2_o21ai_1 _22011_ (.B1(_07707_),
    .Y(_08399_),
    .A1(net6762),
    .A2(_08398_));
 sg13g2_and2_1 _22012_ (.A(net5940),
    .B(_08392_),
    .X(_08400_));
 sg13g2_and2_1 _22013_ (.A(_01735_),
    .B(_08400_),
    .X(_08401_));
 sg13g2_nand2_1 _22014_ (.Y(_08402_),
    .A(_01736_),
    .B(_08401_));
 sg13g2_xor2_1 _22015_ (.B(_08402_),
    .A(_01737_),
    .X(_08403_));
 sg13g2_o21ai_1 _22016_ (.B1(_07722_),
    .Y(_08404_),
    .A1(net6762),
    .A2(_08403_));
 sg13g2_xnor2_1 _22017_ (.Y(_08405_),
    .A(_01736_),
    .B(_08401_));
 sg13g2_a21oi_1 _22018_ (.A1(net6771),
    .A2(_08405_),
    .Y(_08406_),
    .B1(_07729_));
 sg13g2_xnor2_1 _22019_ (.Y(_08407_),
    .A(_01735_),
    .B(_08400_));
 sg13g2_a21oi_1 _22020_ (.A1(net6771),
    .A2(_08407_),
    .Y(_08408_),
    .B1(_07740_));
 sg13g2_nor2_1 _22021_ (.A(_07093_),
    .B(_08400_),
    .Y(_08409_));
 sg13g2_nor2_1 _22022_ (.A(_01734_),
    .B(_08396_),
    .Y(_08410_));
 sg13g2_or2_1 _22023_ (.X(_08411_),
    .B(_08391_),
    .A(_01734_));
 sg13g2_a22oi_1 _22024_ (.Y(_08412_),
    .B1(_08409_),
    .B2(_08411_),
    .A2(_07754_),
    .A1(_07744_));
 sg13g2_nor2_1 _22025_ (.A(_08410_),
    .B(_08412_),
    .Y(_08413_));
 sg13g2_inv_1 _22026_ (.Y(_08414_),
    .A(_01918_));
 sg13g2_nand2_1 _22027_ (.Y(_08415_),
    .A(_01729_),
    .B(_08066_));
 sg13g2_nand3_1 _22028_ (.B(_01729_),
    .C(_08066_),
    .A(_01732_),
    .Y(_08416_));
 sg13g2_mux4_1 _22029_ (.S0(net7749),
    .A0(_01063_),
    .A1(_01098_),
    .A2(_01133_),
    .A3(_01168_),
    .S1(net7721),
    .X(_08417_));
 sg13g2_xor2_1 _22030_ (.B(_08416_),
    .A(_01733_),
    .X(_08418_));
 sg13g2_a21oi_1 _22031_ (.A1(net6771),
    .A2(_08418_),
    .Y(_08419_),
    .B1(_07767_));
 sg13g2_nand2b_1 _22032_ (.Y(_08420_),
    .B(net7433),
    .A_N(_08417_));
 sg13g2_xor2_1 _22033_ (.B(_08415_),
    .A(_01732_),
    .X(_08421_));
 sg13g2_a21oi_1 _22034_ (.A1(net6771),
    .A2(_08421_),
    .Y(_08422_),
    .B1(_07793_));
 sg13g2_nand3_1 _22035_ (.B(_01717_),
    .C(_01716_),
    .A(_01719_),
    .Y(_08423_));
 sg13g2_nand3b_1 _22036_ (.B(net7712),
    .C(net7691),
    .Y(_08424_),
    .A_N(net7697));
 sg13g2_and4_1 _22037_ (.A(_01711_),
    .B(_01710_),
    .C(_01709_),
    .D(_01708_),
    .X(_08425_));
 sg13g2_and4_1 _22038_ (.A(_01714_),
    .B(_01713_),
    .C(_01712_),
    .D(_08425_),
    .X(_08426_));
 sg13g2_nand3_1 _22039_ (.B(_08394_),
    .C(_08426_),
    .A(_01715_),
    .Y(_08427_));
 sg13g2_nor2_1 _22040_ (.A(_08423_),
    .B(_08427_),
    .Y(_08428_));
 sg13g2_nand3_1 _22041_ (.B(_01720_),
    .C(_08428_),
    .A(_01721_),
    .Y(_08429_));
 sg13g2_nor2_1 _22042_ (.A(_15030_),
    .B(_08429_),
    .Y(_08430_));
 sg13g2_and2_1 _22043_ (.A(_01723_),
    .B(_08430_),
    .X(_08431_));
 sg13g2_nand2_1 _22044_ (.Y(_08432_),
    .A(_01724_),
    .B(_08431_));
 sg13g2_nand3_1 _22045_ (.B(_01726_),
    .C(_01725_),
    .A(_01727_),
    .Y(_08433_));
 sg13g2_nor2_1 _22046_ (.A(_08432_),
    .B(_08433_),
    .Y(_08434_));
 sg13g2_nor3_1 _22047_ (.A(_14860_),
    .B(_08432_),
    .C(_08433_),
    .Y(_08435_));
 sg13g2_nand2_1 _22048_ (.Y(_08436_),
    .A(_01730_),
    .B(_08435_));
 sg13g2_nand2_1 _22049_ (.Y(_08437_),
    .A(_07803_),
    .B(_08436_));
 sg13g2_nand2_1 _22050_ (.Y(_08438_),
    .A(net5868),
    .B(_08437_));
 sg13g2_nand3_1 _22051_ (.B(net5938),
    .C(_08435_),
    .A(_01730_),
    .Y(_08439_));
 sg13g2_o21ai_1 _22052_ (.B1(net6769),
    .Y(_08440_),
    .A1(_14784_),
    .A2(_08439_));
 sg13g2_a22oi_1 _22053_ (.Y(_08441_),
    .B1(_08440_),
    .B2(_07803_),
    .A2(_08438_),
    .A1(_14784_));
 sg13g2_o21ai_1 _22054_ (.B1(net5868),
    .Y(_08442_),
    .A1(_07817_),
    .A2(_08435_));
 sg13g2_a21oi_1 _22055_ (.A1(net6769),
    .A2(_08439_),
    .Y(_08443_),
    .B1(_07817_));
 sg13g2_inv_1 _22056_ (.Y(_08444_),
    .A(net7665));
 sg13g2_a21oi_1 _22057_ (.A1(_14814_),
    .A2(_08442_),
    .Y(_08445_),
    .B1(_08443_));
 sg13g2_nand2_1 _22058_ (.Y(_08446_),
    .A(_07843_),
    .B(_08064_));
 sg13g2_a21oi_1 _22059_ (.A1(_08396_),
    .A2(_08446_),
    .Y(_08447_),
    .B1(_01729_));
 sg13g2_nand2_1 _22060_ (.Y(_08448_),
    .A(net6771),
    .B(_08415_));
 sg13g2_a21oi_1 _22061_ (.A1(_07843_),
    .A2(_08448_),
    .Y(_08449_),
    .B1(_08447_));
 sg13g2_o21ai_1 _22062_ (.B1(net5868),
    .Y(_08450_),
    .A1(_07853_),
    .A2(_08434_));
 sg13g2_a21oi_1 _22063_ (.A1(net5938),
    .A2(_08435_),
    .Y(_08451_),
    .B1(net6767));
 sg13g2_nor2_1 _22064_ (.A(_07853_),
    .B(_08451_),
    .Y(_08452_));
 sg13g2_a21oi_1 _22065_ (.A1(_14860_),
    .A2(_08450_),
    .Y(_08453_),
    .B1(_08452_));
 sg13g2_nor2_1 _22066_ (.A(_07045_),
    .B(_08432_),
    .Y(_08454_));
 sg13g2_nand3_1 _22067_ (.B(_01725_),
    .C(_08454_),
    .A(_01726_),
    .Y(_08455_));
 sg13g2_mux4_1 _22068_ (.S0(net7749),
    .A0(_01204_),
    .A1(_01239_),
    .A2(_01274_),
    .A3(_01309_),
    .S1(net7721),
    .X(_08456_));
 sg13g2_xnor2_1 _22069_ (.Y(_08457_),
    .A(_01727_),
    .B(_08455_));
 sg13g2_a21o_1 _22070_ (.A2(_08457_),
    .A1(net6769),
    .B1(_07862_),
    .X(_08458_));
 sg13g2_nand2_1 _22071_ (.Y(_08459_),
    .A(_01725_),
    .B(_08454_));
 sg13g2_or2_1 _22072_ (.X(_08460_),
    .B(_08456_),
    .A(net7586));
 sg13g2_xor2_1 _22073_ (.B(_08459_),
    .A(_01726_),
    .X(_08461_));
 sg13g2_nand2_1 _22074_ (.Y(_08462_),
    .A(_01902_),
    .B(net7697));
 sg13g2_o21ai_1 _22075_ (.B1(_07873_),
    .Y(_08463_),
    .A1(net6763),
    .A2(_08461_));
 sg13g2_nand2b_1 _22076_ (.Y(_08464_),
    .B(net7744),
    .A_N(net7715));
 sg13g2_xor2_1 _22077_ (.B(_08454_),
    .A(_01725_),
    .X(_08465_));
 sg13g2_a21o_1 _22078_ (.A2(_08465_),
    .A1(net6769),
    .B1(_07882_),
    .X(_08466_));
 sg13g2_nor2_1 _22079_ (.A(net6763),
    .B(_08454_),
    .Y(_08467_));
 sg13g2_nor2_1 _22080_ (.A(_01724_),
    .B(net5868),
    .Y(_08468_));
 sg13g2_or2_1 _22081_ (.X(_08469_),
    .B(_08431_),
    .A(_01724_));
 sg13g2_a21oi_1 _22082_ (.A1(_08467_),
    .A2(_08469_),
    .Y(_08470_),
    .B1(_07892_));
 sg13g2_nor2_1 _22083_ (.A(_08468_),
    .B(_08470_),
    .Y(_08471_));
 sg13g2_nand2_1 _22084_ (.Y(_08472_),
    .A(net5938),
    .B(_08430_));
 sg13g2_xor2_1 _22085_ (.B(_08472_),
    .A(_01723_),
    .X(_08473_));
 sg13g2_o21ai_1 _22086_ (.B1(_07902_),
    .Y(_08474_),
    .A1(net6763),
    .A2(_08473_));
 sg13g2_nand2b_1 _22087_ (.Y(_08475_),
    .B(_08429_),
    .A_N(_07912_));
 sg13g2_a21oi_1 _22088_ (.A1(net5868),
    .A2(_08475_),
    .Y(_08476_),
    .B1(_01722_));
 sg13g2_a21oi_1 _22089_ (.A1(net6769),
    .A2(_08472_),
    .Y(_08477_),
    .B1(_07912_));
 sg13g2_nor2_1 _22090_ (.A(_08476_),
    .B(_08477_),
    .Y(_08478_));
 sg13g2_mux2_1 _22091_ (.A0(_01415_),
    .A1(_01450_),
    .S(net7757),
    .X(_08479_));
 sg13g2_nand3_1 _22092_ (.B(_01720_),
    .C(_08428_),
    .A(net5939),
    .Y(_08480_));
 sg13g2_nor3_1 _22093_ (.A(net7584),
    .B(net7568),
    .C(_08479_),
    .Y(_08481_));
 sg13g2_xnor2_1 _22094_ (.Y(_08482_),
    .A(_01721_),
    .B(_08480_));
 sg13g2_a21o_1 _22095_ (.A2(_08482_),
    .A1(net6770),
    .B1(_07921_),
    .X(_08483_));
 sg13g2_o21ai_1 _22096_ (.B1(net5868),
    .Y(_08484_),
    .A1(_07931_),
    .A2(_08428_));
 sg13g2_nand2b_1 _22097_ (.Y(_08485_),
    .B(net7714),
    .A_N(net7744));
 sg13g2_a21oi_1 _22098_ (.A1(net6770),
    .A2(_08480_),
    .Y(_08486_),
    .B1(_07931_));
 sg13g2_a21oi_1 _22099_ (.A1(_15108_),
    .A2(_08484_),
    .Y(_08487_),
    .B1(_08486_));
 sg13g2_nor2_1 _22100_ (.A(_07045_),
    .B(_08427_),
    .Y(_08488_));
 sg13g2_nand3_1 _22101_ (.B(_01716_),
    .C(_08488_),
    .A(_01717_),
    .Y(_08489_));
 sg13g2_xnor2_1 _22102_ (.Y(_08490_),
    .A(_01719_),
    .B(_08489_));
 sg13g2_a21o_1 _22103_ (.A2(_08490_),
    .A1(net6769),
    .B1(_07941_),
    .X(_08491_));
 sg13g2_o21ai_1 _22104_ (.B1(net7976),
    .Y(_08492_),
    .A1(_07012_),
    .A2(net5922));
 sg13g2_a21oi_1 _22105_ (.A1(net5953),
    .A2(_08064_),
    .Y(_08493_),
    .B1(_07093_));
 sg13g2_nand2_1 _22106_ (.Y(_08494_),
    .A(\alu_adder_result_ex[1] ),
    .B(net6886));
 sg13g2_a221oi_1 _22107_ (.B2(_00259_),
    .C1(net6770),
    .B1(_07695_),
    .A1(_00361_),
    .Y(_08495_),
    .A2(_07686_));
 sg13g2_a22oi_1 _22108_ (.Y(_08496_),
    .B1(_08494_),
    .B2(_08495_),
    .A2(_08493_),
    .A1(_08492_));
 sg13g2_mux2_1 _22109_ (.A0(_01485_),
    .A1(_01520_),
    .S(net7756),
    .X(_08497_));
 sg13g2_nor3_1 _22110_ (.A(net7584),
    .B(net7565),
    .C(_08497_),
    .Y(_08498_));
 sg13g2_nand2_1 _22111_ (.Y(_08499_),
    .A(_01716_),
    .B(_08488_));
 sg13g2_xnor2_1 _22112_ (.Y(_08500_),
    .A(_01717_),
    .B(_08499_));
 sg13g2_a21o_1 _22113_ (.A2(_08500_),
    .A1(net6769),
    .B1(_07951_),
    .X(_08501_));
 sg13g2_xor2_1 _22114_ (.B(_08488_),
    .A(_01716_),
    .X(_08502_));
 sg13g2_or2_1 _22115_ (.X(_08503_),
    .B(net7731),
    .A(net7706));
 sg13g2_a21o_1 _22116_ (.A2(_08502_),
    .A1(net6769),
    .B1(_07962_),
    .X(_08504_));
 sg13g2_a21o_1 _22117_ (.A2(_08426_),
    .A1(_08394_),
    .B1(_07974_),
    .X(_08505_));
 sg13g2_a21oi_1 _22118_ (.A1(net5868),
    .A2(_08505_),
    .Y(_08506_),
    .B1(_01715_));
 sg13g2_nand4_1 _22119_ (.B(net5935),
    .C(_08394_),
    .A(_01715_),
    .Y(_08507_),
    .D(_08426_));
 sg13g2_a21oi_1 _22120_ (.A1(net6770),
    .A2(_08507_),
    .Y(_08508_),
    .B1(_07974_));
 sg13g2_nor2_1 _22121_ (.A(_08506_),
    .B(_08508_),
    .Y(_08509_));
 sg13g2_inv_1 _22122_ (.Y(_08510_),
    .A(_01915_));
 sg13g2_nand2_1 _22123_ (.Y(_08511_),
    .A(_08395_),
    .B(_08425_));
 sg13g2_nand4_1 _22124_ (.B(_01712_),
    .C(_08395_),
    .A(_01713_),
    .Y(_08512_),
    .D(_08425_));
 sg13g2_xnor2_1 _22125_ (.Y(_08513_),
    .A(_01714_),
    .B(_08512_));
 sg13g2_a21o_1 _22126_ (.A2(_08513_),
    .A1(net6771),
    .B1(_07986_),
    .X(_08514_));
 sg13g2_nand3_1 _22127_ (.B(_08395_),
    .C(_08425_),
    .A(_01712_),
    .Y(_08515_));
 sg13g2_mux2_1 _22128_ (.A0(_01344_),
    .A1(_01380_),
    .S(net7757),
    .X(_08516_));
 sg13g2_xor2_1 _22129_ (.B(_08515_),
    .A(_01713_),
    .X(_08517_));
 sg13g2_o21ai_1 _22130_ (.B1(_07996_),
    .Y(_08518_),
    .A1(net6767),
    .A2(_08517_));
 sg13g2_nor3_1 _22131_ (.A(net7584),
    .B(net7560),
    .C(_08516_),
    .Y(_08519_));
 sg13g2_xor2_1 _22132_ (.B(_08511_),
    .A(_01712_),
    .X(_08520_));
 sg13g2_o21ai_1 _22133_ (.B1(_08006_),
    .Y(_08521_),
    .A1(net6760),
    .A2(_08520_));
 sg13g2_nand2_1 _22134_ (.Y(_08522_),
    .A(net7711),
    .B(net7745));
 sg13g2_nand4_1 _22135_ (.B(_01709_),
    .C(_01708_),
    .A(_01710_),
    .Y(_08523_),
    .D(_08394_));
 sg13g2_nand2b_1 _22136_ (.Y(_08524_),
    .B(_08523_),
    .A_N(net6554));
 sg13g2_a21oi_1 _22137_ (.A1(net5868),
    .A2(_08524_),
    .Y(_08525_),
    .B1(_01711_));
 sg13g2_a21oi_1 _22138_ (.A1(net6771),
    .A2(_08511_),
    .Y(_08526_),
    .B1(net6554));
 sg13g2_nand4_1 _22139_ (.B(net7697),
    .C(net7712),
    .A(net7691),
    .Y(_08527_),
    .D(net7747));
 sg13g2_nor2_1 _22140_ (.A(_08525_),
    .B(_08526_),
    .Y(_08528_));
 sg13g2_nand2_1 _22141_ (.Y(_08529_),
    .A(_01708_),
    .B(_08395_));
 sg13g2_nand3_1 _22142_ (.B(_01708_),
    .C(_08395_),
    .A(_01709_),
    .Y(_08530_));
 sg13g2_xnor2_1 _22143_ (.Y(_08531_),
    .A(_01710_),
    .B(_08530_));
 sg13g2_a21o_1 _22144_ (.A2(_08531_),
    .A1(net6776),
    .B1(net6553),
    .X(_08532_));
 sg13g2_inv_1 _22145_ (.Y(_08533_),
    .A(_01914_));
 sg13g2_xor2_1 _22146_ (.B(_08529_),
    .A(_01709_),
    .X(_08534_));
 sg13g2_o21ai_1 _22147_ (.B1(_08043_),
    .Y(_08535_),
    .A1(net6760),
    .A2(_08534_));
 sg13g2_xnor2_1 _22148_ (.Y(_08536_),
    .A(_01708_),
    .B(_08395_));
 sg13g2_o21ai_1 _22149_ (.B1(_08052_),
    .Y(_08537_),
    .A1(net6760),
    .A2(_08536_));
 sg13g2_mux2_1 _22150_ (.A0(_01556_),
    .A1(_01591_),
    .S(net7756),
    .X(_08538_));
 sg13g2_mux2_1 _22151_ (.A0(_01707_),
    .A1(net383),
    .S(_08081_),
    .X(_08539_));
 sg13g2_nor2b_1 _22152_ (.A(_01837_),
    .B_N(net383),
    .Y(_08540_));
 sg13g2_a21oi_1 _22153_ (.A1(_01837_),
    .A2(_01707_),
    .Y(_08541_),
    .B1(_08540_));
 sg13g2_nor2_1 _22154_ (.A(net7552),
    .B(_08538_),
    .Y(_08542_));
 sg13g2_nand2_2 _22155_ (.Y(_08543_),
    .A(_08122_),
    .B(_01706_));
 sg13g2_o21ai_1 _22156_ (.B1(_08543_),
    .Y(_08544_),
    .A1(net5869),
    .A2(_08541_));
 sg13g2_nor2_1 _22157_ (.A(_01705_),
    .B(net5819),
    .Y(_08545_));
 sg13g2_a21oi_1 _22158_ (.A1(net7956),
    .A2(_01706_),
    .Y(_08546_),
    .B1(_07627_));
 sg13g2_a21oi_1 _22159_ (.A1(net5810),
    .A2(_08546_),
    .Y(_08547_),
    .B1(_08545_));
 sg13g2_nor2_1 _22160_ (.A(_07711_),
    .B(_07845_),
    .Y(_08548_));
 sg13g2_nor3_1 _22161_ (.A(_07711_),
    .B(_07795_),
    .C(_07845_),
    .Y(_08549_));
 sg13g2_nand3_1 _22162_ (.B(_07768_),
    .C(_08549_),
    .A(_07756_),
    .Y(_08550_));
 sg13g2_nor2_1 _22163_ (.A(_07742_),
    .B(_08550_),
    .Y(_08551_));
 sg13g2_and2_1 _22164_ (.A(_07730_),
    .B(_08551_),
    .X(_08552_));
 sg13g2_a21oi_1 _22165_ (.A1(_07724_),
    .A2(_08552_),
    .Y(_08553_),
    .B1(_07709_));
 sg13g2_nand3_1 _22166_ (.B(_07730_),
    .C(_07741_),
    .A(_07709_),
    .Y(_08554_));
 sg13g2_or3_1 _22167_ (.A(_07723_),
    .B(_08550_),
    .C(_08554_),
    .X(_08555_));
 sg13g2_nor2b_1 _22168_ (.A(_08553_),
    .B_N(_08555_),
    .Y(_08556_));
 sg13g2_nor4_1 _22169_ (.A(_08481_),
    .B(_08498_),
    .C(_08519_),
    .D(_08542_),
    .Y(_08557_));
 sg13g2_xnor2_1 _22170_ (.Y(_08558_),
    .A(_07723_),
    .B(_08552_));
 sg13g2_xor2_1 _22171_ (.B(_08551_),
    .A(_07730_),
    .X(_08559_));
 sg13g2_xnor2_1 _22172_ (.Y(_08560_),
    .A(_07741_),
    .B(_08550_));
 sg13g2_a21o_1 _22173_ (.A2(_08549_),
    .A1(_07768_),
    .B1(_07756_),
    .X(_08561_));
 sg13g2_and2_1 _22174_ (.A(_08550_),
    .B(_08561_),
    .X(_08562_));
 sg13g2_inv_1 _22175_ (.Y(_08563_),
    .A(net7674));
 sg13g2_xor2_1 _22176_ (.B(_08549_),
    .A(_07768_),
    .X(_08564_));
 sg13g2_xnor2_1 _22177_ (.Y(_08565_),
    .A(_07795_),
    .B(_08548_));
 sg13g2_and2_1 _22178_ (.A(_01676_),
    .B(_01675_),
    .X(_08566_));
 sg13g2_nor4_1 _22179_ (.A(net6773),
    .B(_08042_),
    .C(_08046_),
    .D(_08051_),
    .Y(_08567_));
 sg13g2_a21oi_1 _22180_ (.A1(net6772),
    .A2(_08566_),
    .Y(_08568_),
    .B1(_08567_));
 sg13g2_nor2_1 _22181_ (.A(_08555_),
    .B(_08568_),
    .Y(_08569_));
 sg13g2_nor2_1 _22182_ (.A(_01677_),
    .B(net6553),
    .Y(_08570_));
 sg13g2_nor2_1 _22183_ (.A(_01678_),
    .B(net6554),
    .Y(_08571_));
 sg13g2_a21oi_1 _22184_ (.A1(net6554),
    .A2(net6553),
    .Y(_08572_),
    .B1(net6775));
 sg13g2_nor3_1 _22185_ (.A(_08570_),
    .B(_08571_),
    .C(_08572_),
    .Y(_08573_));
 sg13g2_nor2_1 _22186_ (.A(_07975_),
    .B(_07987_),
    .Y(_08574_));
 sg13g2_nand4_1 _22187_ (.B(_08007_),
    .C(_08573_),
    .A(_07997_),
    .Y(_08575_),
    .D(_08574_));
 sg13g2_nor3_1 _22188_ (.A(_08555_),
    .B(_08568_),
    .C(_08575_),
    .Y(_08576_));
 sg13g2_nor2_1 _22189_ (.A(_07952_),
    .B(_07963_),
    .Y(_08577_));
 sg13g2_and4_1 _22190_ (.A(_07932_),
    .B(_07942_),
    .C(_08576_),
    .D(_08577_),
    .X(_08578_));
 sg13g2_and2_1 _22191_ (.A(_07922_),
    .B(_08578_),
    .X(_08579_));
 sg13g2_and3_1 _22192_ (.X(_08580_),
    .A(_07893_),
    .B(_07903_),
    .C(_07913_));
 sg13g2_and4_1 _22193_ (.A(_07818_),
    .B(_07854_),
    .C(_07863_),
    .D(_07874_),
    .X(_08581_));
 sg13g2_and4_1 _22194_ (.A(_07883_),
    .B(_08579_),
    .C(_08580_),
    .D(_08581_),
    .X(_08582_));
 sg13g2_nand3_1 _22195_ (.B(_01703_),
    .C(net6775),
    .A(_01704_),
    .Y(_08583_));
 sg13g2_nand3_1 _22196_ (.B(_07706_),
    .C(_07721_),
    .A(net6760),
    .Y(_08584_));
 sg13g2_a21oi_1 _22197_ (.A1(_08583_),
    .A2(_08584_),
    .Y(_08585_),
    .B1(_08568_));
 sg13g2_nand4_1 _22198_ (.B(_08420_),
    .C(_08460_),
    .A(_08381_),
    .Y(_08586_),
    .D(_08557_));
 sg13g2_nand4_1 _22199_ (.B(_08552_),
    .C(_08573_),
    .A(_08007_),
    .Y(_08587_),
    .D(_08585_));
 sg13g2_nand2b_1 _22200_ (.Y(_08588_),
    .B(_07997_),
    .A_N(_08587_));
 sg13g2_nor4_1 _22201_ (.A(_07963_),
    .B(_07975_),
    .C(_07987_),
    .D(_08588_),
    .Y(_08589_));
 sg13g2_and2_1 _22202_ (.A(_07953_),
    .B(_08589_),
    .X(_08590_));
 sg13g2_nand3_1 _22203_ (.B(_07953_),
    .C(_08589_),
    .A(_07942_),
    .Y(_08591_));
 sg13g2_nor2b_1 _22204_ (.A(_08591_),
    .B_N(_07932_),
    .Y(_08592_));
 sg13g2_and4_1 _22205_ (.A(_07883_),
    .B(_07922_),
    .C(_08580_),
    .D(_08592_),
    .X(_08593_));
 sg13g2_nand2_1 _22206_ (.Y(_08594_),
    .A(_07874_),
    .B(_08593_));
 sg13g2_nand3_1 _22207_ (.B(_07874_),
    .C(_08593_),
    .A(_07863_),
    .Y(_08595_));
 sg13g2_nand4_1 _22208_ (.B(_07863_),
    .C(_07874_),
    .A(_07854_),
    .Y(_08596_),
    .D(_08593_));
 sg13g2_o21ai_1 _22209_ (.B1(net7672),
    .Y(_08597_),
    .A1(net7675),
    .A2(_07557_));
 sg13g2_nor2_1 _22210_ (.A(net7672),
    .B(net7675),
    .Y(_08598_));
 sg13g2_xor2_1 _22211_ (.B(_08582_),
    .A(_07803_),
    .X(_08599_));
 sg13g2_nand2_1 _22212_ (.Y(_08600_),
    .A(_09244_),
    .B(_08598_));
 sg13g2_nand3_1 _22213_ (.B(_07710_),
    .C(_08582_),
    .A(_01697_),
    .Y(_08601_));
 sg13g2_o21ai_1 _22214_ (.B1(_08601_),
    .Y(_08602_),
    .A1(_01697_),
    .A2(_07710_));
 sg13g2_a22oi_1 _22215_ (.Y(_08603_),
    .B1(_08602_),
    .B2(net6774),
    .A2(_08599_),
    .A1(_07804_));
 sg13g2_nand2_1 _22216_ (.Y(_08604_),
    .A(_07913_),
    .B(_08579_));
 sg13g2_nand3_1 _22217_ (.B(_07913_),
    .C(_08579_),
    .A(_07903_),
    .Y(_08605_));
 sg13g2_and2_1 _22218_ (.A(_08579_),
    .B(_08580_),
    .X(_08606_));
 sg13g2_xnor2_1 _22219_ (.Y(_08607_),
    .A(_07818_),
    .B(_08596_));
 sg13g2_xnor2_1 _22220_ (.Y(_08608_),
    .A(_07710_),
    .B(_07845_));
 sg13g2_xnor2_1 _22221_ (.Y(_08609_),
    .A(_07854_),
    .B(_08595_));
 sg13g2_xnor2_1 _22222_ (.Y(_08610_),
    .A(_07863_),
    .B(_08594_));
 sg13g2_nor2_1 _22223_ (.A(_08563_),
    .B(net7676),
    .Y(_08611_));
 sg13g2_xor2_1 _22224_ (.B(_08593_),
    .A(_07874_),
    .X(_08612_));
 sg13g2_xor2_1 _22225_ (.B(_08606_),
    .A(_07883_),
    .X(_08613_));
 sg13g2_and4_1 _22226_ (.A(_07946_),
    .B(_08597_),
    .C(_08600_),
    .D(_08611_),
    .X(_08614_));
 sg13g2_xnor2_1 _22227_ (.Y(_08615_),
    .A(_07893_),
    .B(_08605_));
 sg13g2_nand4_1 _22228_ (.B(_08597_),
    .C(_08600_),
    .A(_07946_),
    .Y(_08616_),
    .D(_08611_));
 sg13g2_xnor2_1 _22229_ (.Y(_08617_),
    .A(_07903_),
    .B(_08604_));
 sg13g2_nand2b_1 _22230_ (.Y(_08618_),
    .B(_01983_),
    .A_N(\load_store_unit_i.handle_misaligned_q ));
 sg13g2_xor2_1 _22231_ (.B(_08579_),
    .A(_07913_),
    .X(_08619_));
 sg13g2_xor2_1 _22232_ (.B(_08578_),
    .A(_07922_),
    .X(_08620_));
 sg13g2_xnor2_1 _22233_ (.Y(_08621_),
    .A(_07932_),
    .B(_08591_));
 sg13g2_inv_1 _22234_ (.Y(_08622_),
    .A(net7676));
 sg13g2_nor2b_1 _22235_ (.A(_01985_),
    .B_N(_01984_),
    .Y(_08623_));
 sg13g2_xor2_1 _22236_ (.B(_08590_),
    .A(_07942_),
    .X(_08624_));
 sg13g2_and2_1 _22237_ (.A(_08618_),
    .B(_08623_),
    .X(_08625_));
 sg13g2_xnor2_1 _22238_ (.Y(_08626_),
    .A(_07952_),
    .B(_08589_));
 sg13g2_nor2_1 _22239_ (.A(net7659),
    .B(_01983_),
    .Y(_08627_));
 sg13g2_xnor2_1 _22240_ (.Y(_08628_),
    .A(_07963_),
    .B(_08576_));
 sg13g2_nand2_1 _22241_ (.Y(_08629_),
    .A(_08569_),
    .B(_08573_));
 sg13g2_nand3_1 _22242_ (.B(_08569_),
    .C(_08573_),
    .A(_08007_),
    .Y(_08630_));
 sg13g2_o21ai_1 _22243_ (.B1(_07975_),
    .Y(_08631_),
    .A1(_07987_),
    .A2(_08588_));
 sg13g2_nor2b_1 _22244_ (.A(_08576_),
    .B_N(_08631_),
    .Y(_08632_));
 sg13g2_xnor2_1 _22245_ (.Y(_08633_),
    .A(_07988_),
    .B(_08588_));
 sg13g2_a22oi_1 _22246_ (.Y(_08634_),
    .B1(_08627_),
    .B2(_01985_),
    .A2(_08623_),
    .A1(_08618_));
 sg13g2_xnor2_1 _22247_ (.Y(_08635_),
    .A(_07997_),
    .B(_08630_));
 sg13g2_a21o_1 _22248_ (.A2(_08627_),
    .A1(net7657),
    .B1(_08625_),
    .X(_08636_));
 sg13g2_xnor2_1 _22249_ (.Y(_08637_),
    .A(_08007_),
    .B(_08629_));
 sg13g2_nand2_1 _22250_ (.Y(_08638_),
    .A(_08034_),
    .B(_08569_));
 sg13g2_nor2_1 _22251_ (.A(_08616_),
    .B(net7362),
    .Y(_08639_));
 sg13g2_xnor2_1 _22252_ (.Y(_08640_),
    .A(_08023_),
    .B(_08638_));
 sg13g2_nand2_1 _22253_ (.Y(_08641_),
    .A(_08614_),
    .B(_08634_));
 sg13g2_xor2_1 _22254_ (.B(_08569_),
    .A(_08034_),
    .X(_08642_));
 sg13g2_nand2b_1 _22255_ (.Y(_08643_),
    .B(_08053_),
    .A_N(_08555_));
 sg13g2_xnor2_1 _22256_ (.Y(_08644_),
    .A(_08044_),
    .B(_08643_));
 sg13g2_and3_1 _22257_ (.X(_08645_),
    .A(net7679),
    .B(_01897_),
    .C(_01886_));
 sg13g2_xnor2_1 _22258_ (.Y(_08646_),
    .A(_08053_),
    .B(_08555_));
 sg13g2_a21oi_1 _22259_ (.A1(_02033_),
    .A2(net6775),
    .Y(_08647_),
    .B1(net7455));
 sg13g2_nand2_1 _22260_ (.Y(_08648_),
    .A(net7679),
    .B(_07559_));
 sg13g2_a21oi_1 _22261_ (.A1(_01839_),
    .A2(net6761),
    .Y(_08649_),
    .B1(_01674_));
 sg13g2_nand3_1 _22262_ (.B(net7937),
    .C(_08647_),
    .A(net384),
    .Y(_08650_));
 sg13g2_a22oi_1 _22263_ (.Y(_08651_),
    .B1(_08649_),
    .B2(_08650_),
    .A2(net7937),
    .A1(net417));
 sg13g2_nand2b_1 _22264_ (.Y(_08652_),
    .B(_08649_),
    .A_N(_07006_));
 sg13g2_o21ai_1 _22265_ (.B1(net7937),
    .Y(_08653_),
    .A1(net417),
    .A2(net6761));
 sg13g2_nand2b_1 _22266_ (.Y(_08654_),
    .B(_08653_),
    .A_N(_01673_));
 sg13g2_a22oi_1 _22267_ (.Y(_08655_),
    .B1(_08652_),
    .B2(_08654_),
    .A2(_08647_),
    .A1(net384));
 sg13g2_inv_1 _22268_ (.Y(_08656_),
    .A(_08655_));
 sg13g2_nor2_1 _22269_ (.A(net7482),
    .B(_08242_),
    .Y(_08657_));
 sg13g2_and2_1 _22270_ (.A(_06767_),
    .B(net7289),
    .X(_08658_));
 sg13g2_nand2_1 _22271_ (.Y(_08659_),
    .A(_06767_),
    .B(net7289));
 sg13g2_nand2_1 _22272_ (.Y(_08660_),
    .A(_00540_),
    .B(_08658_));
 sg13g2_nor2_1 _22273_ (.A(net7482),
    .B(net7370),
    .Y(_08661_));
 sg13g2_nand2_1 _22274_ (.Y(_08662_),
    .A(net7923),
    .B(net7383));
 sg13g2_nor2_1 _22275_ (.A(_06768_),
    .B(_08662_),
    .Y(_08663_));
 sg13g2_nand2_1 _22276_ (.Y(_08664_),
    .A(_01672_),
    .B(net6818));
 sg13g2_nand3_1 _22277_ (.B(_07608_),
    .C(_08645_),
    .A(_08622_),
    .Y(_08665_));
 sg13g2_nor2_1 _22278_ (.A(_02104_),
    .B(net7127),
    .Y(_08666_));
 sg13g2_nor4_1 _22279_ (.A(_01891_),
    .B(_07701_),
    .C(_07872_),
    .D(_07884_),
    .Y(_08667_));
 sg13g2_a21oi_1 _22280_ (.A1(net469),
    .A2(net7123),
    .Y(_08668_),
    .B1(_08666_));
 sg13g2_nand4_1 _22281_ (.B(_07780_),
    .C(_07870_),
    .A(net7929),
    .Y(_08669_),
    .D(_07881_));
 sg13g2_o21ai_1 _22282_ (.B1(_08664_),
    .Y(_08670_),
    .A1(net6818),
    .A2(_08668_));
 sg13g2_nand2_1 _22283_ (.Y(_08671_),
    .A(_01671_),
    .B(net6815));
 sg13g2_nor2_1 _22284_ (.A(net7271),
    .B(net7128),
    .Y(_08672_));
 sg13g2_nor2_1 _22285_ (.A(_07555_),
    .B(net7608),
    .Y(_08673_));
 sg13g2_a21oi_1 _22286_ (.A1(net468),
    .A2(net7124),
    .Y(_08674_),
    .B1(_08672_));
 sg13g2_o21ai_1 _22287_ (.B1(_08671_),
    .Y(_08675_),
    .A1(net6817),
    .A2(_08674_));
 sg13g2_nand2_1 _22288_ (.Y(_08676_),
    .A(_01670_),
    .B(net6814));
 sg13g2_nor2_1 _22289_ (.A(_15462_),
    .B(net7125),
    .Y(_08677_));
 sg13g2_a21oi_1 _22290_ (.A1(net6627),
    .A2(net7122),
    .Y(_08678_),
    .B1(_08677_));
 sg13g2_o21ai_1 _22291_ (.B1(_08676_),
    .Y(_08679_),
    .A1(net6814),
    .A2(_08678_));
 sg13g2_nand2_1 _22292_ (.Y(_08680_),
    .A(_01669_),
    .B(net6820));
 sg13g2_o21ai_1 _22293_ (.B1(_08645_),
    .Y(_08681_),
    .A1(_08667_),
    .A2(_08673_));
 sg13g2_nor2_1 _22294_ (.A(_14725_),
    .B(net7125),
    .Y(_08682_));
 sg13g2_a21oi_1 _22295_ (.A1(net6628),
    .A2(net7122),
    .Y(_08683_),
    .B1(_08682_));
 sg13g2_o21ai_1 _22296_ (.B1(_08680_),
    .Y(_08684_),
    .A1(net6820),
    .A2(_08683_));
 sg13g2_nand2_1 _22297_ (.Y(_08685_),
    .A(_05174_),
    .B(_00005_));
 sg13g2_nor3_1 _22298_ (.A(net7993),
    .B(net7427),
    .C(_08685_),
    .Y(_08686_));
 sg13g2_nor2_1 _22299_ (.A(_03628_),
    .B(_04792_),
    .Y(_08687_));
 sg13g2_nand2_1 _22300_ (.Y(_08688_),
    .A(_03629_),
    .B(_04791_));
 sg13g2_nor3_1 _22301_ (.A(net7482),
    .B(net7926),
    .C(_08242_),
    .Y(_08689_));
 sg13g2_nand2_1 _22302_ (.Y(_08690_),
    .A(net7477),
    .B(_08657_));
 sg13g2_nand3_1 _22303_ (.B(_08688_),
    .C(_08689_),
    .A(net7129),
    .Y(_08691_));
 sg13g2_o21ai_1 _22304_ (.B1(_08691_),
    .Y(_08692_),
    .A1(net7129),
    .A2(_08688_));
 sg13g2_a22oi_1 _22305_ (.Y(_08693_),
    .B1(_08692_),
    .B2(_05213_),
    .A2(_08690_),
    .A1(_08687_));
 sg13g2_nor2_1 _22306_ (.A(net7926),
    .B(_08662_),
    .Y(_08694_));
 sg13g2_nand2_1 _22307_ (.Y(_08695_),
    .A(net7477),
    .B(_08661_));
 sg13g2_nand3_1 _22308_ (.B(net7609),
    .C(_08598_),
    .A(_07559_),
    .Y(_08696_));
 sg13g2_nor2b_1 _22309_ (.A(net7924),
    .B_N(net7674),
    .Y(_08697_));
 sg13g2_a21oi_1 _22310_ (.A1(net7993),
    .A2(_08693_),
    .Y(_08698_),
    .B1(_08686_));
 sg13g2_nand2b_1 _22311_ (.Y(_08699_),
    .B(net7923),
    .A_N(_08698_));
 sg13g2_nand3_1 _22312_ (.B(_06767_),
    .C(_08699_),
    .A(net7385),
    .Y(_08700_));
 sg13g2_nand3_1 _22313_ (.B(_06767_),
    .C(_08699_),
    .A(net7381),
    .Y(_08701_));
 sg13g2_nor2b_1 _22314_ (.A(net8016),
    .B_N(_00004_),
    .Y(_08702_));
 sg13g2_nor2_1 _22315_ (.A(_00537_),
    .B(_00536_),
    .Y(_08703_));
 sg13g2_nand4_1 _22316_ (.B(net7609),
    .C(_08598_),
    .A(net7610),
    .Y(_08704_),
    .D(_08697_));
 sg13g2_o21ai_1 _22317_ (.B1(_08702_),
    .Y(_08705_),
    .A1(_03816_),
    .A2(_08703_));
 sg13g2_nor2_1 _22318_ (.A(net7924),
    .B(_08242_),
    .Y(_08706_));
 sg13g2_and2_1 _22319_ (.A(_08705_),
    .B(_08706_),
    .X(_08707_));
 sg13g2_nor2_1 _22320_ (.A(net7924),
    .B(net7370),
    .Y(_08708_));
 sg13g2_and2_1 _22321_ (.A(_08705_),
    .B(_08708_),
    .X(_08709_));
 sg13g2_a22oi_1 _22322_ (.Y(_08710_),
    .B1(net7083),
    .B2(_00104_),
    .A2(net7096),
    .A1(net7629));
 sg13g2_inv_1 _22323_ (.Y(_08711_),
    .A(_01909_));
 sg13g2_nand2_1 _22324_ (.Y(_08712_),
    .A(_01668_),
    .B(net6805));
 sg13g2_o21ai_1 _22325_ (.B1(_08712_),
    .Y(_08713_),
    .A1(net6805),
    .A2(_08710_));
 sg13g2_nand3_1 _22326_ (.B(net7285),
    .C(_08705_),
    .A(_00103_),
    .Y(_08714_));
 sg13g2_and2_1 _22327_ (.A(_08665_),
    .B(_08704_),
    .X(_08715_));
 sg13g2_nand2_1 _22328_ (.Y(_08716_),
    .A(net7923),
    .B(net7977));
 sg13g2_nor2_1 _22329_ (.A(_05162_),
    .B(_08716_),
    .Y(_08717_));
 sg13g2_a221oi_1 _22330_ (.B2(net6568),
    .C1(net6808),
    .B1(_08717_),
    .A1(net7629),
    .Y(_08718_),
    .A2(_08689_));
 sg13g2_a22oi_1 _22331_ (.Y(_08719_),
    .B1(_08714_),
    .B2(_08718_),
    .A2(net6807),
    .A1(_02055_));
 sg13g2_nand2_1 _22332_ (.Y(_08720_),
    .A(net7977),
    .B(net6808));
 sg13g2_a21oi_1 _22333_ (.A1(_07792_),
    .A2(net7385),
    .Y(_08721_),
    .B1(_08703_));
 sg13g2_o21ai_1 _22334_ (.B1(_03816_),
    .Y(_08722_),
    .A1(_00537_),
    .A2(_00536_));
 sg13g2_nor2_1 _22335_ (.A(net7922),
    .B(_08722_),
    .Y(_08723_));
 sg13g2_nand3_1 _22336_ (.B(net6568),
    .C(net7092),
    .A(net7977),
    .Y(_08724_));
 sg13g2_nor2_1 _22337_ (.A(_05199_),
    .B(_05201_),
    .Y(_08725_));
 sg13g2_nand2_1 _22338_ (.Y(_08726_),
    .A(_01631_),
    .B(net6568));
 sg13g2_nor2_1 _22339_ (.A(_01631_),
    .B(net6568),
    .Y(_08727_));
 sg13g2_o21ai_1 _22340_ (.B1(_08726_),
    .Y(_08728_),
    .A1(net7977),
    .A2(_08727_));
 sg13g2_nand2b_1 _22341_ (.Y(_08729_),
    .B(_00535_),
    .A_N(net6474));
 sg13g2_nand2_1 _22342_ (.Y(_08730_),
    .A(net8020),
    .B(_00531_));
 sg13g2_nor2_1 _22343_ (.A(_08729_),
    .B(_08730_),
    .Y(_08731_));
 sg13g2_a21oi_1 _22344_ (.A1(_08725_),
    .A2(_08731_),
    .Y(_08732_),
    .B1(_00600_));
 sg13g2_o21ai_1 _22345_ (.B1(_08724_),
    .Y(_08733_),
    .A1(net7092),
    .A2(_08732_));
 sg13g2_nand2_1 _22346_ (.Y(_08734_),
    .A(net8010),
    .B(_08733_));
 sg13g2_mux2_1 _22347_ (.A0(net6569),
    .A1(_01665_),
    .S(net6470),
    .X(_08735_));
 sg13g2_a21oi_1 _22348_ (.A1(_03628_),
    .A2(net7098),
    .Y(_08736_),
    .B1(net8012));
 sg13g2_a221oi_1 _22349_ (.B2(net7990),
    .C1(_08736_),
    .B1(_08735_),
    .A1(net7995),
    .Y(_08737_),
    .A2(net6568));
 sg13g2_a21oi_1 _22350_ (.A1(_08734_),
    .A2(_08737_),
    .Y(_08738_),
    .B1(net7482));
 sg13g2_and2_1 _22351_ (.A(net7482),
    .B(_08705_),
    .X(_08739_));
 sg13g2_a221oi_1 _22352_ (.B2(_00102_),
    .C1(_08738_),
    .B1(_08739_),
    .A1(net5970),
    .Y(_08740_),
    .A2(_08723_));
 sg13g2_o21ai_1 _22353_ (.B1(_08720_),
    .Y(_08741_),
    .A1(net6808),
    .A2(_08740_));
 sg13g2_and2_1 _22354_ (.A(_08706_),
    .B(_08721_),
    .X(_08742_));
 sg13g2_nand2b_1 _22355_ (.Y(_08743_),
    .B(_00532_),
    .A_N(_00531_));
 sg13g2_nor2_1 _22356_ (.A(_08729_),
    .B(_08743_),
    .Y(_08744_));
 sg13g2_nor2_1 _22357_ (.A(_08694_),
    .B(_08735_),
    .Y(_08745_));
 sg13g2_a21oi_1 _22358_ (.A1(net7431),
    .A2(_08744_),
    .Y(_08746_),
    .B1(_00599_));
 sg13g2_a21oi_1 _22359_ (.A1(_08694_),
    .A2(_08746_),
    .Y(_08747_),
    .B1(_08745_));
 sg13g2_mux2_1 _22360_ (.A0(net6571),
    .A1(_01664_),
    .S(net6472),
    .X(_08748_));
 sg13g2_nand2_1 _22361_ (.Y(_08749_),
    .A(net7328),
    .B(net7092));
 sg13g2_a22oi_1 _22362_ (.Y(_08750_),
    .B1(_08748_),
    .B2(net7987),
    .A2(net6569),
    .A1(net7996));
 sg13g2_a22oi_1 _22363_ (.Y(_08751_),
    .B1(_08749_),
    .B2(net7629),
    .A2(_08747_),
    .A1(net8010));
 sg13g2_a21oi_1 _22364_ (.A1(_08750_),
    .A2(_08751_),
    .Y(_08752_),
    .B1(_08662_));
 sg13g2_and2_1 _22365_ (.A(_08708_),
    .B(_08721_),
    .X(_08753_));
 sg13g2_a221oi_1 _22366_ (.B2(net6057),
    .C1(_08752_),
    .B1(net7080),
    .A1(net5923),
    .Y(_08754_),
    .A2(net7083));
 sg13g2_nand2_1 _22367_ (.Y(_08755_),
    .A(_01665_),
    .B(net6805));
 sg13g2_o21ai_1 _22368_ (.B1(_08755_),
    .Y(_08756_),
    .A1(net6805),
    .A2(_08754_));
 sg13g2_nand2_1 _22369_ (.Y(_08757_),
    .A(_00099_),
    .B(_08739_));
 sg13g2_inv_1 _22370_ (.Y(_08758_),
    .A(_08759_));
 sg13g2_nand2b_1 _22371_ (.Y(_08759_),
    .B(net8021),
    .A_N(net8019));
 sg13g2_nor2_1 _22372_ (.A(_08729_),
    .B(_08759_),
    .Y(_08760_));
 sg13g2_a21oi_1 _22373_ (.A1(net7431),
    .A2(_08760_),
    .Y(_08761_),
    .B1(_00597_));
 sg13g2_nor2_1 _22374_ (.A(net7095),
    .B(_08761_),
    .Y(_08762_));
 sg13g2_a21oi_1 _22375_ (.A1(net7095),
    .A2(_08748_),
    .Y(_08763_),
    .B1(_08762_));
 sg13g2_mux2_1 _22376_ (.A0(net6572),
    .A1(_01663_),
    .S(net6471),
    .X(_08764_));
 sg13g2_a21oi_1 _22377_ (.A1(net7329),
    .A2(net7099),
    .Y(_08765_),
    .B1(net8012));
 sg13g2_a221oi_1 _22378_ (.B2(net7990),
    .C1(_08765_),
    .B1(_08764_),
    .A1(net7995),
    .Y(_08766_),
    .A2(net6571));
 sg13g2_o21ai_1 _22379_ (.B1(_08766_),
    .Y(_08767_),
    .A1(net7631),
    .A2(_08763_));
 sg13g2_a22oi_1 _22380_ (.Y(_08768_),
    .B1(_08767_),
    .B2(net7922),
    .A2(_08723_),
    .A1(net6058));
 sg13g2_a21oi_1 _22381_ (.A1(_08757_),
    .A2(_08768_),
    .Y(_08769_),
    .B1(net6807));
 sg13g2_a21o_1 _22382_ (.A2(net6807),
    .A1(_01664_),
    .B1(_08769_),
    .X(_08770_));
 sg13g2_nand2_1 _22383_ (.Y(_08771_),
    .A(_01663_),
    .B(net6807));
 sg13g2_nor2_1 _22384_ (.A(net8020),
    .B(_00531_),
    .Y(_08772_));
 sg13g2_or2_1 _22385_ (.X(_08773_),
    .B(net8022),
    .A(net8020));
 sg13g2_nor2_1 _22386_ (.A(_08729_),
    .B(_08773_),
    .Y(_08774_));
 sg13g2_nor2_1 _22387_ (.A(_08694_),
    .B(_08764_),
    .Y(_08775_));
 sg13g2_a21oi_1 _22388_ (.A1(net7431),
    .A2(_08774_),
    .Y(_08776_),
    .B1(_00596_));
 sg13g2_a21oi_1 _22389_ (.A1(_08681_),
    .A2(_08715_),
    .Y(_08777_),
    .B1(_08636_));
 sg13g2_a21oi_1 _22390_ (.A1(net7097),
    .A2(_08776_),
    .Y(_08778_),
    .B1(_08775_));
 sg13g2_nand2_1 _22391_ (.Y(_08779_),
    .A(net8009),
    .B(_08778_));
 sg13g2_mux2_1 _22392_ (.A0(net6575),
    .A1(_01662_),
    .S(net6472),
    .X(_08780_));
 sg13g2_a21o_1 _22393_ (.A2(_08715_),
    .A1(_08681_),
    .B1(net7360),
    .X(_08781_));
 sg13g2_a21oi_1 _22394_ (.A1(net7331),
    .A2(net7098),
    .Y(_08782_),
    .B1(net8012));
 sg13g2_a221oi_1 _22395_ (.B2(net7987),
    .C1(_08782_),
    .B1(_08780_),
    .A1(net7996),
    .Y(_08783_),
    .A2(net6572));
 sg13g2_or4_1 _22396_ (.A(_07555_),
    .B(_07562_),
    .C(_07570_),
    .D(net7608),
    .X(_08784_));
 sg13g2_and2_1 _22397_ (.A(_08634_),
    .B(_08784_),
    .X(_08785_));
 sg13g2_a21oi_1 _22398_ (.A1(_08779_),
    .A2(_08783_),
    .Y(_08786_),
    .B1(_08662_));
 sg13g2_a221oi_1 _22399_ (.B2(net6397),
    .C1(_08786_),
    .B1(net7080),
    .A1(_00098_),
    .Y(_08787_),
    .A2(net7083));
 sg13g2_o21ai_1 _22400_ (.B1(_08771_),
    .Y(_08788_),
    .A1(net6806),
    .A2(_08787_));
 sg13g2_nand2_1 _22401_ (.Y(_08789_),
    .A(_01662_),
    .B(net6807));
 sg13g2_nor2_1 _22402_ (.A(_05199_),
    .B(net8018),
    .Y(_08790_));
 sg13g2_nand2_1 _22403_ (.Y(_08791_),
    .A(_00534_),
    .B(_05201_));
 sg13g2_nor2_1 _22404_ (.A(_08694_),
    .B(_08780_),
    .Y(_08792_));
 sg13g2_a21oi_1 _22405_ (.A1(_08731_),
    .A2(_08790_),
    .Y(_08793_),
    .B1(_00595_));
 sg13g2_a21oi_1 _22406_ (.A1(net7097),
    .A2(_08793_),
    .Y(_08794_),
    .B1(_08792_));
 sg13g2_nand2_1 _22407_ (.Y(_08795_),
    .A(net8009),
    .B(_08794_));
 sg13g2_mux2_1 _22408_ (.A0(net6576),
    .A1(_01661_),
    .S(net6470),
    .X(_08796_));
 sg13g2_nand3_1 _22409_ (.B(_08665_),
    .C(_08784_),
    .A(_08634_),
    .Y(_08797_));
 sg13g2_a21oi_1 _22410_ (.A1(_03367_),
    .A2(net7098),
    .Y(_08798_),
    .B1(net8012));
 sg13g2_a221oi_1 _22411_ (.B2(net7987),
    .C1(_08798_),
    .B1(_08796_),
    .A1(net7996),
    .Y(_08799_),
    .A2(net6575));
 sg13g2_nor2_1 _22412_ (.A(_08777_),
    .B(_08797_),
    .Y(_08800_));
 sg13g2_a21oi_1 _22413_ (.A1(_08795_),
    .A2(_08799_),
    .Y(_08801_),
    .B1(net7285));
 sg13g2_a221oi_1 _22414_ (.B2(net6398),
    .C1(_08801_),
    .B1(net7080),
    .A1(_00097_),
    .Y(_08802_),
    .A2(net7083));
 sg13g2_o21ai_1 _22415_ (.B1(_08789_),
    .Y(_08803_),
    .A1(net6806),
    .A2(_08802_));
 sg13g2_a21o_1 _22416_ (.A2(_07555_),
    .A1(_08622_),
    .B1(net7608),
    .X(_08804_));
 sg13g2_nor2_1 _22417_ (.A(net7097),
    .B(_08796_),
    .Y(_08805_));
 sg13g2_a21oi_1 _22418_ (.A1(_08744_),
    .A2(_08790_),
    .Y(_08806_),
    .B1(_00594_));
 sg13g2_a21oi_1 _22419_ (.A1(net7097),
    .A2(_08806_),
    .Y(_08807_),
    .B1(_08805_));
 sg13g2_a21oi_1 _22420_ (.A1(_08669_),
    .A2(_08804_),
    .Y(_08808_),
    .B1(_08648_));
 sg13g2_mux2_1 _22421_ (.A0(net6579),
    .A1(_01659_),
    .S(net6470),
    .X(_08809_));
 sg13g2_nand2_1 _22422_ (.Y(_08810_),
    .A(net7332),
    .B(net7092));
 sg13g2_a22oi_1 _22423_ (.Y(_08811_),
    .B1(_08809_),
    .B2(net7991),
    .A2(net6576),
    .A1(net7997));
 sg13g2_a22oi_1 _22424_ (.Y(_08812_),
    .B1(_08810_),
    .B2(net7629),
    .A2(_08807_),
    .A1(net8009));
 sg13g2_a21oi_1 _22425_ (.A1(_08811_),
    .A2(_08812_),
    .Y(_08813_),
    .B1(_08662_));
 sg13g2_a221oi_1 _22426_ (.B2(net6399),
    .C1(_08813_),
    .B1(net7080),
    .A1(net5924),
    .Y(_08814_),
    .A2(_08709_));
 sg13g2_nand2_1 _22427_ (.Y(_08815_),
    .A(_01661_),
    .B(net6804));
 sg13g2_o21ai_1 _22428_ (.B1(_08815_),
    .Y(_08816_),
    .A1(net6804),
    .A2(_08814_));
 sg13g2_nand2_1 _22429_ (.Y(_08817_),
    .A(_01660_),
    .B(net6814));
 sg13g2_nor2_1 _22430_ (.A(net7074),
    .B(net7125),
    .Y(_08818_));
 sg13g2_nand2b_1 _22431_ (.Y(_08819_),
    .B(_08634_),
    .A_N(_08808_));
 sg13g2_a21oi_1 _22432_ (.A1(net6636),
    .A2(net7122),
    .Y(_08820_),
    .B1(_08818_));
 sg13g2_o21ai_1 _22433_ (.B1(_08817_),
    .Y(_08821_),
    .A1(net6823),
    .A2(_08820_));
 sg13g2_nor2_1 _22434_ (.A(net7096),
    .B(_08809_),
    .Y(_08822_));
 sg13g2_a21oi_1 _22435_ (.A1(_08760_),
    .A2(_08790_),
    .Y(_08823_),
    .B1(_00593_));
 sg13g2_a21oi_1 _22436_ (.A1(net7096),
    .A2(_08823_),
    .Y(_08824_),
    .B1(_08822_));
 sg13g2_nand2_1 _22437_ (.Y(_08825_),
    .A(net8009),
    .B(_08824_));
 sg13g2_nor3_1 _22438_ (.A(_09041_),
    .B(_08797_),
    .C(_08808_),
    .Y(_08826_));
 sg13g2_mux2_1 _22439_ (.A0(net6582),
    .A1(_01658_),
    .S(net6473),
    .X(_08827_));
 sg13g2_a21oi_1 _22440_ (.A1(net7333),
    .A2(net7098),
    .Y(_08828_),
    .B1(net8012));
 sg13g2_a221oi_1 _22441_ (.B2(net7987),
    .C1(_08828_),
    .B1(_08827_),
    .A1(net7996),
    .Y(_08829_),
    .A2(net6579));
 sg13g2_a21oi_1 _22442_ (.A1(_08825_),
    .A2(_08829_),
    .Y(_08830_),
    .B1(net7285));
 sg13g2_a221oi_1 _22443_ (.B2(net6400),
    .C1(_08830_),
    .B1(net7080),
    .A1(_00095_),
    .Y(_08831_),
    .A2(net7083));
 sg13g2_nand2_1 _22444_ (.Y(_08832_),
    .A(_01659_),
    .B(net6806));
 sg13g2_o21ai_1 _22445_ (.B1(_08832_),
    .Y(_08833_),
    .A1(net6806),
    .A2(_08831_));
 sg13g2_nor2_1 _22446_ (.A(net7097),
    .B(_08827_),
    .Y(_08834_));
 sg13g2_a21oi_1 _22447_ (.A1(_08774_),
    .A2(_08790_),
    .Y(_08835_),
    .B1(_00592_));
 sg13g2_a21oi_1 _22448_ (.A1(_08681_),
    .A2(_08704_),
    .Y(_08836_),
    .B1(_08797_));
 sg13g2_a21oi_1 _22449_ (.A1(net7097),
    .A2(_08835_),
    .Y(_08837_),
    .B1(_08834_));
 sg13g2_a21o_1 _22450_ (.A2(_08704_),
    .A1(_08681_),
    .B1(_08797_),
    .X(_08838_));
 sg13g2_mux2_1 _22451_ (.A0(net6603),
    .A1(_01657_),
    .S(net6473),
    .X(_08839_));
 sg13g2_nor3_1 _22452_ (.A(_08510_),
    .B(net7360),
    .C(_08808_),
    .Y(_08840_));
 sg13g2_nand2_1 _22453_ (.Y(_08841_),
    .A(net7334),
    .B(_08695_));
 sg13g2_a22oi_1 _22454_ (.Y(_08842_),
    .B1(_08839_),
    .B2(net7991),
    .A2(net6582),
    .A1(net7997));
 sg13g2_a22oi_1 _22455_ (.Y(_08843_),
    .B1(_08841_),
    .B2(net7629),
    .A2(_08837_),
    .A1(net8009));
 sg13g2_a21oi_1 _22456_ (.A1(_08842_),
    .A2(_08843_),
    .Y(_08844_),
    .B1(_08662_));
 sg13g2_a22oi_1 _22457_ (.Y(_08845_),
    .B1(_08836_),
    .B2(_08840_),
    .A2(_08826_),
    .A1(_08781_));
 sg13g2_a221oi_1 _22458_ (.B2(net6478),
    .C1(_08844_),
    .B1(net7080),
    .A1(_00094_),
    .Y(_08846_),
    .A2(_08709_));
 sg13g2_nand2_1 _22459_ (.Y(_08847_),
    .A(_01658_),
    .B(net6804));
 sg13g2_o21ai_1 _22460_ (.B1(_08847_),
    .Y(_08848_),
    .A1(net6804),
    .A2(_08846_));
 sg13g2_nand2_1 _22461_ (.Y(_08849_),
    .A(net7978),
    .B(net6807));
 sg13g2_nor2_1 _22462_ (.A(_00534_),
    .B(_05201_),
    .Y(_08850_));
 sg13g2_nor2_1 _22463_ (.A(_08614_),
    .B(net7362),
    .Y(_08851_));
 sg13g2_a21oi_1 _22464_ (.A1(_08731_),
    .A2(net7430),
    .Y(_08852_),
    .B1(_00591_));
 sg13g2_nor2_1 _22465_ (.A(net7094),
    .B(_08852_),
    .Y(_08853_));
 sg13g2_a21oi_1 _22466_ (.A1(net7095),
    .A2(_08839_),
    .Y(_08854_),
    .B1(_08853_));
 sg13g2_nand2b_1 _22467_ (.Y(_08855_),
    .B(_08851_),
    .A_N(_08845_));
 sg13g2_mux2_1 _22468_ (.A0(net6605),
    .A1(_01656_),
    .S(net6470),
    .X(_08856_));
 sg13g2_a21oi_1 _22469_ (.A1(net7336),
    .A2(net7098),
    .Y(_08857_),
    .B1(net8012));
 sg13g2_a221oi_1 _22470_ (.B2(net7987),
    .C1(_08857_),
    .B1(_08856_),
    .A1(net7996),
    .Y(_08858_),
    .A2(net6603));
 sg13g2_o21ai_1 _22471_ (.B1(_08858_),
    .Y(_08859_),
    .A1(_05180_),
    .A2(_08854_));
 sg13g2_and2_1 _22472_ (.A(net6557),
    .B(_08723_),
    .X(_08860_));
 sg13g2_a221oi_1 _22473_ (.B2(net7922),
    .C1(_08860_),
    .B1(_08859_),
    .A1(_00093_),
    .Y(_08861_),
    .A2(_08739_));
 sg13g2_o21ai_1 _22474_ (.B1(_08849_),
    .Y(_08862_),
    .A1(net6807),
    .A2(_08861_));
 sg13g2_nand2_1 _22475_ (.Y(_08863_),
    .A(_00092_),
    .B(net7084));
 sg13g2_a21oi_1 _22476_ (.A1(_08744_),
    .A2(net7430),
    .Y(_08864_),
    .B1(_00590_));
 sg13g2_nor2_1 _22477_ (.A(net7095),
    .B(_08864_),
    .Y(_08865_));
 sg13g2_a21oi_1 _22478_ (.A1(net7092),
    .A2(_08856_),
    .Y(_08866_),
    .B1(_08865_));
 sg13g2_mux2_1 _22479_ (.A0(net6584),
    .A1(net7979),
    .S(net6470),
    .X(_08867_));
 sg13g2_a21oi_1 _22480_ (.A1(net7338),
    .A2(net7099),
    .Y(_08868_),
    .B1(net8015));
 sg13g2_a221oi_1 _22481_ (.B2(net7991),
    .C1(_08868_),
    .B1(_08867_),
    .A1(net7997),
    .Y(_08869_),
    .A2(net6605));
 sg13g2_o21ai_1 _22482_ (.B1(_08869_),
    .Y(_08870_),
    .A1(_05180_),
    .A2(_08866_));
 sg13g2_nand2_1 _22483_ (.Y(_08871_),
    .A(net6479),
    .B(net7082));
 sg13g2_a221oi_1 _22484_ (.B2(net7289),
    .C1(net6812),
    .B1(_08870_),
    .A1(net6479),
    .Y(_08872_),
    .A2(_08742_));
 sg13g2_o21ai_1 _22485_ (.B1(_08855_),
    .Y(_08873_),
    .A1(_08641_),
    .A2(net7103));
 sg13g2_inv_1 _22486_ (.Y(_08874_),
    .A(net6977));
 sg13g2_a22oi_1 _22487_ (.Y(_08875_),
    .B1(_08863_),
    .B2(_08872_),
    .A2(net6812),
    .A1(_02081_));
 sg13g2_nor2_1 _22488_ (.A(net7096),
    .B(_08867_),
    .Y(_08876_));
 sg13g2_a21oi_1 _22489_ (.A1(_08760_),
    .A2(net7430),
    .Y(_08877_),
    .B1(_00589_));
 sg13g2_a21oi_1 _22490_ (.A1(net7096),
    .A2(_08877_),
    .Y(_08878_),
    .B1(_08876_));
 sg13g2_nand2_1 _22491_ (.Y(_08879_),
    .A(net8009),
    .B(_08878_));
 sg13g2_mux2_1 _22492_ (.A0(net6586),
    .A1(net7980),
    .S(net6470),
    .X(_08880_));
 sg13g2_a21oi_1 _22493_ (.A1(net7340),
    .A2(net7099),
    .Y(_08881_),
    .B1(net8015));
 sg13g2_a221oi_1 _22494_ (.B2(net7991),
    .C1(_08881_),
    .B1(_08880_),
    .A1(net7997),
    .Y(_08882_),
    .A2(net6584));
 sg13g2_a21oi_1 _22495_ (.A1(_08879_),
    .A2(_08882_),
    .Y(_08883_),
    .B1(net7285));
 sg13g2_a221oi_1 _22496_ (.B2(_00107_),
    .C1(_08883_),
    .B1(net7080),
    .A1(_00091_),
    .Y(_08884_),
    .A2(net7083));
 sg13g2_nand2_1 _22497_ (.Y(_08885_),
    .A(_01655_),
    .B(net6806));
 sg13g2_o21ai_1 _22498_ (.B1(_08885_),
    .Y(_08886_),
    .A1(net6806),
    .A2(_08884_));
 sg13g2_nor2_1 _22499_ (.A(net7097),
    .B(_08880_),
    .Y(_08887_));
 sg13g2_a21oi_1 _22500_ (.A1(_08774_),
    .A2(_08850_),
    .Y(_08888_),
    .B1(_00588_));
 sg13g2_nor2b_1 _22501_ (.A(net7806),
    .B_N(_01895_),
    .Y(_08889_));
 sg13g2_a21oi_1 _22502_ (.A1(net7096),
    .A2(_08888_),
    .Y(_08890_),
    .B1(_08887_));
 sg13g2_nand2_1 _22503_ (.Y(_08891_),
    .A(net8009),
    .B(_08890_));
 sg13g2_nand2b_1 _22504_ (.Y(_08892_),
    .B(net7808),
    .A_N(_01896_));
 sg13g2_mux2_1 _22505_ (.A0(net6607),
    .A1(_01653_),
    .S(net6470),
    .X(_08893_));
 sg13g2_inv_1 _22506_ (.Y(_08894_),
    .A(_01903_));
 sg13g2_a21oi_1 _22507_ (.A1(net7341),
    .A2(net7099),
    .Y(_08895_),
    .B1(net8015));
 sg13g2_a221oi_1 _22508_ (.B2(net7987),
    .C1(_08895_),
    .B1(_08893_),
    .A1(net7996),
    .Y(_08896_),
    .A2(net6586));
 sg13g2_a21oi_1 _22509_ (.A1(_08891_),
    .A2(_08896_),
    .Y(_08897_),
    .B1(net7285));
 sg13g2_a221oi_1 _22510_ (.B2(net6620),
    .C1(_08897_),
    .B1(_08753_),
    .A1(net5954),
    .Y(_08898_),
    .A2(_08709_));
 sg13g2_nand2_1 _22511_ (.Y(_08899_),
    .A(net7980),
    .B(net6804));
 sg13g2_o21ai_1 _22512_ (.B1(_08899_),
    .Y(_08900_),
    .A1(net6804),
    .A2(_08898_));
 sg13g2_nor2_1 _22513_ (.A(_00534_),
    .B(_00533_),
    .Y(_08901_));
 sg13g2_nand2_1 _22514_ (.Y(_08902_),
    .A(_05199_),
    .B(_05201_));
 sg13g2_nor2_1 _22515_ (.A(net7096),
    .B(_08893_),
    .Y(_08903_));
 sg13g2_a21oi_1 _22516_ (.A1(_08731_),
    .A2(_08901_),
    .Y(_08904_),
    .B1(_00586_));
 sg13g2_a21oi_1 _22517_ (.A1(net7096),
    .A2(_08904_),
    .Y(_08905_),
    .B1(_08903_));
 sg13g2_nand2_1 _22518_ (.Y(_08906_),
    .A(net8009),
    .B(_08905_));
 sg13g2_mux2_1 _22519_ (.A0(net6608),
    .A1(_01652_),
    .S(net6470),
    .X(_08907_));
 sg13g2_a21oi_1 _22520_ (.A1(_02818_),
    .A2(net7098),
    .Y(_08908_),
    .B1(net8012));
 sg13g2_a221oi_1 _22521_ (.B2(net7987),
    .C1(_08908_),
    .B1(_08907_),
    .A1(net7995),
    .Y(_08909_),
    .A2(net6607));
 sg13g2_a21oi_1 _22522_ (.A1(_08906_),
    .A2(_08909_),
    .Y(_08910_),
    .B1(net7285));
 sg13g2_a221oi_1 _22523_ (.B2(net6635),
    .C1(_08910_),
    .B1(net7080),
    .A1(net5955),
    .Y(_08911_),
    .A2(net7083));
 sg13g2_nand2_1 _22524_ (.Y(_08912_),
    .A(_01653_),
    .B(net6805));
 sg13g2_o21ai_1 _22525_ (.B1(_08912_),
    .Y(_08913_),
    .A1(net6805),
    .A2(_08911_));
 sg13g2_nand2_1 _22526_ (.Y(_08914_),
    .A(net5969),
    .B(_08739_));
 sg13g2_a21oi_1 _22527_ (.A1(_08744_),
    .A2(_08901_),
    .Y(_08915_),
    .B1(_00585_));
 sg13g2_nor2_1 _22528_ (.A(net7094),
    .B(_08915_),
    .Y(_08916_));
 sg13g2_a21oi_1 _22529_ (.A1(net7091),
    .A2(_08907_),
    .Y(_08917_),
    .B1(_08916_));
 sg13g2_mux2_1 _22530_ (.A0(net6609),
    .A1(_01651_),
    .S(net6471),
    .X(_08918_));
 sg13g2_a21oi_1 _22531_ (.A1(net7343),
    .A2(net7099),
    .Y(_08919_),
    .B1(net8015));
 sg13g2_a221oi_1 _22532_ (.B2(net7990),
    .C1(_08919_),
    .B1(_08918_),
    .A1(net7995),
    .Y(_08920_),
    .A2(net6608));
 sg13g2_o21ai_1 _22533_ (.B1(_08920_),
    .Y(_08921_),
    .A1(net7631),
    .A2(_08917_));
 sg13g2_a22oi_1 _22534_ (.Y(_08922_),
    .B1(_08921_),
    .B2(net7922),
    .A2(_08723_),
    .A1(_00100_));
 sg13g2_mux4_1 _22535_ (.S0(net7906),
    .A0(_00922_),
    .A1(_00957_),
    .A2(_00992_),
    .A3(_01028_),
    .S1(net7827),
    .X(_08923_));
 sg13g2_a21oi_1 _22536_ (.A1(_08914_),
    .A2(_08922_),
    .Y(_08924_),
    .B1(net6808));
 sg13g2_a21o_1 _22537_ (.A2(net6807),
    .A1(_01652_),
    .B1(_08924_),
    .X(_08925_));
 sg13g2_nand2_1 _22538_ (.Y(_08926_),
    .A(_00086_),
    .B(net7084));
 sg13g2_a21oi_1 _22539_ (.A1(_08760_),
    .A2(_08901_),
    .Y(_08927_),
    .B1(_00584_));
 sg13g2_nor2_1 _22540_ (.A(net7094),
    .B(_08927_),
    .Y(_08928_));
 sg13g2_a21oi_1 _22541_ (.A1(net7091),
    .A2(_08918_),
    .Y(_08929_),
    .B1(_08928_));
 sg13g2_mux2_1 _22542_ (.A0(net6611),
    .A1(_01650_),
    .S(net6471),
    .X(_08930_));
 sg13g2_a21oi_1 _22543_ (.A1(net7344),
    .A2(net7098),
    .Y(_08931_),
    .B1(net8013));
 sg13g2_a221oi_1 _22544_ (.B2(net7990),
    .C1(_08931_),
    .B1(_08930_),
    .A1(net7995),
    .Y(_08932_),
    .A2(net6609));
 sg13g2_o21ai_1 _22545_ (.B1(_08932_),
    .Y(_08933_),
    .A1(net7631),
    .A2(_08929_));
 sg13g2_a221oi_1 _22546_ (.B2(net7290),
    .C1(net6812),
    .B1(_08933_),
    .A1(_00089_),
    .Y(_08934_),
    .A2(net7081));
 sg13g2_a22oi_1 _22547_ (.Y(_08935_),
    .B1(_08926_),
    .B2(_08934_),
    .A2(net6808),
    .A1(_02089_));
 sg13g2_nor2_1 _22548_ (.A(_08694_),
    .B(_08930_),
    .Y(_08936_));
 sg13g2_nand2_1 _22549_ (.Y(_08937_),
    .A(_05201_),
    .B(_08772_));
 sg13g2_nand2_1 _22550_ (.Y(_08938_),
    .A(_08772_),
    .B(_08901_));
 sg13g2_nor2_1 _22551_ (.A(_08729_),
    .B(_08938_),
    .Y(_08939_));
 sg13g2_nor3_1 _22552_ (.A(_00583_),
    .B(_08695_),
    .C(_08939_),
    .Y(_08940_));
 sg13g2_nor2_1 _22553_ (.A(_08936_),
    .B(_08940_),
    .Y(_08941_));
 sg13g2_mux2_1 _22554_ (.A0(net6612),
    .A1(_01648_),
    .S(net6472),
    .X(_08942_));
 sg13g2_nand2_1 _22555_ (.Y(_08943_),
    .A(net7993),
    .B(net6611));
 sg13g2_o21ai_1 _22556_ (.B1(net7629),
    .Y(_08944_),
    .A1(_02616_),
    .A2(_08689_));
 sg13g2_nand3_1 _22557_ (.B(_08943_),
    .C(_08944_),
    .A(net7922),
    .Y(_08945_));
 sg13g2_inv_1 _22558_ (.Y(_08946_),
    .A(net7693));
 sg13g2_a221oi_1 _22559_ (.B2(net7990),
    .C1(_08945_),
    .B1(_08942_),
    .A1(net8010),
    .Y(_08947_),
    .A2(_08941_));
 sg13g2_a221oi_1 _22560_ (.B2(_00078_),
    .C1(net7922),
    .B1(_08721_),
    .A1(_00085_),
    .Y(_08948_),
    .A2(_08705_));
 sg13g2_nor4_1 _22561_ (.A(net7370),
    .B(_08701_),
    .C(_08947_),
    .D(_08948_),
    .Y(_08949_));
 sg13g2_a21o_1 _22562_ (.A2(_08701_),
    .A1(_01650_),
    .B1(_08949_),
    .X(_08950_));
 sg13g2_nand2_1 _22563_ (.Y(_08951_),
    .A(_01649_),
    .B(net6821));
 sg13g2_nor2_1 _22564_ (.A(_12791_),
    .B(net7129),
    .Y(_08952_));
 sg13g2_a21oi_1 _22565_ (.A1(net6638),
    .A2(net7121),
    .Y(_08953_),
    .B1(_08952_));
 sg13g2_o21ai_1 _22566_ (.B1(_08951_),
    .Y(_08954_),
    .A1(net6821),
    .A2(_08953_));
 sg13g2_nor2_1 _22567_ (.A(_02098_),
    .B(_08722_),
    .Y(_08955_));
 sg13g2_a21o_1 _22568_ (.A2(_08705_),
    .A1(_00084_),
    .B1(_08955_),
    .X(_08956_));
 sg13g2_nor3_1 _22569_ (.A(_00535_),
    .B(net6474),
    .C(_08730_),
    .Y(_08957_));
 sg13g2_mux4_1 _22570_ (.S0(net7906),
    .A0(_00788_),
    .A1(_00820_),
    .A2(_00852_),
    .A3(_00887_),
    .S1(net7827),
    .X(_08958_));
 sg13g2_a21oi_1 _22571_ (.A1(net7431),
    .A2(_08957_),
    .Y(_08959_),
    .B1(_00582_));
 sg13g2_nor2_1 _22572_ (.A(net7095),
    .B(_08959_),
    .Y(_08960_));
 sg13g2_a21oi_1 _22573_ (.A1(net7092),
    .A2(_08942_),
    .Y(_08961_),
    .B1(_08960_));
 sg13g2_mux2_1 _22574_ (.A0(net6614),
    .A1(_01647_),
    .S(net6469),
    .X(_08962_));
 sg13g2_a21oi_1 _22575_ (.A1(_02549_),
    .A2(net7100),
    .Y(_08963_),
    .B1(net8014));
 sg13g2_a221oi_1 _22576_ (.B2(net7989),
    .C1(_08963_),
    .B1(_08962_),
    .A1(net7994),
    .Y(_08964_),
    .A2(net6612));
 sg13g2_o21ai_1 _22577_ (.B1(_08964_),
    .Y(_08965_),
    .A1(_05180_),
    .A2(_08961_));
 sg13g2_a221oi_1 _22578_ (.B2(net7290),
    .C1(net6812),
    .B1(_08965_),
    .A1(_08706_),
    .Y(_08966_),
    .A2(net5933));
 sg13g2_mux2_1 _22579_ (.A0(_08923_),
    .A1(_08958_),
    .S(net7486),
    .X(_08967_));
 sg13g2_a21oi_1 _22580_ (.A1(_02098_),
    .A2(net6812),
    .Y(_08968_),
    .B1(_08966_));
 sg13g2_or2_1 _22581_ (.X(_08969_),
    .B(net7081),
    .A(net6812));
 sg13g2_nand2_1 _22582_ (.Y(_08970_),
    .A(_01647_),
    .B(_08969_));
 sg13g2_nand2_1 _22583_ (.Y(_08971_),
    .A(_00083_),
    .B(net7087));
 sg13g2_nor3_1 _22584_ (.A(_00535_),
    .B(net6474),
    .C(_08743_),
    .Y(_08972_));
 sg13g2_nor2_1 _22585_ (.A(net7806),
    .B(_01895_),
    .Y(_08973_));
 sg13g2_or2_1 _22586_ (.X(_08974_),
    .B(_01895_),
    .A(net7806));
 sg13g2_a21oi_1 _22587_ (.A1(net7431),
    .A2(_08972_),
    .Y(_08975_),
    .B1(_00581_));
 sg13g2_nor2_1 _22588_ (.A(net7094),
    .B(_08975_),
    .Y(_08976_));
 sg13g2_a21oi_1 _22589_ (.A1(net7090),
    .A2(_08962_),
    .Y(_08977_),
    .B1(_08976_));
 sg13g2_mux2_1 _22590_ (.A0(net6599),
    .A1(_01646_),
    .S(net6469),
    .X(_08978_));
 sg13g2_a21oi_1 _22591_ (.A1(net7347),
    .A2(net7101),
    .Y(_08979_),
    .B1(net8011));
 sg13g2_a221oi_1 _22592_ (.B2(net7988),
    .C1(_08979_),
    .B1(_08978_),
    .A1(net7992),
    .Y(_08980_),
    .A2(net6614));
 sg13g2_o21ai_1 _22593_ (.B1(_08980_),
    .Y(_08981_),
    .A1(net7630),
    .A2(_08977_));
 sg13g2_a22oi_1 _22594_ (.Y(_08982_),
    .B1(_08981_),
    .B2(net7287),
    .A2(net7086),
    .A1(net6057));
 sg13g2_mux2_1 _22595_ (.A0(_01214_),
    .A1(_01566_),
    .S(net7837),
    .X(_08983_));
 sg13g2_o21ai_1 _22596_ (.B1(_08970_),
    .Y(_08984_),
    .A1(net6809),
    .A2(_08982_));
 sg13g2_nand2_1 _22597_ (.Y(_08985_),
    .A(_01646_),
    .B(_08969_));
 sg13g2_nor3_1 _22598_ (.A(_00535_),
    .B(net6473),
    .C(_08759_),
    .Y(_08986_));
 sg13g2_a21oi_1 _22599_ (.A1(net7431),
    .A2(_08986_),
    .Y(_08987_),
    .B1(_00580_));
 sg13g2_nor2b_1 _22600_ (.A(net7835),
    .B_N(net7895),
    .Y(_08988_));
 sg13g2_nor2_1 _22601_ (.A(net7094),
    .B(_08987_),
    .Y(_08989_));
 sg13g2_a21oi_1 _22602_ (.A1(net7090),
    .A2(_08978_),
    .Y(_08990_),
    .B1(_08989_));
 sg13g2_mux2_1 _22603_ (.A0(net6602),
    .A1(_01645_),
    .S(_08728_),
    .X(_08991_));
 sg13g2_a21oi_1 _22604_ (.A1(_02439_),
    .A2(net7101),
    .Y(_08992_),
    .B1(net8011));
 sg13g2_a221oi_1 _22605_ (.B2(net7988),
    .C1(_08992_),
    .B1(_08991_),
    .A1(net7992),
    .Y(_08993_),
    .A2(net6599));
 sg13g2_o21ai_1 _22606_ (.B1(_08993_),
    .Y(_08994_),
    .A1(net7630),
    .A2(_08990_));
 sg13g2_a22oi_1 _22607_ (.Y(_08995_),
    .B1(_08994_),
    .B2(net7290),
    .A2(net7089),
    .A1(net6058));
 sg13g2_o21ai_1 _22608_ (.B1(_08985_),
    .Y(_08996_),
    .A1(net6811),
    .A2(_08995_));
 sg13g2_nand2_1 _22609_ (.Y(_08997_),
    .A(_01645_),
    .B(net6759));
 sg13g2_a221oi_1 _22610_ (.B2(_00862_),
    .C1(net7810),
    .B1(_08988_),
    .A1(net7820),
    .Y(_08998_),
    .A2(_08983_));
 sg13g2_nor3_1 _22611_ (.A(_00535_),
    .B(net6473),
    .C(_08773_),
    .Y(_08999_));
 sg13g2_a21oi_1 _22612_ (.A1(net7431),
    .A2(_08999_),
    .Y(_09000_),
    .B1(_00579_));
 sg13g2_and2_1 _22613_ (.A(net7815),
    .B(net7835),
    .X(_09001_));
 sg13g2_nor2_1 _22614_ (.A(net7093),
    .B(_09000_),
    .Y(_09002_));
 sg13g2_a21oi_1 _22615_ (.A1(net7090),
    .A2(_08991_),
    .Y(_09003_),
    .B1(_09002_));
 sg13g2_nand2_1 _22616_ (.Y(_09004_),
    .A(net7816),
    .B(net7835));
 sg13g2_mux2_1 _22617_ (.A0(net6621),
    .A1(_01644_),
    .S(_08728_),
    .X(_09005_));
 sg13g2_a21oi_1 _22618_ (.A1(_02361_),
    .A2(net7101),
    .Y(_09006_),
    .B1(net8011));
 sg13g2_a221oi_1 _22619_ (.B2(net7989),
    .C1(_09006_),
    .B1(_09005_),
    .A1(net7994),
    .Y(_09007_),
    .A2(net6602));
 sg13g2_o21ai_1 _22620_ (.B1(_09007_),
    .Y(_09008_),
    .A1(net7630),
    .A2(_09003_));
 sg13g2_a22oi_1 _22621_ (.Y(_09009_),
    .B1(_09008_),
    .B2(net7286),
    .A2(net7085),
    .A1(net6397));
 sg13g2_o21ai_1 _22622_ (.B1(_08997_),
    .Y(_09010_),
    .A1(net6809),
    .A2(_09009_));
 sg13g2_inv_1 _22623_ (.Y(_09011_),
    .A(net7735));
 sg13g2_nand2_1 _22624_ (.Y(_09012_),
    .A(_01644_),
    .B(net6759));
 sg13g2_a21oi_1 _22625_ (.A1(_08790_),
    .A2(_08957_),
    .Y(_09013_),
    .B1(_00578_));
 sg13g2_nor2_1 _22626_ (.A(net7093),
    .B(_09013_),
    .Y(_09014_));
 sg13g2_a21oi_1 _22627_ (.A1(net7090),
    .A2(_09005_),
    .Y(_09015_),
    .B1(_09014_));
 sg13g2_mux2_1 _22628_ (.A0(net6623),
    .A1(_01643_),
    .S(_08728_),
    .X(_09016_));
 sg13g2_a21oi_1 _22629_ (.A1(_02283_),
    .A2(_08690_),
    .Y(_09017_),
    .B1(net8014));
 sg13g2_a221oi_1 _22630_ (.B2(net7989),
    .C1(_09017_),
    .B1(_09016_),
    .A1(net7994),
    .Y(_09018_),
    .A2(net6621));
 sg13g2_o21ai_1 _22631_ (.B1(_09018_),
    .Y(_09019_),
    .A1(net7630),
    .A2(_09015_));
 sg13g2_mux2_1 _22632_ (.A0(_00724_),
    .A1(_00756_),
    .S(net7837),
    .X(_09020_));
 sg13g2_a22oi_1 _22633_ (.Y(_09021_),
    .B1(_09019_),
    .B2(net7286),
    .A2(net7085),
    .A1(net6398));
 sg13g2_o21ai_1 _22634_ (.B1(_09012_),
    .Y(_09022_),
    .A1(net6810),
    .A2(_09021_));
 sg13g2_nor2_1 _22635_ (.A(net7522),
    .B(_09020_),
    .Y(_09023_));
 sg13g2_a221oi_1 _22636_ (.B2(_01643_),
    .C1(net7922),
    .B1(_08721_),
    .A1(_00079_),
    .Y(_09024_),
    .A2(_08705_));
 sg13g2_nor2_1 _22637_ (.A(_08694_),
    .B(_09016_),
    .Y(_09025_));
 sg13g2_nor2b_1 _22638_ (.A(net7835),
    .B_N(net7816),
    .Y(_09026_));
 sg13g2_a21oi_1 _22639_ (.A1(_08790_),
    .A2(_08972_),
    .Y(_09027_),
    .B1(_00577_));
 sg13g2_nand2b_1 _22640_ (.Y(_09028_),
    .B(net7816),
    .A_N(net7832));
 sg13g2_a21oi_1 _22641_ (.A1(_08694_),
    .A2(_09027_),
    .Y(_09029_),
    .B1(_09025_));
 sg13g2_mux2_1 _22642_ (.A0(net6625),
    .A1(_01642_),
    .S(net6469),
    .X(_09030_));
 sg13g2_nand2_1 _22643_ (.Y(_09031_),
    .A(net7993),
    .B(net6623));
 sg13g2_o21ai_1 _22644_ (.B1(net7629),
    .Y(_09032_),
    .A1(_02205_),
    .A2(_08689_));
 sg13g2_nand3_1 _22645_ (.B(_09031_),
    .C(_09032_),
    .A(net7922),
    .Y(_09033_));
 sg13g2_a221oi_1 _22646_ (.B2(net7989),
    .C1(_09033_),
    .B1(_09030_),
    .A1(net8010),
    .Y(_09034_),
    .A2(_09029_));
 sg13g2_nor3_1 _22647_ (.A(_08700_),
    .B(_09024_),
    .C(_09034_),
    .Y(_09035_));
 sg13g2_a21o_1 _22648_ (.A2(_08700_),
    .A1(_01643_),
    .B1(_09035_),
    .X(_09036_));
 sg13g2_nand2_1 _22649_ (.Y(_09037_),
    .A(_01642_),
    .B(net6759));
 sg13g2_a21oi_1 _22650_ (.A1(_08790_),
    .A2(_08986_),
    .Y(_09038_),
    .B1(_00607_));
 sg13g2_nor2_1 _22651_ (.A(net7094),
    .B(_09038_),
    .Y(_09039_));
 sg13g2_a21oi_1 _22652_ (.A1(net7091),
    .A2(_09030_),
    .Y(_09040_),
    .B1(_09039_));
 sg13g2_inv_1 _22653_ (.Y(_09041_),
    .A(_01898_));
 sg13g2_mux2_1 _22654_ (.A0(net6626),
    .A1(_01641_),
    .S(_08728_),
    .X(_09042_));
 sg13g2_a21oi_1 _22655_ (.A1(net7349),
    .A2(net7101),
    .Y(_09043_),
    .B1(net8011));
 sg13g2_mux2_1 _22656_ (.A0(_00660_),
    .A1(_00692_),
    .S(net7837),
    .X(_09044_));
 sg13g2_a221oi_1 _22657_ (.B2(net7989),
    .C1(_09043_),
    .B1(_09042_),
    .A1(net7994),
    .Y(_09045_),
    .A2(net6625));
 sg13g2_o21ai_1 _22658_ (.B1(_09045_),
    .Y(_09046_),
    .A1(net7630),
    .A2(_09040_));
 sg13g2_a22oi_1 _22659_ (.Y(_09047_),
    .B1(_09046_),
    .B2(net7286),
    .A2(net7085),
    .A1(net6400));
 sg13g2_o21ai_1 _22660_ (.B1(_09037_),
    .Y(_09048_),
    .A1(net6810),
    .A2(_09047_));
 sg13g2_nand2_1 _22661_ (.Y(_09049_),
    .A(_01641_),
    .B(net6759));
 sg13g2_a21oi_1 _22662_ (.A1(_08790_),
    .A2(_08999_),
    .Y(_09050_),
    .B1(_00606_));
 sg13g2_nor2_1 _22663_ (.A(net7093),
    .B(_09050_),
    .Y(_09051_));
 sg13g2_a21oi_1 _22664_ (.A1(net7091),
    .A2(_09042_),
    .Y(_09052_),
    .B1(_09051_));
 sg13g2_mux2_1 _22665_ (.A0(net6627),
    .A1(_01640_),
    .S(net6469),
    .X(_09053_));
 sg13g2_a21oi_1 _22666_ (.A1(_02067_),
    .A2(net7100),
    .Y(_09054_),
    .B1(net8013));
 sg13g2_a221oi_1 _22667_ (.B2(net7988),
    .C1(_09054_),
    .B1(_09053_),
    .A1(net7992),
    .Y(_09055_),
    .A2(net6626));
 sg13g2_o21ai_1 _22668_ (.B1(_09055_),
    .Y(_09056_),
    .A1(net7631),
    .A2(_09052_));
 sg13g2_a22oi_1 _22669_ (.Y(_09057_),
    .B1(_09056_),
    .B2(net7287),
    .A2(net7086),
    .A1(net6478));
 sg13g2_o21ai_1 _22670_ (.B1(_09049_),
    .Y(_09058_),
    .A1(net6810),
    .A2(_09057_));
 sg13g2_nand2_1 _22671_ (.Y(_09059_),
    .A(_01640_),
    .B(_08969_));
 sg13g2_o21ai_1 _22672_ (.B1(_08973_),
    .Y(_09060_),
    .A1(net7506),
    .A2(_09044_));
 sg13g2_a21oi_1 _22673_ (.A1(net7430),
    .A2(_08957_),
    .Y(_09061_),
    .B1(_00605_));
 sg13g2_nor2_1 _22674_ (.A(net7093),
    .B(_09061_),
    .Y(_09062_));
 sg13g2_a21oi_1 _22675_ (.A1(net7091),
    .A2(_09053_),
    .Y(_09063_),
    .B1(_09062_));
 sg13g2_mux2_1 _22676_ (.A0(net6628),
    .A1(_01639_),
    .S(net6469),
    .X(_09064_));
 sg13g2_or3_1 _22677_ (.A(_08998_),
    .B(_09023_),
    .C(_09060_),
    .X(_09065_));
 sg13g2_a21oi_1 _22678_ (.A1(_15563_),
    .A2(net7100),
    .Y(_09066_),
    .B1(net8013));
 sg13g2_a221oi_1 _22679_ (.B2(net7988),
    .C1(_09066_),
    .B1(_09064_),
    .A1(net7992),
    .Y(_09067_),
    .A2(net6627));
 sg13g2_o21ai_1 _22680_ (.B1(_09067_),
    .Y(_09068_),
    .A1(net7631),
    .A2(_09063_));
 sg13g2_a22oi_1 _22681_ (.Y(_09069_),
    .B1(_09068_),
    .B2(net7290),
    .A2(net7089),
    .A1(net6557));
 sg13g2_nor2b_1 _22682_ (.A(net7808),
    .B_N(net7806),
    .Y(_09070_));
 sg13g2_o21ai_1 _22683_ (.B1(_09059_),
    .Y(_09071_),
    .A1(net6811),
    .A2(_09069_));
 sg13g2_nand2_1 _22684_ (.Y(_09072_),
    .A(_01639_),
    .B(_08969_));
 sg13g2_nand2b_1 _22685_ (.Y(_09073_),
    .B(net7806),
    .A_N(net7808));
 sg13g2_a21oi_1 _22686_ (.A1(net7430),
    .A2(_08972_),
    .Y(_09074_),
    .B1(_00604_));
 sg13g2_nor2_1 _22687_ (.A(net7093),
    .B(_09074_),
    .Y(_09075_));
 sg13g2_a21oi_1 _22688_ (.A1(net7091),
    .A2(_09064_),
    .Y(_09076_),
    .B1(_09075_));
 sg13g2_mux2_1 _22689_ (.A0(net6636),
    .A1(_01637_),
    .S(net6469),
    .X(_09077_));
 sg13g2_a21oi_1 _22690_ (.A1(net7273),
    .A2(net7101),
    .Y(_09078_),
    .B1(net8011));
 sg13g2_a221oi_1 _22691_ (.B2(net7988),
    .C1(_09078_),
    .B1(_09077_),
    .A1(net7992),
    .Y(_09079_),
    .A2(net6628));
 sg13g2_o21ai_1 _22692_ (.B1(_09079_),
    .Y(_09080_),
    .A1(net7631),
    .A2(_09076_));
 sg13g2_a22oi_1 _22693_ (.Y(_09081_),
    .B1(_09080_),
    .B2(net7290),
    .A2(net7089),
    .A1(net6479));
 sg13g2_o21ai_1 _22694_ (.B1(_09072_),
    .Y(_09082_),
    .A1(net6811),
    .A2(_09081_));
 sg13g2_nand2_1 _22695_ (.Y(_09083_),
    .A(_01638_),
    .B(net6818));
 sg13g2_nor2b_1 _22696_ (.A(net7127),
    .B_N(_11665_),
    .Y(_09084_));
 sg13g2_a21oi_1 _22697_ (.A1(net6639),
    .A2(net7123),
    .Y(_09085_),
    .B1(_09084_));
 sg13g2_o21ai_1 _22698_ (.B1(_09083_),
    .Y(_09086_),
    .A1(net6818),
    .A2(_09085_));
 sg13g2_nand2_1 _22699_ (.Y(_09087_),
    .A(_01637_),
    .B(_08969_));
 sg13g2_a21oi_1 _22700_ (.A1(net7430),
    .A2(_08986_),
    .Y(_09088_),
    .B1(_00603_));
 sg13g2_nor2_1 _22701_ (.A(net7093),
    .B(_09088_),
    .Y(_09089_));
 sg13g2_a21oi_1 _22702_ (.A1(net7091),
    .A2(_09077_),
    .Y(_09090_),
    .B1(_09089_));
 sg13g2_mux2_1 _22703_ (.A0(net6638),
    .A1(_01636_),
    .S(net6469),
    .X(_09091_));
 sg13g2_a21oi_1 _22704_ (.A1(net7275),
    .A2(net7100),
    .Y(_09092_),
    .B1(net8011));
 sg13g2_a221oi_1 _22705_ (.B2(net7988),
    .C1(_09092_),
    .B1(_09091_),
    .A1(net7992),
    .Y(_09093_),
    .A2(net6636));
 sg13g2_o21ai_1 _22706_ (.B1(_09093_),
    .Y(_09094_),
    .A1(net7631),
    .A2(_09090_));
 sg13g2_a22oi_1 _22707_ (.Y(_09095_),
    .B1(_09094_),
    .B2(net7290),
    .A2(net7089),
    .A1(_00107_));
 sg13g2_o21ai_1 _22708_ (.B1(_09087_),
    .Y(_09096_),
    .A1(net6811),
    .A2(_09095_));
 sg13g2_nand2_1 _22709_ (.Y(_09097_),
    .A(_01636_),
    .B(_08969_));
 sg13g2_a21oi_1 _22710_ (.A1(net7430),
    .A2(_08999_),
    .Y(_09098_),
    .B1(_00602_));
 sg13g2_nor2_1 _22711_ (.A(net7093),
    .B(_09098_),
    .Y(_09099_));
 sg13g2_a21oi_1 _22712_ (.A1(net7090),
    .A2(_09091_),
    .Y(_09100_),
    .B1(_09099_));
 sg13g2_mux2_1 _22713_ (.A0(net6639),
    .A1(_01635_),
    .S(_08728_),
    .X(_09101_));
 sg13g2_mux4_1 _22714_ (.S0(net7899),
    .A0(_01204_),
    .A1(_01239_),
    .A2(_01274_),
    .A3(_01309_),
    .S1(net7819),
    .X(_09102_));
 sg13g2_a21oi_1 _22715_ (.A1(_13358_),
    .A2(net7101),
    .Y(_09103_),
    .B1(net8011));
 sg13g2_a221oi_1 _22716_ (.B2(net7988),
    .C1(_09103_),
    .B1(_09101_),
    .A1(net7992),
    .Y(_09104_),
    .A2(net6638));
 sg13g2_o21ai_1 _22717_ (.B1(_09104_),
    .Y(_09105_),
    .A1(net7630),
    .A2(_09100_));
 sg13g2_a22oi_1 _22718_ (.Y(_09106_),
    .B1(_09105_),
    .B2(net7287),
    .A2(net7086),
    .A1(net6620));
 sg13g2_o21ai_1 _22719_ (.B1(_09097_),
    .Y(_09107_),
    .A1(net6809),
    .A2(_09106_));
 sg13g2_nand2_1 _22720_ (.Y(_09108_),
    .A(_01635_),
    .B(net6759));
 sg13g2_a21oi_1 _22721_ (.A1(_08901_),
    .A2(_08957_),
    .Y(_09109_),
    .B1(_00601_));
 sg13g2_nor2_1 _22722_ (.A(net7094),
    .B(_09109_),
    .Y(_09110_));
 sg13g2_a21oi_1 _22723_ (.A1(net7090),
    .A2(_09101_),
    .Y(_09111_),
    .B1(_09110_));
 sg13g2_mux2_1 _22724_ (.A0(net6640),
    .A1(_01634_),
    .S(_08728_),
    .X(_09112_));
 sg13g2_a21oi_1 _22725_ (.A1(net7282),
    .A2(net7101),
    .Y(_09113_),
    .B1(net8011));
 sg13g2_a221oi_1 _22726_ (.B2(net7988),
    .C1(_09113_),
    .B1(_09112_),
    .A1(net7992),
    .Y(_09114_),
    .A2(net6639));
 sg13g2_o21ai_1 _22727_ (.B1(_09114_),
    .Y(_09115_),
    .A1(net7630),
    .A2(_09111_));
 sg13g2_a22oi_1 _22728_ (.Y(_09116_),
    .B1(_09115_),
    .B2(net7287),
    .A2(net7086),
    .A1(net6635));
 sg13g2_o21ai_1 _22729_ (.B1(_09108_),
    .Y(_09117_),
    .A1(net6809),
    .A2(_09116_));
 sg13g2_nand2_1 _22730_ (.Y(_09118_),
    .A(_01634_),
    .B(_08969_));
 sg13g2_a21oi_1 _22731_ (.A1(_08901_),
    .A2(_08972_),
    .Y(_09119_),
    .B1(_00598_));
 sg13g2_nor2_1 _22732_ (.A(net7093),
    .B(_09119_),
    .Y(_09120_));
 sg13g2_a21oi_1 _22733_ (.A1(net7090),
    .A2(_09112_),
    .Y(_09121_),
    .B1(_09120_));
 sg13g2_mux2_1 _22734_ (.A0(net6717),
    .A1(_01633_),
    .S(net6472),
    .X(_09122_));
 sg13g2_a21oi_1 _22735_ (.A1(net7283),
    .A2(_08690_),
    .Y(_09123_),
    .B1(net8014));
 sg13g2_a221oi_1 _22736_ (.B2(net7989),
    .C1(_09123_),
    .B1(_09122_),
    .A1(net7994),
    .Y(_09124_),
    .A2(net6640));
 sg13g2_o21ai_1 _22737_ (.B1(_09124_),
    .Y(_09125_),
    .A1(net7630),
    .A2(_09121_));
 sg13g2_a22oi_1 _22738_ (.Y(_09126_),
    .B1(_09125_),
    .B2(net7287),
    .A2(net7086),
    .A1(_00100_));
 sg13g2_o21ai_1 _22739_ (.B1(_09118_),
    .Y(_09127_),
    .A1(net6810),
    .A2(_09126_));
 sg13g2_nand2_1 _22740_ (.Y(_09128_),
    .A(_01633_),
    .B(net6759));
 sg13g2_or4_1 _22741_ (.A(_00535_),
    .B(net6473),
    .C(_08759_),
    .D(_08902_),
    .X(_09129_));
 sg13g2_nor2b_1 _22742_ (.A(_00587_),
    .B_N(_09129_),
    .Y(_09130_));
 sg13g2_nor2_1 _22743_ (.A(net7095),
    .B(_09130_),
    .Y(_09131_));
 sg13g2_a21oi_1 _22744_ (.A1(net7092),
    .A2(_09122_),
    .Y(_09132_),
    .B1(_09131_));
 sg13g2_nand2_1 _22745_ (.Y(_09133_),
    .A(_01632_),
    .B(net6472));
 sg13g2_o21ai_1 _22746_ (.B1(_09133_),
    .Y(_09134_),
    .A1(net6735),
    .A2(net6472));
 sg13g2_a21oi_1 _22747_ (.A1(net7076),
    .A2(_08690_),
    .Y(_09135_),
    .B1(net8014));
 sg13g2_a221oi_1 _22748_ (.B2(net7989),
    .C1(_09135_),
    .B1(_09134_),
    .A1(net7994),
    .Y(_09136_),
    .A2(net6717));
 sg13g2_o21ai_1 _22749_ (.B1(_09136_),
    .Y(_09137_),
    .A1(_05180_),
    .A2(_09132_));
 sg13g2_mux4_1 _22750_ (.S0(net7899),
    .A0(_01063_),
    .A1(_01098_),
    .A2(_01133_),
    .A3(_01168_),
    .S1(net7819),
    .X(_09138_));
 sg13g2_a22oi_1 _22751_ (.Y(_09139_),
    .B1(_09137_),
    .B2(net7286),
    .A2(net7085),
    .A1(_00089_));
 sg13g2_nand2_1 _22752_ (.Y(_09140_),
    .A(_00089_),
    .B(_08709_));
 sg13g2_o21ai_1 _22753_ (.B1(_09128_),
    .Y(_09141_),
    .A1(net6809),
    .A2(_09139_));
 sg13g2_nand2_1 _22754_ (.Y(_09142_),
    .A(_01632_),
    .B(net6759));
 sg13g2_nand2b_1 _22755_ (.Y(_09143_),
    .B(_08695_),
    .A_N(_09134_));
 sg13g2_nor3_1 _22756_ (.A(_00535_),
    .B(net6473),
    .C(_08938_),
    .Y(_09144_));
 sg13g2_or3_1 _22757_ (.A(_00576_),
    .B(_08695_),
    .C(_09144_),
    .X(_09145_));
 sg13g2_nand3_1 _22758_ (.B(_09143_),
    .C(_09145_),
    .A(net8010),
    .Y(_09146_));
 sg13g2_mux2_1 _22759_ (.A0(_09102_),
    .A1(_09138_),
    .S(net7486),
    .X(_09147_));
 sg13g2_mux2_1 _22760_ (.A0(_00575_),
    .A1(_00545_),
    .S(net8021),
    .X(_09148_));
 sg13g2_a221oi_1 _22761_ (.B2(net8020),
    .C1(_08791_),
    .B1(_09148_),
    .A1(_00574_),
    .Y(_09149_),
    .A2(_08758_));
 sg13g2_and2_1 _22762_ (.A(_01896_),
    .B(_01895_),
    .X(_09150_));
 sg13g2_a21oi_1 _22763_ (.A1(_05199_),
    .A2(_08937_),
    .Y(_09151_),
    .B1(_09149_));
 sg13g2_nand2_1 _22764_ (.Y(_09152_),
    .A(_01896_),
    .B(net7808));
 sg13g2_inv_1 _22765_ (.Y(_09153_),
    .A(net7813));
 sg13g2_mux4_1 _22766_ (.S0(net8021),
    .A0(_00546_),
    .A1(_00547_),
    .A2(_00548_),
    .A3(_00549_),
    .S1(net8019),
    .X(_09154_));
 sg13g2_o21ai_1 _22767_ (.B1(_09151_),
    .Y(_09155_),
    .A1(_05201_),
    .A2(_09154_));
 sg13g2_o21ai_1 _22768_ (.B1(net8017),
    .Y(_09156_),
    .A1(_00550_),
    .A2(_08938_));
 sg13g2_o21ai_1 _22769_ (.B1(_09156_),
    .Y(_09157_),
    .A1(net8017),
    .A2(_09155_));
 sg13g2_nand3b_1 _22770_ (.B(net8018),
    .C(_08772_),
    .Y(_09158_),
    .A_N(_00569_));
 sg13g2_nand2b_1 _22771_ (.Y(_09159_),
    .B(net8021),
    .A_N(_00566_));
 sg13g2_o21ai_1 _22772_ (.B1(_09159_),
    .Y(_09160_),
    .A1(_00555_),
    .A2(net8021));
 sg13g2_a22oi_1 _22773_ (.Y(_09161_),
    .B1(_09160_),
    .B2(net8019),
    .A2(_08758_),
    .A1(_05159_));
 sg13g2_o21ai_1 _22774_ (.B1(_09158_),
    .Y(_09162_),
    .A1(net8018),
    .A2(_09161_));
 sg13g2_nand2b_1 _22775_ (.Y(_09163_),
    .B(net8019),
    .A_N(_00572_));
 sg13g2_o21ai_1 _22776_ (.B1(_09163_),
    .Y(_09164_),
    .A1(_00570_),
    .A2(net8019));
 sg13g2_o21ai_1 _22777_ (.B1(net8018),
    .Y(_09165_),
    .A1(_00571_),
    .A2(_08743_));
 sg13g2_a21o_1 _22778_ (.A2(_09164_),
    .A1(net8022),
    .B1(_09165_),
    .X(_09166_));
 sg13g2_o21ai_1 _22779_ (.B1(_09166_),
    .Y(_09167_),
    .A1(net8018),
    .A2(_08772_));
 sg13g2_nor2_1 _22780_ (.A(_05199_),
    .B(_08937_),
    .Y(_09168_));
 sg13g2_a22oi_1 _22781_ (.Y(_09169_),
    .B1(_09168_),
    .B2(_00573_),
    .A2(_09167_),
    .A1(_05199_));
 sg13g2_nor2_1 _22782_ (.A(_09162_),
    .B(_09169_),
    .Y(_09170_));
 sg13g2_o21ai_1 _22783_ (.B1(_00543_),
    .Y(_09171_),
    .A1(_09157_),
    .A2(_09170_));
 sg13g2_nor2_1 _22784_ (.A(_00559_),
    .B(_05199_),
    .Y(_09172_));
 sg13g2_o21ai_1 _22785_ (.B1(net8017),
    .Y(_09173_),
    .A1(_08937_),
    .A2(_09172_));
 sg13g2_mux4_1 _22786_ (.S0(net8020),
    .A0(_00568_),
    .A1(_00565_),
    .A2(_00564_),
    .A3(_00567_),
    .S1(net8021),
    .X(_09174_));
 sg13g2_or3_1 _22787_ (.A(net8017),
    .B(_08938_),
    .C(_09174_),
    .X(_09175_));
 sg13g2_mux4_1 _22788_ (.S0(_00532_),
    .A0(_00563_),
    .A1(_00561_),
    .A2(_00560_),
    .A3(_00562_),
    .S1(net8022),
    .X(_09176_));
 sg13g2_nand2_1 _22789_ (.Y(_09177_),
    .A(net8018),
    .B(_08773_));
 sg13g2_nand3_1 _22790_ (.B(_09176_),
    .C(_09177_),
    .A(_08937_),
    .Y(_09178_));
 sg13g2_nand3_1 _22791_ (.B(_08773_),
    .C(_09174_),
    .A(net8018),
    .Y(_09179_));
 sg13g2_nand2_1 _22792_ (.Y(_09180_),
    .A(_09178_),
    .B(_09179_));
 sg13g2_mux4_1 _22793_ (.S0(net7905),
    .A0(_01485_),
    .A1(_01520_),
    .A2(_01556_),
    .A3(_01591_),
    .S1(net7817),
    .X(_09181_));
 sg13g2_mux4_1 _22794_ (.S0(net8020),
    .A0(_00554_),
    .A1(_00552_),
    .A2(_00551_),
    .A3(_00553_),
    .S1(net8021),
    .X(_09182_));
 sg13g2_a21oi_1 _22795_ (.A1(_08773_),
    .A2(_09182_),
    .Y(_09183_),
    .B1(net8018));
 sg13g2_nor2_1 _22796_ (.A(_08773_),
    .B(_09182_),
    .Y(_09184_));
 sg13g2_nand2b_1 _22797_ (.Y(_09185_),
    .B(net8022),
    .A_N(_00558_));
 sg13g2_o21ai_1 _22798_ (.B1(_09185_),
    .Y(_09186_),
    .A1(_00557_),
    .A2(net8022));
 sg13g2_a22oi_1 _22799_ (.Y(_09187_),
    .B1(_09186_),
    .B2(net8020),
    .A2(_08758_),
    .A1(_05113_));
 sg13g2_nor2_1 _22800_ (.A(_05201_),
    .B(_09187_),
    .Y(_09188_));
 sg13g2_nor4_1 _22801_ (.A(_00534_),
    .B(_09183_),
    .C(_09184_),
    .D(_09188_),
    .Y(_09189_));
 sg13g2_a221oi_1 _22802_ (.B2(_00534_),
    .C1(_09189_),
    .B1(_09180_),
    .A1(_09173_),
    .Y(_09190_),
    .A2(_09175_));
 sg13g2_or2_1 _22803_ (.X(_09191_),
    .B(_09190_),
    .A(_09171_));
 sg13g2_o21ai_1 _22804_ (.B1(_05186_),
    .Y(_09192_),
    .A1(net7477),
    .A2(net7284));
 sg13g2_a22oi_1 _22805_ (.Y(_09193_),
    .B1(net6743),
    .B2(net7997),
    .A2(_00540_),
    .A1(_00568_));
 sg13g2_nand4_1 _22806_ (.B(_09191_),
    .C(_09192_),
    .A(_09146_),
    .Y(_09194_),
    .D(_09193_));
 sg13g2_a22oi_1 _22807_ (.Y(_09195_),
    .B1(_09194_),
    .B2(net7286),
    .A2(net7085),
    .A1(_00078_));
 sg13g2_o21ai_1 _22808_ (.B1(_09142_),
    .Y(_09196_),
    .A1(net6810),
    .A2(_09195_));
 sg13g2_or3_1 _22809_ (.A(_08242_),
    .B(_03608_),
    .C(net6823),
    .X(_09197_));
 sg13g2_a21oi_1 _22810_ (.A1(_08032_),
    .A2(_07152_),
    .Y(_09198_),
    .B1(_09197_));
 sg13g2_a21o_1 _22811_ (.A2(net6822),
    .A1(_01631_),
    .B1(_09198_),
    .X(_09199_));
 sg13g2_nand2_1 _22812_ (.Y(_09200_),
    .A(_01630_),
    .B(net6821));
 sg13g2_nor2_1 _22813_ (.A(net7259),
    .B(net7126),
    .Y(_09201_));
 sg13g2_a21oi_1 _22814_ (.A1(net6569),
    .A2(net7121),
    .Y(_09202_),
    .B1(_09201_));
 sg13g2_o21ai_1 _22815_ (.B1(_09200_),
    .Y(_09203_),
    .A1(net6821),
    .A2(_09202_));
 sg13g2_nand2_1 _22816_ (.Y(_09204_),
    .A(_01629_),
    .B(net6818));
 sg13g2_nor2b_1 _22817_ (.A(net7127),
    .B_N(_10750_),
    .Y(_09205_));
 sg13g2_a21oi_1 _22818_ (.A1(net6640),
    .A2(net7123),
    .Y(_09206_),
    .B1(_09205_));
 sg13g2_o21ai_1 _22819_ (.B1(_09204_),
    .Y(_09207_),
    .A1(net6818),
    .A2(_09206_));
 sg13g2_nand2_1 _22820_ (.Y(_09208_),
    .A(_01628_),
    .B(net6822));
 sg13g2_nor2_1 _22821_ (.A(_03473_),
    .B(net7126),
    .Y(_09209_));
 sg13g2_a21oi_1 _22822_ (.A1(net459),
    .A2(_04742_),
    .Y(_09210_),
    .B1(_09209_));
 sg13g2_o21ai_1 _22823_ (.B1(_09208_),
    .Y(_09211_),
    .A1(net6822),
    .A2(_09210_));
 sg13g2_nand2_1 _22824_ (.Y(_09212_),
    .A(_01627_),
    .B(net6813));
 sg13g2_nor2_1 _22825_ (.A(net7260),
    .B(net7126),
    .Y(_09213_));
 sg13g2_a21oi_1 _22826_ (.A1(net6572),
    .A2(net7121),
    .Y(_09214_),
    .B1(_09213_));
 sg13g2_o21ai_1 _22827_ (.B1(_09212_),
    .Y(_09215_),
    .A1(net6813),
    .A2(_09214_));
 sg13g2_nand2_1 _22828_ (.Y(_09216_),
    .A(_01626_),
    .B(net6816));
 sg13g2_nor2b_1 _22829_ (.A(net7125),
    .B_N(_03327_),
    .Y(_09217_));
 sg13g2_a21oi_1 _22830_ (.A1(net6574),
    .A2(net7122),
    .Y(_09218_),
    .B1(_09217_));
 sg13g2_o21ai_1 _22831_ (.B1(_09216_),
    .Y(_09219_),
    .A1(net6816),
    .A2(_09218_));
 sg13g2_nand2_1 _22832_ (.Y(_09220_),
    .A(_01625_),
    .B(net6814));
 sg13g2_nor2b_1 _22833_ (.A(net7125),
    .B_N(_03256_),
    .Y(_09221_));
 sg13g2_mux4_1 _22834_ (.S0(net7905),
    .A0(_01344_),
    .A1(_01380_),
    .A2(_01415_),
    .A3(_01450_),
    .S1(net7817),
    .X(_09222_));
 sg13g2_a21oi_1 _22835_ (.A1(net456),
    .A2(net7122),
    .Y(_09223_),
    .B1(_09221_));
 sg13g2_o21ai_1 _22836_ (.B1(_09220_),
    .Y(_09224_),
    .A1(net6814),
    .A2(_09223_));
 sg13g2_nand2_1 _22837_ (.Y(_09225_),
    .A(_01624_),
    .B(net6820));
 sg13g2_nor2_1 _22838_ (.A(_03192_),
    .B(net7126),
    .Y(_09226_));
 sg13g2_a21oi_1 _22839_ (.A1(net6578),
    .A2(net7121),
    .Y(_09227_),
    .B1(_09226_));
 sg13g2_o21ai_1 _22840_ (.B1(_09225_),
    .Y(_09228_),
    .A1(net6820),
    .A2(_09227_));
 sg13g2_nand2_1 _22841_ (.Y(_09229_),
    .A(_01623_),
    .B(net6823));
 sg13g2_nor2_1 _22842_ (.A(_03122_),
    .B(net7125),
    .Y(_09230_));
 sg13g2_mux2_1 _22843_ (.A0(_09181_),
    .A1(_09222_),
    .S(net7486),
    .X(_09231_));
 sg13g2_a21oi_1 _22844_ (.A1(net6581),
    .A2(net7122),
    .Y(_09232_),
    .B1(_09230_));
 sg13g2_o21ai_1 _22845_ (.B1(_09229_),
    .Y(_09233_),
    .A1(net6823),
    .A2(_09232_));
 sg13g2_nand2_1 _22846_ (.Y(_09234_),
    .A(_01622_),
    .B(net6821));
 sg13g2_nand2_1 _22847_ (.Y(_09235_),
    .A(net7498),
    .B(_09231_));
 sg13g2_nor2_1 _22848_ (.A(_03053_),
    .B(net7129),
    .Y(_09236_));
 sg13g2_a21oi_1 _22849_ (.A1(net453),
    .A2(net7121),
    .Y(_09237_),
    .B1(_09236_));
 sg13g2_o21ai_1 _22850_ (.B1(_09234_),
    .Y(_09238_),
    .A1(net6821),
    .A2(_09237_));
 sg13g2_nand2_1 _22851_ (.Y(_09239_),
    .A(_01621_),
    .B(net6813));
 sg13g2_nor2_1 _22852_ (.A(_02986_),
    .B(net7125),
    .Y(_09240_));
 sg13g2_a21oi_1 _22853_ (.A1(net452),
    .A2(net7122),
    .Y(_09241_),
    .B1(_09240_));
 sg13g2_o21ai_1 _22854_ (.B1(_09239_),
    .Y(_09242_),
    .A1(net6813),
    .A2(_09241_));
 sg13g2_nand2_1 _22855_ (.Y(_09243_),
    .A(_01620_),
    .B(net6822));
 sg13g2_inv_1 _22856_ (.Y(_09244_),
    .A(net7925));
 sg13g2_a22oi_1 _22857_ (.Y(_09245_),
    .B1(net7503),
    .B2(_09147_),
    .A2(_08967_),
    .A1(net7541));
 sg13g2_nor2_1 _22858_ (.A(_02919_),
    .B(net7126),
    .Y(_09246_));
 sg13g2_a21oi_1 _22859_ (.A1(net451),
    .A2(net7121),
    .Y(_09247_),
    .B1(_09246_));
 sg13g2_o21ai_1 _22860_ (.B1(_09243_),
    .Y(_09248_),
    .A1(net6820),
    .A2(_09247_));
 sg13g2_nand2_1 _22861_ (.Y(_09249_),
    .A(_01619_),
    .B(net6822));
 sg13g2_nor2_1 _22862_ (.A(net7261),
    .B(net7126),
    .Y(_09250_));
 sg13g2_a21oi_1 _22863_ (.A1(net6585),
    .A2(net7121),
    .Y(_09251_),
    .B1(_09250_));
 sg13g2_and3_1 _22864_ (.X(_09252_),
    .A(_09065_),
    .B(_09235_),
    .C(_09245_));
 sg13g2_o21ai_1 _22865_ (.B1(_09249_),
    .Y(_09253_),
    .A1(net6822),
    .A2(_09251_));
 sg13g2_nand3_1 _22866_ (.B(_09235_),
    .C(_09245_),
    .A(_09065_),
    .Y(_09254_));
 sg13g2_nand2_1 _22867_ (.Y(_09255_),
    .A(_01618_),
    .B(net6815));
 sg13g2_nor2_1 _22868_ (.A(net7077),
    .B(net7128),
    .Y(_09256_));
 sg13g2_a21oi_1 _22869_ (.A1(net6725),
    .A2(net7124),
    .Y(_09257_),
    .B1(_09256_));
 sg13g2_o21ai_1 _22870_ (.B1(_09255_),
    .Y(_09258_),
    .A1(net6815),
    .A2(_09257_));
 sg13g2_nand2_1 _22871_ (.Y(_09259_),
    .A(_01617_),
    .B(net6814));
 sg13g2_nor2_1 _22872_ (.A(_00543_),
    .B(_00539_),
    .Y(_09260_));
 sg13g2_nor2_1 _22873_ (.A(net7262),
    .B(net7125),
    .Y(_09261_));
 sg13g2_a21oi_1 _22874_ (.A1(net449),
    .A2(net7122),
    .Y(_09262_),
    .B1(_09261_));
 sg13g2_nand2_1 _22875_ (.Y(_09263_),
    .A(_05162_),
    .B(_05180_));
 sg13g2_o21ai_1 _22876_ (.B1(_09259_),
    .Y(_09264_),
    .A1(net6814),
    .A2(_09262_));
 sg13g2_nand2_1 _22877_ (.Y(_09265_),
    .A(_01616_),
    .B(net6817));
 sg13g2_nor2_1 _22878_ (.A(net7263),
    .B(net7127),
    .Y(_09266_));
 sg13g2_a21oi_1 _22879_ (.A1(net448),
    .A2(net7123),
    .Y(_09267_),
    .B1(_09266_));
 sg13g2_o21ai_1 _22880_ (.B1(_09265_),
    .Y(_09268_),
    .A1(net6817),
    .A2(_09267_));
 sg13g2_nand2_1 _22881_ (.Y(_09269_),
    .A(_01615_),
    .B(net6815));
 sg13g2_nor2_1 _22882_ (.A(_02652_),
    .B(net7128),
    .Y(_09270_));
 sg13g2_a21oi_1 _22883_ (.A1(net447),
    .A2(net7124),
    .Y(_09271_),
    .B1(_09270_));
 sg13g2_o21ai_1 _22884_ (.B1(_09269_),
    .Y(_09272_),
    .A1(net6815),
    .A2(_09271_));
 sg13g2_nand2_1 _22885_ (.Y(_09273_),
    .A(_01614_),
    .B(net6815));
 sg13g2_nor2_1 _22886_ (.A(_02585_),
    .B(net7128),
    .Y(_09274_));
 sg13g2_nor3_1 _22887_ (.A(_00542_),
    .B(_00541_),
    .C(_09263_),
    .Y(_09275_));
 sg13g2_a21oi_1 _22888_ (.A1(net6611),
    .A2(net7124),
    .Y(_09276_),
    .B1(_09274_));
 sg13g2_or3_1 _22889_ (.A(net8001),
    .B(_00541_),
    .C(_09263_),
    .X(_09277_));
 sg13g2_o21ai_1 _22890_ (.B1(_09273_),
    .Y(_09278_),
    .A1(net6815),
    .A2(_09276_));
 sg13g2_nand2_1 _22891_ (.Y(_09279_),
    .A(_01613_),
    .B(net6813));
 sg13g2_nor2_1 _22892_ (.A(_02534_),
    .B(net7126),
    .Y(_09280_));
 sg13g2_a21oi_1 _22893_ (.A1(net6612),
    .A2(net7121),
    .Y(_09281_),
    .B1(_09280_));
 sg13g2_inv_1 _22894_ (.Y(_09282_),
    .A(net7927));
 sg13g2_o21ai_1 _22895_ (.B1(_09279_),
    .Y(_09283_),
    .A1(net6813),
    .A2(_09281_));
 sg13g2_nand2_1 _22896_ (.Y(_09284_),
    .A(_01612_),
    .B(net6816));
 sg13g2_nor2_1 _22897_ (.A(_02476_),
    .B(net7128),
    .Y(_09285_));
 sg13g2_a21oi_1 _22898_ (.A1(net6614),
    .A2(net7124),
    .Y(_09286_),
    .B1(_09285_));
 sg13g2_o21ai_1 _22899_ (.B1(_09284_),
    .Y(_09287_),
    .A1(net6816),
    .A2(_09286_));
 sg13g2_nand2b_1 _22900_ (.Y(_09288_),
    .B(net8000),
    .A_N(_01632_));
 sg13g2_nand2_1 _22901_ (.Y(_09289_),
    .A(_01611_),
    .B(net6816));
 sg13g2_nor2_1 _22902_ (.A(net7265),
    .B(net7128),
    .Y(_09290_));
 sg13g2_a21oi_1 _22903_ (.A1(net6599),
    .A2(net7124),
    .Y(_09291_),
    .B1(_09290_));
 sg13g2_o21ai_1 _22904_ (.B1(_09288_),
    .Y(_09292_),
    .A1(_01607_),
    .A2(net7479));
 sg13g2_o21ai_1 _22905_ (.B1(_09289_),
    .Y(_09293_),
    .A1(net6816),
    .A2(_09291_));
 sg13g2_nand2_1 _22906_ (.Y(_09294_),
    .A(_01610_),
    .B(net6815));
 sg13g2_nor2_1 _22907_ (.A(net7266),
    .B(net7128),
    .Y(_09295_));
 sg13g2_a21oi_1 _22908_ (.A1(net6602),
    .A2(net7124),
    .Y(_09296_),
    .B1(_09295_));
 sg13g2_o21ai_1 _22909_ (.B1(_09294_),
    .Y(_09297_),
    .A1(net6817),
    .A2(_09296_));
 sg13g2_nand2_1 _22910_ (.Y(_09298_),
    .A(_01609_),
    .B(net6817));
 sg13g2_nor2_1 _22911_ (.A(net7269),
    .B(net7127),
    .Y(_09299_));
 sg13g2_a21oi_1 _22912_ (.A1(net441),
    .A2(net7123),
    .Y(_09300_),
    .B1(_09299_));
 sg13g2_o21ai_1 _22913_ (.B1(_09298_),
    .Y(_09301_),
    .A1(net6817),
    .A2(_09300_));
 sg13g2_nand2_1 _22914_ (.Y(_09302_),
    .A(_01608_),
    .B(net6817));
 sg13g2_nor2b_1 _22915_ (.A(net7127),
    .B_N(_02171_),
    .Y(_09303_));
 sg13g2_a221oi_1 _22916_ (.B2(net7103),
    .C1(_09292_),
    .B1(net7354),
    .A1(net8006),
    .Y(_09304_),
    .A2(_09252_));
 sg13g2_a21oi_1 _22917_ (.A1(net6623),
    .A2(net7123),
    .Y(_09305_),
    .B1(_09303_));
 sg13g2_o21ai_1 _22918_ (.B1(_09302_),
    .Y(_09306_),
    .A1(net6819),
    .A2(_09305_));
 sg13g2_nand2_1 _22919_ (.Y(_09307_),
    .A(_01607_),
    .B(net6818));
 sg13g2_nor2_1 _22920_ (.A(net7103),
    .B(net7127),
    .Y(_09308_));
 sg13g2_a21oi_1 _22921_ (.A1(net6747),
    .A2(net7123),
    .Y(_09309_),
    .B1(_09308_));
 sg13g2_nand2b_1 _22922_ (.Y(_09310_),
    .B(net7385),
    .A_N(_09304_));
 sg13g2_o21ai_1 _22923_ (.B1(_09307_),
    .Y(_09311_),
    .A1(net6818),
    .A2(_09309_));
 sg13g2_nand2_1 _22924_ (.Y(_09312_),
    .A(_02201_),
    .B(_07024_));
 sg13g2_nor3_1 _22925_ (.A(_07035_),
    .B(_07039_),
    .C(_09312_),
    .Y(_09313_));
 sg13g2_o21ai_1 _22926_ (.B1(_09310_),
    .Y(_09314_),
    .A1(net6981),
    .A2(_08873_));
 sg13g2_nor3_1 _22927_ (.A(_02201_),
    .B(_08696_),
    .C(_06960_),
    .Y(_09315_));
 sg13g2_o21ai_1 _22928_ (.B1(_06641_),
    .Y(_09316_),
    .A1(_06600_),
    .A2(_09315_));
 sg13g2_o21ai_1 _22929_ (.B1(net7981),
    .Y(_09317_),
    .A1(_06599_),
    .A2(_07030_));
 sg13g2_a21oi_1 _22930_ (.A1(_09316_),
    .A2(_09317_),
    .Y(_09318_),
    .B1(_09313_));
 sg13g2_and2_1 _22931_ (.A(\load_store_unit_i.data_we_q ),
    .B(_06963_),
    .X(_09319_));
 sg13g2_and2_1 _22932_ (.A(net7313),
    .B(_07691_),
    .X(_09320_));
 sg13g2_nand2_1 _22933_ (.Y(_09321_),
    .A(net7313),
    .B(_07691_));
 sg13g2_nand2_1 _22934_ (.Y(_09322_),
    .A(net7985),
    .B(net7078));
 sg13g2_nand3_1 _22935_ (.B(_02226_),
    .C(_09322_),
    .A(net434),
    .Y(_09323_));
 sg13g2_inv_1 _22936_ (.Y(_09324_),
    .A(net7929));
 sg13g2_a21oi_1 _22937_ (.A1(net7983),
    .A2(net7078),
    .Y(_09325_),
    .B1(\id_stage_i.controller_i.nmi_mode_d ));
 sg13g2_a21oi_1 _22938_ (.A1(_02211_),
    .A2(_09323_),
    .Y(_09326_),
    .B1(_09325_));
 sg13g2_nor2_1 _22939_ (.A(\load_store_unit_i.data_we_q ),
    .B(_06964_),
    .Y(_09327_));
 sg13g2_nor4_1 _22940_ (.A(_01601_),
    .B(_06910_),
    .C(_07091_),
    .D(_07661_),
    .Y(_09328_));
 sg13g2_nor2_1 _22941_ (.A(_06770_),
    .B(_06957_),
    .Y(_09329_));
 sg13g2_nor2_1 _22942_ (.A(_06916_),
    .B(_09329_),
    .Y(_09330_));
 sg13g2_a21oi_1 _22943_ (.A1(_06641_),
    .A2(_09330_),
    .Y(_09331_),
    .B1(_08444_));
 sg13g2_nor2_1 _22944_ (.A(_06781_),
    .B(_09331_),
    .Y(_09332_));
 sg13g2_nor2_1 _22945_ (.A(_09328_),
    .B(_09332_),
    .Y(_09333_));
 sg13g2_a21oi_1 _22946_ (.A1(_06783_),
    .A2(_06958_),
    .Y(_09334_),
    .B1(_09328_));
 sg13g2_a21oi_1 _22947_ (.A1(net7984),
    .A2(_07693_),
    .Y(_09335_),
    .B1(_07657_));
 sg13g2_a22oi_1 _22948_ (.Y(_09336_),
    .B1(_07693_),
    .B2(net7985),
    .A2(_06908_),
    .A1(_01600_));
 sg13g2_nor2_1 _22949_ (.A(net7984),
    .B(_09336_),
    .Y(_09337_));
 sg13g2_nor2_1 _22950_ (.A(_09335_),
    .B(_09337_),
    .Y(_09338_));
 sg13g2_a21oi_1 _22951_ (.A1(_07017_),
    .A2(_07041_),
    .Y(_09339_),
    .B1(_01601_));
 sg13g2_nand2_1 _22952_ (.Y(_09340_),
    .A(_06977_),
    .B(_07004_));
 sg13g2_nor2_1 _22953_ (.A(_09339_),
    .B(_09340_),
    .Y(_09341_));
 sg13g2_nor4_1 _22954_ (.A(net349),
    .B(net7984),
    .C(\cs_registers_i.debug_single_step_o ),
    .D(_07002_),
    .Y(_09342_));
 sg13g2_a21o_1 _22955_ (.A2(_09342_),
    .A1(_01606_),
    .B1(_01602_),
    .X(_09343_));
 sg13g2_nor2_1 _22956_ (.A(_07005_),
    .B(net5968),
    .Y(_09344_));
 sg13g2_nand2_1 _22957_ (.Y(_09345_),
    .A(_06966_),
    .B(_07691_));
 sg13g2_a21o_1 _22958_ (.A2(_08873_),
    .A1(net6917),
    .B1(_09314_),
    .X(_09346_));
 sg13g2_o21ai_1 _22959_ (.B1(_09345_),
    .Y(_09347_),
    .A1(_06978_),
    .A2(_07086_));
 sg13g2_o21ai_1 _22960_ (.B1(_06978_),
    .Y(_09348_),
    .A1(_06899_),
    .A2(_06906_));
 sg13g2_a21oi_1 _22961_ (.A1(_09347_),
    .A2(_09348_),
    .Y(_09349_),
    .B1(_07659_));
 sg13g2_a21oi_1 _22962_ (.A1(_01601_),
    .A2(_07043_),
    .Y(_09350_),
    .B1(_07017_));
 sg13g2_o21ai_1 _22963_ (.B1(_09349_),
    .Y(_09351_),
    .A1(_09344_),
    .A2(_09350_));
 sg13g2_nor3_1 _22964_ (.A(_06900_),
    .B(_06906_),
    .C(_07673_),
    .Y(_09352_));
 sg13g2_and3_1 _22965_ (.X(_09353_),
    .A(_06779_),
    .B(_07691_),
    .C(_09348_));
 sg13g2_nand2_1 _22966_ (.Y(_09354_),
    .A(_01601_),
    .B(_07005_));
 sg13g2_nand2b_1 _22967_ (.Y(_09355_),
    .B(_01606_),
    .A_N(_09342_));
 sg13g2_nor2b_1 _22968_ (.A(_01604_),
    .B_N(_09355_),
    .Y(_09356_));
 sg13g2_o21ai_1 _22969_ (.B1(_09356_),
    .Y(_09357_),
    .A1(_07043_),
    .A2(_09354_));
 sg13g2_o21ai_1 _22970_ (.B1(net7985),
    .Y(_09358_),
    .A1(_06899_),
    .A2(_06906_));
 sg13g2_a21oi_1 _22971_ (.A1(_09339_),
    .A2(_09358_),
    .Y(_09359_),
    .B1(_06979_));
 sg13g2_a22oi_1 _22972_ (.Y(_09360_),
    .B1(_08673_),
    .B2(net7679),
    .A2(_07608_),
    .A1(_08622_));
 sg13g2_o21ai_1 _22973_ (.B1(_06770_),
    .Y(_09361_),
    .A1(_07562_),
    .A2(_09360_));
 sg13g2_nand2_1 _22974_ (.Y(_09362_),
    .A(_07031_),
    .B(_09361_));
 sg13g2_nand2_1 _22975_ (.Y(_09363_),
    .A(_08819_),
    .B(_08836_));
 sg13g2_nor4_2 _22976_ (.A(_06768_),
    .B(_06916_),
    .C(_09329_),
    .Y(_09364_),
    .D(_09362_));
 sg13g2_or4_1 _22977_ (.A(_06768_),
    .B(_06916_),
    .C(_09329_),
    .D(_09362_),
    .X(_09365_));
 sg13g2_nor2b_1 _22978_ (.A(_01986_),
    .B_N(_01987_),
    .Y(_09366_));
 sg13g2_nor2b_1 _22979_ (.A(net7653),
    .B_N(net341),
    .Y(_09367_));
 sg13g2_a21oi_1 _22980_ (.A1(_01989_),
    .A2(net7652),
    .Y(_09368_),
    .B1(_09367_));
 sg13g2_nor2_1 _22981_ (.A(net7645),
    .B(_09368_),
    .Y(_09369_));
 sg13g2_a21oi_1 _22982_ (.A1(_01997_),
    .A2(net7475),
    .Y(_09370_),
    .B1(_09369_));
 sg13g2_nor2_1 _22983_ (.A(net7664),
    .B(_09370_),
    .Y(_09371_));
 sg13g2_nor2_1 _22984_ (.A(net7661),
    .B(_01981_),
    .Y(_09372_));
 sg13g2_inv_1 _22985_ (.Y(_09373_),
    .A(_01888_));
 sg13g2_a21oi_1 _22986_ (.A1(net318),
    .A2(net7652),
    .Y(_09374_),
    .B1(_09367_));
 sg13g2_nor2_1 _22987_ (.A(net7643),
    .B(_09374_),
    .Y(_09375_));
 sg13g2_a21oi_1 _22988_ (.A1(net326),
    .A2(net7476),
    .Y(_09376_),
    .B1(_09375_));
 sg13g2_and2_1 _22989_ (.A(_01987_),
    .B(net7656),
    .X(_09377_));
 sg13g2_nor2_1 _22990_ (.A(net7661),
    .B(_06077_),
    .Y(_09378_));
 sg13g2_nor2b_1 _22991_ (.A(_09378_),
    .B_N(_09377_),
    .Y(_09379_));
 sg13g2_and3_1 _22992_ (.X(_09380_),
    .A(\id_stage_i.controller_i.instr_is_compressed_i ),
    .B(_08819_),
    .C(_08836_));
 sg13g2_and2_1 _22993_ (.A(_01981_),
    .B(_09377_),
    .X(_09381_));
 sg13g2_a221oi_1 _22994_ (.B2(net335),
    .C1(_09371_),
    .B1(_09381_),
    .A1(_02005_),
    .Y(_09382_),
    .A2(_09379_));
 sg13g2_o21ai_1 _22995_ (.B1(_09382_),
    .Y(_09383_),
    .A1(_09372_),
    .A2(_09376_));
 sg13g2_and2_1 _22996_ (.A(net6984),
    .B(net6639),
    .X(_09384_));
 sg13g2_xor2_1 _22997_ (.B(net7104),
    .A(_08158_),
    .X(_09385_));
 sg13g2_or3_1 _22998_ (.A(_08016_),
    .B(net7046),
    .C(_09385_),
    .X(_09386_));
 sg13g2_and3_1 _22999_ (.X(_09387_),
    .A(net7104),
    .B(_08208_),
    .C(_06749_));
 sg13g2_nand3_1 _23000_ (.B(_08208_),
    .C(_06749_),
    .A(net7104),
    .Y(_09388_));
 sg13g2_nor3_1 _23001_ (.A(net7438),
    .B(_08012_),
    .C(_08153_),
    .Y(_09389_));
 sg13g2_nand2_1 _23002_ (.Y(_09390_),
    .A(_08014_),
    .B(_08158_));
 sg13g2_nand3_1 _23003_ (.B(net7027),
    .C(net6972),
    .A(net6953),
    .Y(_09391_));
 sg13g2_o21ai_1 _23004_ (.B1(_09391_),
    .Y(_09392_),
    .A1(net7027),
    .A2(net6906));
 sg13g2_and2_1 _23005_ (.A(net6912),
    .B(_09388_),
    .X(_09393_));
 sg13g2_nand2_1 _23006_ (.Y(_09394_),
    .A(_09386_),
    .B(_09388_));
 sg13g2_nand2_1 _23007_ (.Y(_09395_),
    .A(net7027),
    .B(net6880));
 sg13g2_a22oi_1 _23008_ (.Y(_09396_),
    .B1(_09395_),
    .B2(_11684_),
    .A2(_09392_),
    .A1(net6908));
 sg13g2_a21oi_1 _23009_ (.A1(_08785_),
    .A2(_08838_),
    .Y(_09397_),
    .B1(_08819_));
 sg13g2_nor2b_1 _23010_ (.A(_08208_),
    .B_N(_08195_),
    .Y(_09398_));
 sg13g2_nor2b_1 _23011_ (.A(_08126_),
    .B_N(_09398_),
    .Y(_09399_));
 sg13g2_nand2b_1 _23012_ (.Y(_09400_),
    .B(_09398_),
    .A_N(net7046));
 sg13g2_and2_1 _23013_ (.A(_07557_),
    .B(_06800_),
    .X(_09401_));
 sg13g2_xnor2_1 _23014_ (.Y(_09402_),
    .A(net6953),
    .B(_09401_));
 sg13g2_xnor2_1 _23015_ (.Y(_09403_),
    .A(_11684_),
    .B(_09401_));
 sg13g2_nor2_1 _23016_ (.A(_07555_),
    .B(_06801_),
    .Y(_09404_));
 sg13g2_xnor2_1 _23017_ (.Y(_09405_),
    .A(net6951),
    .B(_09404_));
 sg13g2_xnor2_1 _23018_ (.Y(_09406_),
    .A(net6949),
    .B(_09404_));
 sg13g2_nand2_1 _23019_ (.Y(_09407_),
    .A(_07557_),
    .B(_06799_));
 sg13g2_xnor2_1 _23020_ (.Y(_09408_),
    .A(_10789_),
    .B(_09407_));
 sg13g2_xnor2_1 _23021_ (.Y(_09409_),
    .A(net6901),
    .B(_09407_));
 sg13g2_nand3_1 _23022_ (.B(_08195_),
    .C(_08202_),
    .A(net7046),
    .Y(_09410_));
 sg13g2_nand2_1 _23023_ (.Y(_09411_),
    .A(_06799_),
    .B(_09410_));
 sg13g2_nand2_1 _23024_ (.Y(_09412_),
    .A(_03811_),
    .B(_09400_));
 sg13g2_o21ai_1 _23025_ (.B1(_09412_),
    .Y(_09413_),
    .A1(net7072),
    .A2(_09400_));
 sg13g2_nor2_1 _23026_ (.A(_09408_),
    .B(_09413_),
    .Y(_09414_));
 sg13g2_nand2_1 _23027_ (.Y(_09415_),
    .A(_07557_),
    .B(net6977));
 sg13g2_inv_1 _23028_ (.Y(_09416_),
    .A(_09417_));
 sg13g2_xor2_1 _23029_ (.B(_09415_),
    .A(_09945_),
    .X(_09417_));
 sg13g2_nand2_1 _23030_ (.Y(_09418_),
    .A(_03795_),
    .B(_09400_));
 sg13g2_o21ai_1 _23031_ (.B1(_09418_),
    .Y(_09419_),
    .A1(net7027),
    .A2(_09400_));
 sg13g2_nand2b_1 _23032_ (.Y(_09420_),
    .B(net6969),
    .A_N(net7026));
 sg13g2_a221oi_1 _23033_ (.B2(_01916_),
    .C1(_09380_),
    .B1(_09397_),
    .A1(net7734),
    .Y(_09421_),
    .A2(_08800_));
 sg13g2_o21ai_1 _23034_ (.B1(_09420_),
    .Y(_09422_),
    .A1(net7008),
    .A2(net6969));
 sg13g2_mux2_1 _23035_ (.A0(_09419_),
    .A1(_09422_),
    .S(net6916),
    .X(_09423_));
 sg13g2_and2_1 _23036_ (.A(net6842),
    .B(_09423_),
    .X(_09424_));
 sg13g2_nand2_1 _23037_ (.Y(_09425_),
    .A(net7029),
    .B(_09399_));
 sg13g2_o21ai_1 _23038_ (.B1(_09425_),
    .Y(_09426_),
    .A1(net7006),
    .A2(net6965));
 sg13g2_nor2_1 _23039_ (.A(net6913),
    .B(_09426_),
    .Y(_09427_));
 sg13g2_nor2b_1 _23040_ (.A(_09421_),
    .B_N(_08851_),
    .Y(_09428_));
 sg13g2_mux2_1 _23041_ (.A0(net7028),
    .A1(net7007),
    .S(net6960),
    .X(_09429_));
 sg13g2_a21oi_1 _23042_ (.A1(net6913),
    .A2(_09429_),
    .Y(_09430_),
    .B1(_09427_));
 sg13g2_a21oi_1 _23043_ (.A1(net6874),
    .A2(_09430_),
    .Y(_09431_),
    .B1(_09424_));
 sg13g2_a22oi_1 _23044_ (.Y(_09432_),
    .B1(_09431_),
    .B2(_09408_),
    .A2(_09414_),
    .A1(_09411_));
 sg13g2_nand2_1 _23045_ (.Y(_09433_),
    .A(net6755),
    .B(_09432_));
 sg13g2_nor2b_1 _23046_ (.A(net7773),
    .B_N(_00725_),
    .Y(_09434_));
 sg13g2_mux2_1 _23047_ (.A0(net7017),
    .A1(net7013),
    .S(net6959),
    .X(_09435_));
 sg13g2_mux2_1 _23048_ (.A0(net7016),
    .A1(net7014),
    .S(net6959),
    .X(_09436_));
 sg13g2_mux2_1 _23049_ (.A0(_09435_),
    .A1(_09436_),
    .S(net6914),
    .X(_09437_));
 sg13g2_xnor2_1 _23050_ (.Y(_09438_),
    .A(net6976),
    .B(net6968));
 sg13g2_nand2_1 _23051_ (.Y(_09439_),
    .A(_03729_),
    .B(_09438_));
 sg13g2_o21ai_1 _23052_ (.B1(_09439_),
    .Y(_09440_),
    .A1(net7015),
    .A2(_09438_));
 sg13g2_nor2_1 _23053_ (.A(net6873),
    .B(_09440_),
    .Y(_09441_));
 sg13g2_a21oi_1 _23054_ (.A1(net6873),
    .A2(_09437_),
    .Y(_09442_),
    .B1(_09441_));
 sg13g2_o21ai_1 _23055_ (.B1(net7705),
    .Y(_09443_),
    .A1(_08285_),
    .A2(_09434_));
 sg13g2_mux2_1 _23056_ (.A0(net7018),
    .A1(net7012),
    .S(net6967),
    .X(_09444_));
 sg13g2_nor2_1 _23057_ (.A(net7019),
    .B(net6967),
    .Y(_09445_));
 sg13g2_a21oi_1 _23058_ (.A1(_03754_),
    .A2(net6967),
    .Y(_09446_),
    .B1(_09445_));
 sg13g2_mux2_1 _23059_ (.A0(_09444_),
    .A1(_09446_),
    .S(net6914),
    .X(_09447_));
 sg13g2_mux2_1 _23060_ (.A0(net7016),
    .A1(net7014),
    .S(net6967),
    .X(_09448_));
 sg13g2_nand2_1 _23061_ (.Y(_09449_),
    .A(net6974),
    .B(_09448_));
 sg13g2_nand2b_1 _23062_ (.Y(_09450_),
    .B(net6967),
    .A_N(net7013));
 sg13g2_o21ai_1 _23063_ (.B1(_09450_),
    .Y(_09451_),
    .A1(net7017),
    .A2(net6967));
 sg13g2_o21ai_1 _23064_ (.B1(_09449_),
    .Y(_09452_),
    .A1(net6974),
    .A2(_09451_));
 sg13g2_mux2_1 _23065_ (.A0(_09447_),
    .A1(_09452_),
    .S(net6872),
    .X(_09453_));
 sg13g2_nor2_1 _23066_ (.A(net6844),
    .B(_09453_),
    .Y(_09454_));
 sg13g2_a21oi_1 _23067_ (.A1(net6844),
    .A2(_09442_),
    .Y(_09455_),
    .B1(_09454_));
 sg13g2_o21ai_1 _23068_ (.B1(_09433_),
    .Y(_09456_),
    .A1(net6755),
    .A2(_09455_));
 sg13g2_nor2_1 _23069_ (.A(net6801),
    .B(_09456_),
    .Y(_09457_));
 sg13g2_nand2_1 _23070_ (.Y(_09458_),
    .A(_03754_),
    .B(net6959));
 sg13g2_o21ai_1 _23071_ (.B1(_09458_),
    .Y(_09459_),
    .A1(net7019),
    .A2(net6959));
 sg13g2_mux2_1 _23072_ (.A0(_00661_),
    .A1(_00693_),
    .S(net7779),
    .X(_09460_));
 sg13g2_nand2b_1 _23073_ (.Y(_09461_),
    .B(net6967),
    .A_N(net7018));
 sg13g2_o21ai_1 _23074_ (.B1(_09461_),
    .Y(_09462_),
    .A1(net7012),
    .A2(net6967));
 sg13g2_mux2_1 _23075_ (.A0(_09459_),
    .A1(_09462_),
    .S(net6914),
    .X(_09463_));
 sg13g2_nand2_1 _23076_ (.Y(_09464_),
    .A(_03764_),
    .B(net6959));
 sg13g2_inv_1 _23077_ (.Y(_09465_),
    .A(_09466_));
 sg13g2_o21ai_1 _23078_ (.B1(_09464_),
    .Y(_09466_),
    .A1(net7021),
    .A2(net6959));
 sg13g2_nor2_1 _23079_ (.A(net7020),
    .B(net6959),
    .Y(_09467_));
 sg13g2_a21oi_1 _23080_ (.A1(_03759_),
    .A2(net6959),
    .Y(_09468_),
    .B1(_09467_));
 sg13g2_nor3_1 _23081_ (.A(net7696),
    .B(net7729),
    .C(_09460_),
    .Y(_09469_));
 sg13g2_mux2_1 _23082_ (.A0(_09465_),
    .A1(_09468_),
    .S(net6915),
    .X(_09470_));
 sg13g2_nor2_1 _23083_ (.A(net6843),
    .B(_09470_),
    .Y(_09471_));
 sg13g2_a21oi_1 _23084_ (.A1(net6843),
    .A2(_09463_),
    .Y(_09472_),
    .B1(_09471_));
 sg13g2_nand2_1 _23085_ (.Y(_09473_),
    .A(_09408_),
    .B(_09472_));
 sg13g2_nand2b_1 _23086_ (.Y(_09474_),
    .B(net6966),
    .A_N(net7023));
 sg13g2_o21ai_1 _23087_ (.B1(_09474_),
    .Y(_09475_),
    .A1(net7010),
    .A2(net6966));
 sg13g2_nor2_1 _23088_ (.A(net6915),
    .B(_09475_),
    .Y(_09476_));
 sg13g2_nor2_1 _23089_ (.A(net7011),
    .B(net6968),
    .Y(_09477_));
 sg13g2_a21oi_1 _23090_ (.A1(net7022),
    .A2(net6966),
    .Y(_09478_),
    .B1(_09477_));
 sg13g2_a21oi_1 _23091_ (.A1(net6915),
    .A2(_09478_),
    .Y(_09479_),
    .B1(_09476_));
 sg13g2_nand2_1 _23092_ (.Y(_09480_),
    .A(net6843),
    .B(_09479_));
 sg13g2_nand2_1 _23093_ (.Y(_09481_),
    .A(_03784_),
    .B(net6960));
 sg13g2_o21ai_1 _23094_ (.B1(_09481_),
    .Y(_09482_),
    .A1(net7025),
    .A2(net6960));
 sg13g2_nor2_1 _23095_ (.A(net7024),
    .B(net6960),
    .Y(_09483_));
 sg13g2_a21oi_1 _23096_ (.A1(net7009),
    .A2(net6960),
    .Y(_09484_),
    .B1(_09483_));
 sg13g2_nand2_1 _23097_ (.Y(_09485_),
    .A(net6915),
    .B(_09484_));
 sg13g2_o21ai_1 _23098_ (.B1(_09485_),
    .Y(_09486_),
    .A1(net6916),
    .A2(_09482_));
 sg13g2_o21ai_1 _23099_ (.B1(_09480_),
    .Y(_09487_),
    .A1(net6842),
    .A2(_09486_));
 sg13g2_inv_1 _23100_ (.Y(_09488_),
    .A(_09489_));
 sg13g2_o21ai_1 _23101_ (.B1(_09473_),
    .Y(_09489_),
    .A1(_09408_),
    .A2(_09487_));
 sg13g2_nor2_1 _23102_ (.A(net7011),
    .B(net6960),
    .Y(_09490_));
 sg13g2_a21oi_1 _23103_ (.A1(net7022),
    .A2(net6960),
    .Y(_09491_),
    .B1(_09490_));
 sg13g2_mux2_1 _23104_ (.A0(net7023),
    .A1(net7010),
    .S(net6968),
    .X(_09492_));
 sg13g2_mux2_1 _23105_ (.A0(_09491_),
    .A1(_09492_),
    .S(net6915),
    .X(_09493_));
 sg13g2_nor2_1 _23106_ (.A(net7020),
    .B(net6965),
    .Y(_09494_));
 sg13g2_a21oi_1 _23107_ (.A1(_03759_),
    .A2(net6969),
    .Y(_09495_),
    .B1(_09494_));
 sg13g2_nand2_1 _23108_ (.Y(_09496_),
    .A(net6973),
    .B(_09495_));
 sg13g2_nand2_1 _23109_ (.Y(_09497_),
    .A(_03764_),
    .B(net6966));
 sg13g2_o21ai_1 _23110_ (.B1(_09497_),
    .Y(_09498_),
    .A1(net7021),
    .A2(net6966));
 sg13g2_o21ai_1 _23111_ (.B1(_09496_),
    .Y(_09499_),
    .A1(net6976),
    .A2(_09498_));
 sg13g2_mux2_1 _23112_ (.A0(_09493_),
    .A1(_09499_),
    .S(net6874),
    .X(_09500_));
 sg13g2_nor2_1 _23113_ (.A(net7024),
    .B(net6969),
    .Y(_09501_));
 sg13g2_a21oi_1 _23114_ (.A1(net7009),
    .A2(net6968),
    .Y(_09502_),
    .B1(_09501_));
 sg13g2_nor2_1 _23115_ (.A(net7025),
    .B(net6969),
    .Y(_09503_));
 sg13g2_a21oi_1 _23116_ (.A1(_03784_),
    .A2(net6969),
    .Y(_09504_),
    .B1(_09503_));
 sg13g2_mux2_1 _23117_ (.A0(_09502_),
    .A1(_09504_),
    .S(net6916),
    .X(_09505_));
 sg13g2_nor2_1 _23118_ (.A(net6842),
    .B(_09505_),
    .Y(_09506_));
 sg13g2_mux2_1 _23119_ (.A0(net7026),
    .A1(net7008),
    .S(net6965),
    .X(_09507_));
 sg13g2_nor2_1 _23120_ (.A(net7027),
    .B(net6965),
    .Y(_09508_));
 sg13g2_a21oi_1 _23121_ (.A1(_03795_),
    .A2(net6965),
    .Y(_09509_),
    .B1(_09508_));
 sg13g2_mux2_1 _23122_ (.A0(_09507_),
    .A1(_09509_),
    .S(net6913),
    .X(_09510_));
 sg13g2_nor2_1 _23123_ (.A(net6874),
    .B(_09510_),
    .Y(_09511_));
 sg13g2_nor3_1 _23124_ (.A(net6847),
    .B(_09506_),
    .C(_09511_),
    .Y(_09512_));
 sg13g2_a21oi_1 _23125_ (.A1(net6847),
    .A2(_09500_),
    .Y(_09513_),
    .B1(_09512_));
 sg13g2_nand2_1 _23126_ (.Y(_09514_),
    .A(net6755),
    .B(_09489_));
 sg13g2_mux2_1 _23127_ (.A0(_00923_),
    .A1(_00958_),
    .S(net7778),
    .X(_09515_));
 sg13g2_o21ai_1 _23128_ (.B1(_09514_),
    .Y(_09516_),
    .A1(net6755),
    .A2(_09513_));
 sg13g2_a21oi_1 _23129_ (.A1(net6801),
    .A2(_09516_),
    .Y(_09517_),
    .B1(_09457_));
 sg13g2_nor2_1 _23130_ (.A(_09410_),
    .B(_09413_),
    .Y(_09518_));
 sg13g2_or2_1 _23131_ (.X(_09519_),
    .B(_09413_),
    .A(_09410_));
 sg13g2_nor2_1 _23132_ (.A(net6798),
    .B(net6755),
    .Y(_09520_));
 sg13g2_nor2_1 _23133_ (.A(_09518_),
    .B(_09520_),
    .Y(_09521_));
 sg13g2_nand2_1 _23134_ (.Y(_09522_),
    .A(net6973),
    .B(_09429_));
 sg13g2_o21ai_1 _23135_ (.B1(_09522_),
    .Y(_09523_),
    .A1(net6973),
    .A2(_09419_));
 sg13g2_nor3_1 _23136_ (.A(net7534),
    .B(net7729),
    .C(_09515_),
    .Y(_09524_));
 sg13g2_mux2_1 _23137_ (.A0(_09413_),
    .A1(_09426_),
    .S(net6913),
    .X(_09525_));
 sg13g2_nand2_1 _23138_ (.Y(_09526_),
    .A(net6876),
    .B(_09525_));
 sg13g2_o21ai_1 _23139_ (.B1(_09526_),
    .Y(_09527_),
    .A1(net6876),
    .A2(_09523_));
 sg13g2_nor2_1 _23140_ (.A(net6847),
    .B(_09527_),
    .Y(_09528_));
 sg13g2_nor2_1 _23141_ (.A(_09408_),
    .B(_09519_),
    .Y(_09529_));
 sg13g2_nor2_1 _23142_ (.A(_09528_),
    .B(_09529_),
    .Y(_09530_));
 sg13g2_a21oi_1 _23143_ (.A1(_09520_),
    .A2(_09530_),
    .Y(_09531_),
    .B1(_09521_));
 sg13g2_o21ai_1 _23144_ (.B1(net7294),
    .Y(_09532_),
    .A1(net6957),
    .A2(_09531_));
 sg13g2_a21oi_1 _23145_ (.A1(net6958),
    .A2(_09517_),
    .Y(_09533_),
    .B1(_09532_));
 sg13g2_nor4_1 _23146_ (.A(net7379),
    .B(_09384_),
    .C(_09396_),
    .D(_09533_),
    .Y(_09534_));
 sg13g2_nand2_1 _23147_ (.Y(_09535_),
    .A(net7482),
    .B(_08722_));
 sg13g2_a221oi_1 _23148_ (.B2(_01635_),
    .C1(net7370),
    .B1(_09535_),
    .A1(_00105_),
    .Y(_09536_),
    .A2(_08739_));
 sg13g2_or2_1 _23149_ (.X(_09537_),
    .B(_09536_),
    .A(_09534_));
 sg13g2_a21oi_1 _23150_ (.A1(net6949),
    .A2(_06784_),
    .Y(_09538_),
    .B1(net6888));
 sg13g2_inv_1 _23151_ (.Y(_09539_),
    .A(_09538_));
 sg13g2_and2_1 _23152_ (.A(net6930),
    .B(_06839_),
    .X(_09540_));
 sg13g2_nand2_1 _23153_ (.Y(_09541_),
    .A(net6931),
    .B(_06799_));
 sg13g2_a22oi_1 _23154_ (.Y(_09542_),
    .B1(net6871),
    .B2(_00147_),
    .A2(net6840),
    .A1(_00211_));
 sg13g2_nand2b_1 _23155_ (.Y(_09543_),
    .B(net6711),
    .A_N(_09542_));
 sg13g2_mux2_1 _23156_ (.A0(_00993_),
    .A1(_01029_),
    .S(net7779),
    .X(_09544_));
 sg13g2_a22oi_1 _23157_ (.Y(_09545_),
    .B1(net6867),
    .B2(_00142_),
    .A2(net6841),
    .A1(_00206_));
 sg13g2_or2_1 _23158_ (.X(_09546_),
    .B(_06836_),
    .A(_06815_));
 sg13g2_nor2_1 _23159_ (.A(net6825),
    .B(_09546_),
    .Y(_09547_));
 sg13g2_nand3_1 _23160_ (.B(_06809_),
    .C(_06813_),
    .A(_08874_),
    .Y(_09548_));
 sg13g2_nor2_1 _23161_ (.A(_06818_),
    .B(_06836_),
    .Y(_09549_));
 sg13g2_nor3_1 _23162_ (.A(net7534),
    .B(net7519),
    .C(_09544_),
    .Y(_09550_));
 sg13g2_nor2_1 _23163_ (.A(net6888),
    .B(_06822_),
    .Y(_09551_));
 sg13g2_nand3_1 _23164_ (.B(net6930),
    .C(_06790_),
    .A(_06784_),
    .Y(_09552_));
 sg13g2_nand4_1 _23165_ (.B(net6900),
    .C(net6931),
    .A(net6975),
    .Y(_09553_),
    .D(_06809_));
 sg13g2_nand2_1 _23166_ (.Y(_09554_),
    .A(_06784_),
    .B(_09540_));
 sg13g2_nor3_1 _23167_ (.A(net6826),
    .B(_06807_),
    .C(_06925_),
    .Y(_09555_));
 sg13g2_inv_1 _23168_ (.Y(_09556_),
    .A(_09557_));
 sg13g2_nand2_1 _23169_ (.Y(_09557_),
    .A(net6930),
    .B(_06881_));
 sg13g2_nor2_1 _23170_ (.A(_09546_),
    .B(_09557_),
    .Y(_09558_));
 sg13g2_or4_1 _23171_ (.A(net6950),
    .B(_06811_),
    .C(_06812_),
    .D(_06836_),
    .X(_09559_));
 sg13g2_nor2_1 _23172_ (.A(_09557_),
    .B(_09559_),
    .Y(_09560_));
 sg13g2_nand3_1 _23173_ (.B(net6931),
    .C(_06809_),
    .A(net6975),
    .Y(_09561_));
 sg13g2_nand2b_1 _23174_ (.Y(_09562_),
    .B(net6900),
    .A_N(_09561_));
 sg13g2_nor2_1 _23175_ (.A(_09559_),
    .B(_09562_),
    .Y(_09563_));
 sg13g2_nor4_1 _23176_ (.A(_09443_),
    .B(_09469_),
    .C(_09524_),
    .D(_09550_),
    .Y(_09564_));
 sg13g2_nor2_1 _23177_ (.A(net6794),
    .B(_09559_),
    .Y(_09565_));
 sg13g2_nor2_1 _23178_ (.A(_06871_),
    .B(_09554_),
    .Y(_09566_));
 sg13g2_nor2_1 _23179_ (.A(_06822_),
    .B(_06871_),
    .Y(_09567_));
 sg13g2_nor2_1 _23180_ (.A(_06871_),
    .B(_09562_),
    .Y(_09568_));
 sg13g2_nor3_1 _23181_ (.A(net6950),
    .B(net6826),
    .C(_06872_),
    .Y(_09569_));
 sg13g2_nor2_1 _23182_ (.A(net6826),
    .B(_09559_),
    .Y(_09570_));
 sg13g2_nand2_1 _23183_ (.Y(_09571_),
    .A(net7704),
    .B(_00757_));
 sg13g2_nor2_1 _23184_ (.A(_09552_),
    .B(_09559_),
    .Y(_09572_));
 sg13g2_nand2b_1 _23185_ (.Y(_09573_),
    .B(_01577_),
    .A_N(net7704));
 sg13g2_nand2_1 _23186_ (.Y(_09574_),
    .A(_06829_),
    .B(_06942_));
 sg13g2_nor2_1 _23187_ (.A(net6825),
    .B(_09574_),
    .Y(_09575_));
 sg13g2_a22oi_1 _23188_ (.Y(_09576_),
    .B1(_09575_),
    .B2(_00425_),
    .A2(net6824),
    .A1(net376));
 sg13g2_nor2_1 _23189_ (.A(_06954_),
    .B(net6794),
    .Y(_09577_));
 sg13g2_nor4_1 _23190_ (.A(_08874_),
    .B(net6901),
    .C(net6888),
    .D(_06810_),
    .Y(_09578_));
 sg13g2_nor2b_1 _23191_ (.A(_06954_),
    .B_N(_09578_),
    .Y(_09579_));
 sg13g2_a21oi_1 _23192_ (.A1(_09571_),
    .A2(_09573_),
    .Y(_09580_),
    .B1(net7601));
 sg13g2_a22oi_1 _23193_ (.Y(_09581_),
    .B1(_09579_),
    .B2(_00273_),
    .A2(_09577_),
    .A1(_00305_));
 sg13g2_nor2b_1 _23194_ (.A(_09574_),
    .B_N(_09578_),
    .Y(_09582_));
 sg13g2_nor2_1 _23195_ (.A(_06822_),
    .B(_06954_),
    .Y(_09583_));
 sg13g2_a22oi_1 _23196_ (.Y(_09584_),
    .B1(_09583_),
    .B2(_00337_),
    .A2(_09582_),
    .A1(_00375_));
 sg13g2_nor3_1 _23197_ (.A(net6826),
    .B(_06807_),
    .C(_06946_),
    .Y(_09585_));
 sg13g2_nor2_1 _23198_ (.A(net6794),
    .B(_09574_),
    .Y(_09586_));
 sg13g2_a21oi_1 _23199_ (.A1(_00347_),
    .A2(_09586_),
    .Y(_09587_),
    .B1(_09585_));
 sg13g2_nand4_1 _23200_ (.B(_09581_),
    .C(_09584_),
    .A(_09576_),
    .Y(_09588_),
    .D(_09587_));
 sg13g2_nor2_1 _23201_ (.A(_09552_),
    .B(_09574_),
    .Y(_09589_));
 sg13g2_nand2b_1 _23202_ (.Y(_09590_),
    .B(_06942_),
    .A_N(_06815_));
 sg13g2_nor2_1 _23203_ (.A(_09548_),
    .B(_09590_),
    .Y(_09591_));
 sg13g2_a22oi_1 _23204_ (.Y(_09592_),
    .B1(_09591_),
    .B2(_00390_),
    .A2(_09589_),
    .A1(_00500_));
 sg13g2_nor2_1 _23205_ (.A(_09548_),
    .B(_09574_),
    .Y(_09593_));
 sg13g2_nor2_1 _23206_ (.A(net6825),
    .B(_09590_),
    .Y(_09594_));
 sg13g2_a22oi_1 _23207_ (.Y(_09595_),
    .B1(_09594_),
    .B2(\cs_registers_i.csr_mstatus_mie_o ),
    .A2(_09593_),
    .A1(net435));
 sg13g2_nand2_1 _23208_ (.Y(_09596_),
    .A(_09592_),
    .B(_09595_));
 sg13g2_nand2b_1 _23209_ (.Y(_09597_),
    .B(_06940_),
    .A_N(_09545_));
 sg13g2_a21oi_1 _23210_ (.A1(_09543_),
    .A2(_09597_),
    .Y(_09598_),
    .B1(_09538_));
 sg13g2_nor3_1 _23211_ (.A(_09588_),
    .B(_09596_),
    .C(_09598_),
    .Y(_09599_));
 sg13g2_nand3_1 _23212_ (.B(_09537_),
    .C(_09599_),
    .A(net6549),
    .Y(_09600_));
 sg13g2_o21ai_1 _23213_ (.B1(net6121),
    .Y(_09601_),
    .A1(net6552),
    .A2(_09383_));
 sg13g2_nor4_1 _23214_ (.A(net314),
    .B(\load_store_unit_i.lsu_err_q ),
    .C(\load_store_unit_i.data_we_q ),
    .D(_06961_),
    .Y(_09602_));
 sg13g2_nor2_1 _23215_ (.A(_09364_),
    .B(_09602_),
    .Y(_09603_));
 sg13g2_or2_1 _23216_ (.X(_09604_),
    .B(_09602_),
    .A(_09364_));
 sg13g2_nor2_1 _23217_ (.A(_08510_),
    .B(_01888_),
    .Y(_09605_));
 sg13g2_nand2_1 _23218_ (.Y(_09606_),
    .A(_01915_),
    .B(_09373_));
 sg13g2_nand2_1 _23219_ (.Y(_09607_),
    .A(_01916_),
    .B(_09604_));
 sg13g2_nor2_1 _23220_ (.A(_09606_),
    .B(_09607_),
    .Y(_09608_));
 sg13g2_nand3_1 _23221_ (.B(_09604_),
    .C(_09605_),
    .A(net7668),
    .Y(_09609_));
 sg13g2_nor2_1 _23222_ (.A(_06620_),
    .B(_09609_),
    .Y(_09610_));
 sg13g2_nand2_1 _23223_ (.Y(_09611_),
    .A(_06619_),
    .B(_09608_));
 sg13g2_nand2_1 _23224_ (.Y(_09612_),
    .A(_01599_),
    .B(net6048));
 sg13g2_o21ai_1 _23225_ (.B1(_09612_),
    .Y(_09613_),
    .A1(net6055),
    .A2(net6048));
 sg13g2_nor2b_1 _23226_ (.A(net7648),
    .B_N(net7654),
    .Y(_09614_));
 sg13g2_a22oi_1 _23227_ (.Y(_09615_),
    .B1(_09614_),
    .B2(net322),
    .A2(_09366_),
    .A1(net331));
 sg13g2_nor2_1 _23228_ (.A(net7647),
    .B(net7655),
    .Y(_09616_));
 sg13g2_a22oi_1 _23229_ (.Y(_09617_),
    .B1(_09616_),
    .B2(net345),
    .A2(_09377_),
    .A1(net340));
 sg13g2_nand2b_1 _23230_ (.Y(_09618_),
    .B(_01981_),
    .A_N(_09617_));
 sg13g2_a21oi_1 _23231_ (.A1(_09615_),
    .A2(_09618_),
    .Y(_09619_),
    .B1(_09372_));
 sg13g2_a22oi_1 _23232_ (.Y(_09620_),
    .B1(_09614_),
    .B2(_01993_),
    .A2(_09366_),
    .A1(_02001_));
 sg13g2_nor2_1 _23233_ (.A(_00007_),
    .B(_09620_),
    .Y(_09621_));
 sg13g2_a22oi_1 _23234_ (.Y(_09622_),
    .B1(_09616_),
    .B2(net345),
    .A2(_09377_),
    .A1(_02009_));
 sg13g2_nor2_1 _23235_ (.A(_09378_),
    .B(_09622_),
    .Y(_09623_));
 sg13g2_nor4_1 _23236_ (.A(net6552),
    .B(_09619_),
    .C(_09621_),
    .D(_09623_),
    .Y(_09624_));
 sg13g2_nand3_1 _23237_ (.B(net7023),
    .C(_09390_),
    .A(_15514_),
    .Y(_09625_));
 sg13g2_o21ai_1 _23238_ (.B1(_09625_),
    .Y(_09626_),
    .A1(net7023),
    .A2(_09387_));
 sg13g2_nand2_1 _23239_ (.Y(_09627_),
    .A(net7023),
    .B(net6879));
 sg13g2_a22oi_1 _23240_ (.Y(_09628_),
    .B1(_09627_),
    .B2(_15516_),
    .A2(_09626_),
    .A1(net6909));
 sg13g2_nand2_1 _23241_ (.Y(_09629_),
    .A(net6847),
    .B(_09472_));
 sg13g2_o21ai_1 _23242_ (.B1(_09629_),
    .Y(_09630_),
    .A1(net6847),
    .A2(_09442_));
 sg13g2_a21o_1 _23243_ (.A2(_09410_),
    .A1(_06800_),
    .B1(_09413_),
    .X(_09631_));
 sg13g2_nor2_1 _23244_ (.A(_09405_),
    .B(_09631_),
    .Y(_09632_));
 sg13g2_a21oi_1 _23245_ (.A1(net6756),
    .A2(_09630_),
    .Y(_09633_),
    .B1(_09632_));
 sg13g2_nand2_1 _23246_ (.Y(_09634_),
    .A(_09409_),
    .B(_09431_));
 sg13g2_o21ai_1 _23247_ (.B1(_09634_),
    .Y(_09635_),
    .A1(_09409_),
    .A2(_09487_));
 sg13g2_nand2b_1 _23248_ (.Y(_09636_),
    .B(net6755),
    .A_N(_09635_));
 sg13g2_nand2_1 _23249_ (.Y(_09637_),
    .A(net6846),
    .B(_09453_));
 sg13g2_nand2_1 _23250_ (.Y(_09638_),
    .A(net6851),
    .B(_09500_));
 sg13g2_nand3_1 _23251_ (.B(_09637_),
    .C(_09638_),
    .A(net6758),
    .Y(_09639_));
 sg13g2_nand3_1 _23252_ (.B(_09636_),
    .C(_09639_),
    .A(net6802),
    .Y(_09640_));
 sg13g2_o21ai_1 _23253_ (.B1(_09640_),
    .Y(_09641_),
    .A1(net6801),
    .A2(_09633_));
 sg13g2_a21oi_1 _23254_ (.A1(net6798),
    .A2(_09519_),
    .Y(_09642_),
    .B1(net6754));
 sg13g2_nand2_1 _23255_ (.Y(_09643_),
    .A(net6973),
    .B(_09484_));
 sg13g2_o21ai_1 _23256_ (.B1(_09643_),
    .Y(_09644_),
    .A1(net6973),
    .A2(_09475_));
 sg13g2_nor2_1 _23257_ (.A(net6873),
    .B(_09644_),
    .Y(_09645_));
 sg13g2_mux2_1 _23258_ (.A0(_09422_),
    .A1(_09482_),
    .S(net6916),
    .X(_09646_));
 sg13g2_a21oi_1 _23259_ (.A1(net6873),
    .A2(_09646_),
    .Y(_09647_),
    .B1(_09645_));
 sg13g2_nand2_1 _23260_ (.Y(_09648_),
    .A(net6851),
    .B(_09647_));
 sg13g2_o21ai_1 _23261_ (.B1(_09648_),
    .Y(_09649_),
    .A1(net6851),
    .A2(_09527_));
 sg13g2_o21ai_1 _23262_ (.B1(_09642_),
    .Y(_09650_),
    .A1(net6798),
    .A2(_09649_));
 sg13g2_nor2_1 _23263_ (.A(net6961),
    .B(_09641_),
    .Y(_09651_));
 sg13g2_a21oi_1 _23264_ (.A1(net6961),
    .A2(_09650_),
    .Y(_09652_),
    .B1(_09651_));
 sg13g2_a221oi_1 _23265_ (.B2(net7296),
    .C1(_09628_),
    .B1(_09652_),
    .A1(net6982),
    .Y(_09653_),
    .A2(net6627));
 sg13g2_or2_1 _23266_ (.X(_09654_),
    .B(_09653_),
    .A(net7378));
 sg13g2_mux4_1 _23267_ (.S0(net7778),
    .A0(_00789_),
    .A1(_00821_),
    .A2(_00853_),
    .A3(_00888_),
    .S1(net7729),
    .X(_09655_));
 sg13g2_a22oi_1 _23268_ (.Y(_09656_),
    .B1(net6870),
    .B2(_00175_),
    .A2(net6839),
    .A1(_00239_));
 sg13g2_a22oi_1 _23269_ (.Y(_09657_),
    .B1(net6871),
    .B2(_00146_),
    .A2(net6840),
    .A1(_00210_));
 sg13g2_nor2_1 _23270_ (.A(net7534),
    .B(_09655_),
    .Y(_09658_));
 sg13g2_and2_1 _23271_ (.A(net436),
    .B(_09560_),
    .X(_09659_));
 sg13g2_a221oi_1 _23272_ (.B2(_00277_),
    .C1(_09659_),
    .B1(net6687),
    .A1(_00389_),
    .Y(_09660_),
    .A2(net6706));
 sg13g2_nor2_1 _23273_ (.A(net6825),
    .B(_06871_),
    .Y(_09661_));
 sg13g2_a22oi_1 _23274_ (.Y(_09662_),
    .B1(_09661_),
    .B2(_00247_),
    .A2(net6691),
    .A1(_00341_));
 sg13g2_inv_1 _23275_ (.Y(_09663_),
    .A(_09662_));
 sg13g2_a221oi_1 _23276_ (.B2(_00429_),
    .C1(_09663_),
    .B1(net6679),
    .A1(_00379_),
    .Y(_09664_),
    .A2(net6700));
 sg13g2_a221oi_1 _23277_ (.B2(_00309_),
    .C1(net6682),
    .B1(net6697),
    .A1(net380),
    .Y(_09665_),
    .A2(net6779));
 sg13g2_a22oi_1 _23278_ (.Y(_09666_),
    .B1(net6675),
    .B2(_00504_),
    .A2(_09547_),
    .A1(_05419_));
 sg13g2_nand4_1 _23279_ (.B(_09664_),
    .C(_09665_),
    .A(_09660_),
    .Y(_09667_),
    .D(_09666_));
 sg13g2_nand2b_1 _23280_ (.Y(_09668_),
    .B(net6712),
    .A_N(_09656_));
 sg13g2_o21ai_1 _23281_ (.B1(_09668_),
    .Y(_09669_),
    .A1(net6652),
    .A2(_09657_));
 sg13g2_a21oi_1 _23282_ (.A1(net6796),
    .A2(_09669_),
    .Y(_09670_),
    .B1(_09667_));
 sg13g2_a21oi_1 _23283_ (.A1(net7482),
    .A2(_08722_),
    .Y(_09671_),
    .B1(_08242_));
 sg13g2_nand2_1 _23284_ (.Y(_09672_),
    .A(_01640_),
    .B(_09671_));
 sg13g2_nand3_1 _23285_ (.B(_09670_),
    .C(_09672_),
    .A(net6549),
    .Y(_09673_));
 sg13g2_a221oi_1 _23286_ (.B2(_01225_),
    .C1(net7696),
    .B1(net7594),
    .A1(_00873_),
    .Y(_09674_),
    .A2(net7597));
 sg13g2_nor2_1 _23287_ (.A(net6825),
    .B(_06954_),
    .Y(_09675_));
 sg13g2_nor3_1 _23288_ (.A(net7703),
    .B(_09658_),
    .C(_09674_),
    .Y(_09676_));
 sg13g2_a21oi_1 _23289_ (.A1(_00109_),
    .A2(net7088),
    .Y(_09677_),
    .B1(_09673_));
 sg13g2_a21o_1 _23290_ (.A2(_09677_),
    .A1(_09654_),
    .B1(_09624_),
    .X(_09678_));
 sg13g2_and2_1 _23291_ (.A(_01917_),
    .B(_01887_),
    .X(_09679_));
 sg13g2_nand2_1 _23292_ (.Y(_09680_),
    .A(_01917_),
    .B(_01887_));
 sg13g2_nor2_1 _23293_ (.A(_08510_),
    .B(_09373_),
    .Y(_09681_));
 sg13g2_nand2_1 _23294_ (.Y(_09682_),
    .A(_01915_),
    .B(_01888_));
 sg13g2_nor2_1 _23295_ (.A(_09607_),
    .B(_09682_),
    .Y(_09683_));
 sg13g2_or4_1 _23296_ (.A(net7686),
    .B(_09564_),
    .C(_09580_),
    .D(_09676_),
    .X(_09684_));
 sg13g2_nor3_1 _23297_ (.A(_09607_),
    .B(_09680_),
    .C(_09682_),
    .Y(_09685_));
 sg13g2_nand2_1 _23298_ (.Y(_09686_),
    .A(net7474),
    .B(_09683_));
 sg13g2_nand2_1 _23299_ (.Y(_09687_),
    .A(_01598_),
    .B(net6034));
 sg13g2_o21ai_1 _23300_ (.B1(_09687_),
    .Y(_09688_),
    .A1(net6119),
    .A2(net6034));
 sg13g2_nor2b_1 _23301_ (.A(net7654),
    .B_N(net344),
    .Y(_09689_));
 sg13g2_a21oi_1 _23302_ (.A1(net321),
    .A2(net7652),
    .Y(_09690_),
    .B1(_09689_));
 sg13g2_nor2_1 _23303_ (.A(net7644),
    .B(_09690_),
    .Y(_09691_));
 sg13g2_a21oi_1 _23304_ (.A1(net330),
    .A2(net7475),
    .Y(_09692_),
    .B1(_09691_));
 sg13g2_a21oi_1 _23305_ (.A1(_01992_),
    .A2(net7654),
    .Y(_09693_),
    .B1(_09689_));
 sg13g2_nor2_1 _23306_ (.A(net7645),
    .B(_09693_),
    .Y(_09694_));
 sg13g2_a21oi_1 _23307_ (.A1(_02000_),
    .A2(net7475),
    .Y(_09695_),
    .B1(_09694_));
 sg13g2_nor2_1 _23308_ (.A(net7664),
    .B(_09695_),
    .Y(_09696_));
 sg13g2_a221oi_1 _23309_ (.B2(net339),
    .C1(_09696_),
    .B1(_09381_),
    .A1(_02008_),
    .Y(_09697_),
    .A2(_09379_));
 sg13g2_o21ai_1 _23310_ (.B1(_09697_),
    .Y(_09698_),
    .A1(_09372_),
    .A2(_09692_));
 sg13g2_a21oi_1 _23311_ (.A1(net6973),
    .A2(_09410_),
    .Y(_09699_),
    .B1(_09413_));
 sg13g2_nand2_1 _23312_ (.Y(_09700_),
    .A(net6877),
    .B(_09699_));
 sg13g2_o21ai_1 _23313_ (.B1(_09700_),
    .Y(_09701_),
    .A1(net6877),
    .A2(_09430_));
 sg13g2_nand2_1 _23314_ (.Y(_09702_),
    .A(net6877),
    .B(_09423_));
 sg13g2_o21ai_1 _23315_ (.B1(_09702_),
    .Y(_09703_),
    .A1(net6877),
    .A2(_09486_));
 sg13g2_nor2_1 _23316_ (.A(net6850),
    .B(_09701_),
    .Y(_09704_));
 sg13g2_a21oi_1 _23317_ (.A1(net6850),
    .A2(_09703_),
    .Y(_09705_),
    .B1(_09704_));
 sg13g2_o21ai_1 _23318_ (.B1(_09642_),
    .Y(_09706_),
    .A1(net6798),
    .A2(_09705_));
 sg13g2_or2_1 _23319_ (.X(_09707_),
    .B(_09706_),
    .A(net6957));
 sg13g2_mux2_1 _23320_ (.A0(_09465_),
    .A1(_09478_),
    .S(net6974),
    .X(_09708_));
 sg13g2_mux2_1 _23321_ (.A0(_09644_),
    .A1(_09708_),
    .S(net6842),
    .X(_09709_));
 sg13g2_nand2_1 _23322_ (.Y(_09710_),
    .A(net6851),
    .B(_09709_));
 sg13g2_nand2_1 _23323_ (.Y(_09711_),
    .A(net6842),
    .B(_09646_));
 sg13g2_o21ai_1 _23324_ (.B1(_09711_),
    .Y(_09712_),
    .A1(net6842),
    .A2(_09523_));
 sg13g2_mux2_1 _23325_ (.A0(_01486_),
    .A1(_01521_),
    .S(net7771),
    .X(_09713_));
 sg13g2_o21ai_1 _23326_ (.B1(_09710_),
    .Y(_09714_),
    .A1(net6848),
    .A2(_09712_));
 sg13g2_nand3b_1 _23327_ (.B(_09416_),
    .C(net6851),
    .Y(_09715_),
    .A_N(_09525_));
 sg13g2_o21ai_1 _23328_ (.B1(_09518_),
    .Y(_09716_),
    .A1(net6845),
    .A2(net6875));
 sg13g2_a21oi_1 _23329_ (.A1(_09715_),
    .A2(_09716_),
    .Y(_09717_),
    .B1(net6803));
 sg13g2_nor3_1 _23330_ (.A(net7578),
    .B(net7563),
    .C(_09713_),
    .Y(_09718_));
 sg13g2_a21oi_1 _23331_ (.A1(net6803),
    .A2(_09714_),
    .Y(_09719_),
    .B1(_09717_));
 sg13g2_nand2_1 _23332_ (.Y(_09720_),
    .A(net6753),
    .B(_09719_));
 sg13g2_nand2_1 _23333_ (.Y(_09721_),
    .A(net7015),
    .B(net6966));
 sg13g2_o21ai_1 _23334_ (.B1(_09721_),
    .Y(_09722_),
    .A1(_03729_),
    .A2(net6966));
 sg13g2_mux2_1 _23335_ (.A0(_09448_),
    .A1(_09722_),
    .S(net6974),
    .X(_09723_));
 sg13g2_nand2_1 _23336_ (.Y(_09724_),
    .A(net6974),
    .B(_09436_));
 sg13g2_nand2_1 _23337_ (.Y(_09725_),
    .A(_03729_),
    .B(net6966));
 sg13g2_o21ai_1 _23338_ (.B1(_09725_),
    .Y(_09726_),
    .A1(net7015),
    .A2(net6968));
 sg13g2_o21ai_1 _23339_ (.B1(_09724_),
    .Y(_09727_),
    .A1(net6974),
    .A2(_09726_));
 sg13g2_mux2_1 _23340_ (.A0(_09723_),
    .A1(_09727_),
    .S(net6876),
    .X(_09728_));
 sg13g2_nand2_1 _23341_ (.Y(_09729_),
    .A(net6848),
    .B(_09728_));
 sg13g2_nand2_1 _23342_ (.Y(_09730_),
    .A(net6914),
    .B(_09435_));
 sg13g2_o21ai_1 _23343_ (.B1(_09730_),
    .Y(_09731_),
    .A1(net6914),
    .A2(_09462_));
 sg13g2_nor2_1 _23344_ (.A(net6974),
    .B(_09459_),
    .Y(_09732_));
 sg13g2_a21oi_1 _23345_ (.A1(net6974),
    .A2(_09468_),
    .Y(_09733_),
    .B1(_09732_));
 sg13g2_nand2_1 _23346_ (.Y(_09734_),
    .A(net6875),
    .B(_09733_));
 sg13g2_o21ai_1 _23347_ (.B1(_09734_),
    .Y(_09735_),
    .A1(net6875),
    .A2(_09731_));
 sg13g2_o21ai_1 _23348_ (.B1(_09729_),
    .Y(_09736_),
    .A1(net6848),
    .A2(_09735_));
 sg13g2_mux2_1 _23349_ (.A0(_09492_),
    .A1(_09502_),
    .S(net6916),
    .X(_09737_));
 sg13g2_nand2_1 _23350_ (.Y(_09738_),
    .A(net6915),
    .B(_09491_));
 sg13g2_o21ai_1 _23351_ (.B1(_09738_),
    .Y(_09739_),
    .A1(net6915),
    .A2(_09498_));
 sg13g2_mux2_1 _23352_ (.A0(_09446_),
    .A1(_09495_),
    .S(net6914),
    .X(_09740_));
 sg13g2_nor2_1 _23353_ (.A(net6875),
    .B(_09740_),
    .Y(_09741_));
 sg13g2_nand2_1 _23354_ (.Y(_09742_),
    .A(net6914),
    .B(_09444_));
 sg13g2_o21ai_1 _23355_ (.B1(_09742_),
    .Y(_09743_),
    .A1(net6914),
    .A2(_09451_));
 sg13g2_nor2_1 _23356_ (.A(_09416_),
    .B(_09743_),
    .Y(_09744_));
 sg13g2_mux2_1 _23357_ (.A0(_01557_),
    .A1(_01592_),
    .S(net7771),
    .X(_09745_));
 sg13g2_mux4_1 _23358_ (.S0(net6875),
    .A0(_09737_),
    .A1(_09739_),
    .A2(_09740_),
    .A3(_09743_),
    .S1(net6846),
    .X(_09746_));
 sg13g2_nor2_1 _23359_ (.A(_09403_),
    .B(_09409_),
    .Y(_09747_));
 sg13g2_nor2_1 _23360_ (.A(net7554),
    .B(_09745_),
    .Y(_09748_));
 sg13g2_mux2_1 _23361_ (.A0(_09736_),
    .A1(_09746_),
    .S(net6803),
    .X(_09749_));
 sg13g2_o21ai_1 _23362_ (.B1(_09720_),
    .Y(_09750_),
    .A1(net6753),
    .A2(_09749_));
 sg13g2_o21ai_1 _23363_ (.B1(_09707_),
    .Y(_09751_),
    .A1(net6962),
    .A2(_09750_));
 sg13g2_nand3_1 _23364_ (.B(net7024),
    .C(net6972),
    .A(net6899),
    .Y(_09752_));
 sg13g2_o21ai_1 _23365_ (.B1(_09752_),
    .Y(_09753_),
    .A1(net7024),
    .A2(net6906));
 sg13g2_a21oi_1 _23366_ (.A1(net7024),
    .A2(net6880),
    .Y(_09754_),
    .B1(net6899));
 sg13g2_a21oi_1 _23367_ (.A1(net6908),
    .A2(_09753_),
    .Y(_09755_),
    .B1(_09754_));
 sg13g2_a221oi_1 _23368_ (.B2(net7295),
    .C1(_09755_),
    .B1(_09751_),
    .A1(net6983),
    .Y(_09756_),
    .A2(net6628));
 sg13g2_or2_1 _23369_ (.X(_09757_),
    .B(_09756_),
    .A(net7382));
 sg13g2_a22oi_1 _23370_ (.Y(_09758_),
    .B1(net6871),
    .B2(_00174_),
    .A2(net6839),
    .A1(_00238_));
 sg13g2_a22oi_1 _23371_ (.Y(_09759_),
    .B1(net6871),
    .B2(_00145_),
    .A2(net6840),
    .A1(_00209_));
 sg13g2_a22oi_1 _23372_ (.Y(_09760_),
    .B1(net6673),
    .B2(_00246_),
    .A2(net6695),
    .A1(_00308_));
 sg13g2_inv_1 _23373_ (.Y(_09761_),
    .A(_09760_));
 sg13g2_a221oi_1 _23374_ (.B2(_00428_),
    .C1(_09761_),
    .B1(net6678),
    .A1(_00276_),
    .Y(_09762_),
    .A2(net6688));
 sg13g2_a221oi_1 _23375_ (.B2(_00503_),
    .C1(net6684),
    .B1(net6675),
    .A1(_00340_),
    .Y(_09763_),
    .A2(net6694));
 sg13g2_nand2_1 _23376_ (.Y(_09764_),
    .A(_00378_),
    .B(net6701));
 sg13g2_mux2_1 _23377_ (.A0(_01345_),
    .A1(_01381_),
    .S(net7770),
    .X(_09765_));
 sg13g2_nand3_1 _23378_ (.B(_09763_),
    .C(_09764_),
    .A(_09762_),
    .Y(_09766_));
 sg13g2_nand2b_1 _23379_ (.Y(_09767_),
    .B(_06850_),
    .A_N(_09758_));
 sg13g2_o21ai_1 _23380_ (.B1(_09767_),
    .Y(_09768_),
    .A1(_06865_),
    .A2(_09759_));
 sg13g2_a221oi_1 _23381_ (.B2(_09768_),
    .C1(_09766_),
    .B1(_09539_),
    .A1(net379),
    .Y(_09769_),
    .A2(net6780));
 sg13g2_nand2_1 _23382_ (.Y(_09770_),
    .A(_01639_),
    .B(_09671_));
 sg13g2_nor3_1 _23383_ (.A(net7578),
    .B(_08503_),
    .C(_09765_),
    .Y(_09771_));
 sg13g2_a21oi_1 _23384_ (.A1(_00108_),
    .A2(_08707_),
    .Y(_09772_),
    .B1(net6547));
 sg13g2_nand4_1 _23385_ (.B(_09769_),
    .C(_09770_),
    .A(_09757_),
    .Y(_09773_),
    .D(_09772_));
 sg13g2_o21ai_1 _23386_ (.B1(net6115),
    .Y(_09774_),
    .A1(net6552),
    .A2(_09698_));
 sg13g2_nand2_1 _23387_ (.Y(_09775_),
    .A(_01597_),
    .B(net6041));
 sg13g2_o21ai_1 _23388_ (.B1(_09775_),
    .Y(_09776_),
    .A1(net6041),
    .A2(net6030));
 sg13g2_nand3_1 _23389_ (.B(net7025),
    .C(net6972),
    .A(_13838_),
    .Y(_09777_));
 sg13g2_o21ai_1 _23390_ (.B1(_09777_),
    .Y(_09778_),
    .A1(net7025),
    .A2(net6907));
 sg13g2_nand2_1 _23391_ (.Y(_09779_),
    .A(net7025),
    .B(net6880));
 sg13g2_a22oi_1 _23392_ (.Y(_09780_),
    .B1(_09779_),
    .B2(net6948),
    .A2(_09778_),
    .A1(net6909));
 sg13g2_a21oi_1 _23393_ (.A1(net6982),
    .A2(net6637),
    .Y(_09781_),
    .B1(_09780_));
 sg13g2_nor2_1 _23394_ (.A(net6874),
    .B(_09470_),
    .Y(_09782_));
 sg13g2_a21oi_1 _23395_ (.A1(net6873),
    .A2(_09479_),
    .Y(_09783_),
    .B1(_09782_));
 sg13g2_nand2_1 _23396_ (.Y(_09784_),
    .A(net6849),
    .B(_09783_));
 sg13g2_o21ai_1 _23397_ (.B1(_09784_),
    .Y(_09785_),
    .A1(net6849),
    .A2(_09703_));
 sg13g2_a21oi_1 _23398_ (.A1(net6851),
    .A2(_09701_),
    .Y(_09786_),
    .B1(_09529_));
 sg13g2_nor2_1 _23399_ (.A(net6800),
    .B(_09786_),
    .Y(_09787_));
 sg13g2_mux2_1 _23400_ (.A0(_01416_),
    .A1(_01451_),
    .S(net7769),
    .X(_09788_));
 sg13g2_a21oi_1 _23401_ (.A1(net6800),
    .A2(_09785_),
    .Y(_09789_),
    .B1(_09787_));
 sg13g2_nor2_1 _23402_ (.A(net6872),
    .B(_09452_),
    .Y(_09790_));
 sg13g2_nor3_1 _23403_ (.A(net7578),
    .B(net7569),
    .C(_09788_),
    .Y(_09791_));
 sg13g2_a21oi_1 _23404_ (.A1(net6872),
    .A2(_09440_),
    .Y(_09792_),
    .B1(_09790_));
 sg13g2_nand2_1 _23405_ (.Y(_09793_),
    .A(net6849),
    .B(_09792_));
 sg13g2_nand2_1 _23406_ (.Y(_09794_),
    .A(net6872),
    .B(_09463_));
 sg13g2_o21ai_1 _23407_ (.B1(_09794_),
    .Y(_09795_),
    .A1(net6872),
    .A2(_09437_));
 sg13g2_o21ai_1 _23408_ (.B1(_09793_),
    .Y(_09796_),
    .A1(net6849),
    .A2(_09795_));
 sg13g2_nor2_1 _23409_ (.A(net6803),
    .B(_09796_),
    .Y(_09797_));
 sg13g2_nand2b_1 _23410_ (.Y(_09798_),
    .B(net6874),
    .A_N(_09493_));
 sg13g2_o21ai_1 _23411_ (.B1(_09798_),
    .Y(_09799_),
    .A1(net6874),
    .A2(_09505_));
 sg13g2_mux2_1 _23412_ (.A0(_09447_),
    .A1(_09499_),
    .S(net6843),
    .X(_09800_));
 sg13g2_nand2_1 _23413_ (.Y(_09801_),
    .A(net6849),
    .B(_09799_));
 sg13g2_o21ai_1 _23414_ (.B1(_09801_),
    .Y(_09802_),
    .A1(net6849),
    .A2(_09800_));
 sg13g2_a21oi_1 _23415_ (.A1(net6803),
    .A2(_09802_),
    .Y(_09803_),
    .B1(_09797_));
 sg13g2_nand2_1 _23416_ (.Y(_09804_),
    .A(net6753),
    .B(_09789_));
 sg13g2_o21ai_1 _23417_ (.B1(_09804_),
    .Y(_09805_),
    .A1(net6753),
    .A2(_09803_));
 sg13g2_nand2_1 _23418_ (.Y(_09806_),
    .A(net6956),
    .B(_09805_));
 sg13g2_nand2_1 _23419_ (.Y(_09807_),
    .A(net6875),
    .B(_09518_));
 sg13g2_o21ai_1 _23420_ (.B1(_09807_),
    .Y(_09808_),
    .A1(net6876),
    .A2(_09525_));
 sg13g2_nand2_1 _23421_ (.Y(_09809_),
    .A(net6844),
    .B(_09808_));
 sg13g2_inv_1 _23422_ (.Y(_09810_),
    .A(_09811_));
 sg13g2_o21ai_1 _23423_ (.B1(_09809_),
    .Y(_09811_),
    .A1(net6844),
    .A2(_09712_));
 sg13g2_o21ai_1 _23424_ (.B1(_09642_),
    .Y(_09812_),
    .A1(net6798),
    .A2(_09811_));
 sg13g2_a21oi_1 _23425_ (.A1(net6961),
    .A2(_09812_),
    .Y(_09813_),
    .B1(_08205_));
 sg13g2_nand2_1 _23426_ (.Y(_09814_),
    .A(_09806_),
    .B(_09813_));
 sg13g2_a21oi_1 _23427_ (.A1(_09781_),
    .A2(_09814_),
    .Y(_09815_),
    .B1(net7378));
 sg13g2_nor4_1 _23428_ (.A(_09718_),
    .B(_09748_),
    .C(_09771_),
    .D(_09791_),
    .Y(_09816_));
 sg13g2_a22oi_1 _23429_ (.Y(_09817_),
    .B1(net6871),
    .B2(_00169_),
    .A2(net6840),
    .A1(_00233_));
 sg13g2_a22oi_1 _23430_ (.Y(_09818_),
    .B1(net6871),
    .B2(_00144_),
    .A2(net6840),
    .A1(_00208_));
 sg13g2_a21oi_1 _23431_ (.A1(_00307_),
    .A2(net6695),
    .Y(_09819_),
    .B1(net6684));
 sg13g2_a22oi_1 _23432_ (.Y(_09820_),
    .B1(net6678),
    .B2(_00427_),
    .A2(net6692),
    .A1(_00339_));
 sg13g2_a22oi_1 _23433_ (.Y(_09821_),
    .B1(net6675),
    .B2(_00502_),
    .A2(net6779),
    .A1(net378));
 sg13g2_a22oi_1 _23434_ (.Y(_09822_),
    .B1(net6688),
    .B2(_00275_),
    .A2(net6701),
    .A1(_00377_));
 sg13g2_nand4_1 _23435_ (.B(_09820_),
    .C(_09821_),
    .A(_09819_),
    .Y(_09823_),
    .D(_09822_));
 sg13g2_nand2b_1 _23436_ (.Y(_09824_),
    .B(net6712),
    .A_N(_09817_));
 sg13g2_o21ai_1 _23437_ (.B1(_09824_),
    .Y(_09825_),
    .A1(net6652),
    .A2(_09818_));
 sg13g2_a21oi_1 _23438_ (.A1(net6796),
    .A2(_09825_),
    .Y(_09826_),
    .B1(_09823_));
 sg13g2_nand2_1 _23439_ (.Y(_09827_),
    .A(_01637_),
    .B(_09671_));
 sg13g2_a21oi_1 _23440_ (.A1(_00107_),
    .A2(net7088),
    .Y(_09828_),
    .B1(_09365_));
 sg13g2_nand3_1 _23441_ (.B(_09827_),
    .C(_09828_),
    .A(_09826_),
    .Y(_09829_));
 sg13g2_nand2_1 _23442_ (.Y(_09830_),
    .A(_01999_),
    .B(_09366_));
 sg13g2_nor2b_1 _23443_ (.A(net7650),
    .B_N(net343),
    .Y(_09831_));
 sg13g2_a21oi_1 _23444_ (.A1(_01991_),
    .A2(_01986_),
    .Y(_09832_),
    .B1(_09831_));
 sg13g2_o21ai_1 _23445_ (.B1(_09830_),
    .Y(_09833_),
    .A1(net7641),
    .A2(_09832_));
 sg13g2_nand2_1 _23446_ (.Y(_09834_),
    .A(net7628),
    .B(_09833_));
 sg13g2_nand2_1 _23447_ (.Y(_09835_),
    .A(net329),
    .B(_09366_));
 sg13g2_a21oi_1 _23448_ (.A1(net320),
    .A2(_01986_),
    .Y(_09836_),
    .B1(_09831_));
 sg13g2_o21ai_1 _23449_ (.B1(_09835_),
    .Y(_09837_),
    .A1(net7641),
    .A2(_09836_));
 sg13g2_nand2b_1 _23450_ (.Y(_09838_),
    .B(_09837_),
    .A_N(_09372_));
 sg13g2_a22oi_1 _23451_ (.Y(_09839_),
    .B1(_09381_),
    .B2(net337),
    .A2(_09379_),
    .A1(_02007_));
 sg13g2_nand4_1 _23452_ (.B(_09834_),
    .C(_09838_),
    .A(_09365_),
    .Y(_09840_),
    .D(_09839_));
 sg13g2_o21ai_1 _23453_ (.B1(_09840_),
    .Y(_09841_),
    .A1(_09815_),
    .A2(_09829_));
 sg13g2_nand2_1 _23454_ (.Y(_09842_),
    .A(_01596_),
    .B(net6034));
 sg13g2_o21ai_1 _23455_ (.B1(_09842_),
    .Y(_09843_),
    .A1(net6034),
    .A2(net6113));
 sg13g2_nor2b_1 _23456_ (.A(net7654),
    .B_N(net342),
    .Y(_09844_));
 sg13g2_a21oi_1 _23457_ (.A1(_01990_),
    .A2(net7654),
    .Y(_09845_),
    .B1(_09844_));
 sg13g2_nor2_1 _23458_ (.A(net7647),
    .B(_09845_),
    .Y(_09846_));
 sg13g2_a21oi_1 _23459_ (.A1(_01998_),
    .A2(net7476),
    .Y(_09847_),
    .B1(_09846_));
 sg13g2_nor2_1 _23460_ (.A(_00007_),
    .B(_09847_),
    .Y(_09848_));
 sg13g2_a21oi_1 _23461_ (.A1(net319),
    .A2(net7654),
    .Y(_09849_),
    .B1(_09844_));
 sg13g2_nor2_1 _23462_ (.A(net7644),
    .B(_09849_),
    .Y(_09850_));
 sg13g2_a21oi_1 _23463_ (.A1(net328),
    .A2(net7476),
    .Y(_09851_),
    .B1(_09850_));
 sg13g2_a221oi_1 _23464_ (.B2(net336),
    .C1(_09848_),
    .B1(_09381_),
    .A1(_02006_),
    .Y(_09852_),
    .A2(_09379_));
 sg13g2_o21ai_1 _23465_ (.B1(_09852_),
    .Y(_09853_),
    .A1(_09372_),
    .A2(_09851_));
 sg13g2_mux4_1 _23466_ (.S0(net7772),
    .A0(_01064_),
    .A1(_01099_),
    .A2(_01134_),
    .A3(_01169_),
    .S1(net7724),
    .X(_09854_));
 sg13g2_nand3_1 _23467_ (.B(net7026),
    .C(net6972),
    .A(net6951),
    .Y(_09855_));
 sg13g2_o21ai_1 _23468_ (.B1(_09855_),
    .Y(_09856_),
    .A1(net7026),
    .A2(net6907));
 sg13g2_inv_1 _23469_ (.Y(_09857_),
    .A(_09854_));
 sg13g2_nand2_1 _23470_ (.Y(_09858_),
    .A(net7026),
    .B(_09394_));
 sg13g2_a22oi_1 _23471_ (.Y(_09859_),
    .B1(_09858_),
    .B2(net6949),
    .A2(_09856_),
    .A1(net6909));
 sg13g2_or2_1 _23472_ (.X(_09860_),
    .B(_09859_),
    .A(_08239_));
 sg13g2_nand2_1 _23473_ (.Y(_09861_),
    .A(net6843),
    .B(_09733_));
 sg13g2_o21ai_1 _23474_ (.B1(_09861_),
    .Y(_09862_),
    .A1(net6843),
    .A2(_09708_));
 sg13g2_nand2_1 _23475_ (.Y(_09863_),
    .A(net6846),
    .B(_09647_));
 sg13g2_o21ai_1 _23476_ (.B1(_09863_),
    .Y(_09864_),
    .A1(net6845),
    .A2(_09862_));
 sg13g2_mux2_1 _23477_ (.A0(_09504_),
    .A1(_09507_),
    .S(net6913),
    .X(_09865_));
 sg13g2_mux2_1 _23478_ (.A0(_09737_),
    .A1(_09865_),
    .S(net6842),
    .X(_09866_));
 sg13g2_nand2_1 _23479_ (.Y(_09867_),
    .A(net6848),
    .B(_09866_));
 sg13g2_mux2_1 _23480_ (.A0(_09739_),
    .A1(_09740_),
    .S(net6875),
    .X(_09868_));
 sg13g2_nand2_1 _23481_ (.Y(_09869_),
    .A(net6845),
    .B(_09868_));
 sg13g2_nand3_1 _23482_ (.B(_09867_),
    .C(_09869_),
    .A(net6757),
    .Y(_09870_));
 sg13g2_o21ai_1 _23483_ (.B1(_09870_),
    .Y(_09871_),
    .A1(net6757),
    .A2(_09864_));
 sg13g2_nand2b_1 _23484_ (.Y(_09872_),
    .B(net6876),
    .A_N(_09723_));
 sg13g2_o21ai_1 _23485_ (.B1(_09872_),
    .Y(_09873_),
    .A1(net6876),
    .A2(_09743_));
 sg13g2_mux2_1 _23486_ (.A0(_09727_),
    .A1(_09731_),
    .S(net6876),
    .X(_09874_));
 sg13g2_nor2_1 _23487_ (.A(net6850),
    .B(_09874_),
    .Y(_09875_));
 sg13g2_a21oi_1 _23488_ (.A1(net6850),
    .A2(_09873_),
    .Y(_09876_),
    .B1(_09875_));
 sg13g2_nor2_1 _23489_ (.A(net6753),
    .B(_09876_),
    .Y(_09877_));
 sg13g2_a21oi_1 _23490_ (.A1(net6754),
    .A2(_09530_),
    .Y(_09878_),
    .B1(_09877_));
 sg13g2_nor2_1 _23491_ (.A(net6799),
    .B(_09878_),
    .Y(_09879_));
 sg13g2_a21oi_1 _23492_ (.A1(net6799),
    .A2(_09871_),
    .Y(_09880_),
    .B1(_09879_));
 sg13g2_a21oi_1 _23493_ (.A1(_09432_),
    .A2(_09520_),
    .Y(_09881_),
    .B1(_09521_));
 sg13g2_mux2_1 _23494_ (.A0(_09880_),
    .A1(_09881_),
    .S(net6964),
    .X(_09882_));
 sg13g2_a221oi_1 _23495_ (.B2(net7296),
    .C1(_09860_),
    .B1(_09882_),
    .A1(_08222_),
    .Y(_09883_),
    .A2(net6638));
 sg13g2_a221oi_1 _23496_ (.B2(_01636_),
    .C1(net7370),
    .B1(_09535_),
    .A1(_00106_),
    .Y(_09884_),
    .A2(_08739_));
 sg13g2_or2_1 _23497_ (.X(_09885_),
    .B(_09884_),
    .A(_09883_));
 sg13g2_a22oi_1 _23498_ (.Y(_09886_),
    .B1(net6871),
    .B2(_00158_),
    .A2(net6840),
    .A1(_00222_));
 sg13g2_nand2b_1 _23499_ (.Y(_09887_),
    .B(net6710),
    .A_N(_09886_));
 sg13g2_a22oi_1 _23500_ (.Y(_09888_),
    .B1(net6867),
    .B2(_00143_),
    .A2(net6841),
    .A1(_00207_));
 sg13g2_mux4_1 _23501_ (.S0(net7772),
    .A0(_01205_),
    .A1(_01240_),
    .A2(_01275_),
    .A3(_01310_),
    .S1(net7724),
    .X(_09889_));
 sg13g2_a22oi_1 _23502_ (.Y(_09890_),
    .B1(_09589_),
    .B2(_00501_),
    .A2(_09583_),
    .A1(_00338_));
 sg13g2_nand2_1 _23503_ (.Y(_09891_),
    .A(_00274_),
    .B(_09579_));
 sg13g2_a22oi_1 _23504_ (.Y(_09892_),
    .B1(_09582_),
    .B2(_00376_),
    .A2(_09577_),
    .A1(_00306_));
 sg13g2_nor2_1 _23505_ (.A(net7588),
    .B(_09889_),
    .Y(_09893_));
 sg13g2_a22oi_1 _23506_ (.Y(_09894_),
    .B1(_09586_),
    .B2(_00348_),
    .A2(_09575_),
    .A1(_00426_));
 sg13g2_nand4_1 _23507_ (.B(_09891_),
    .C(_09892_),
    .A(_09890_),
    .Y(_09895_),
    .D(_09894_));
 sg13g2_and2_1 _23508_ (.A(net377),
    .B(net6824),
    .X(_09896_));
 sg13g2_nand2b_1 _23509_ (.Y(_09897_),
    .B(net6707),
    .A_N(_09888_));
 sg13g2_a21oi_1 _23510_ (.A1(_09887_),
    .A2(_09897_),
    .Y(_09898_),
    .B1(_09538_));
 sg13g2_nor4_1 _23511_ (.A(_09585_),
    .B(_09895_),
    .C(_09896_),
    .D(_09898_),
    .Y(_09899_));
 sg13g2_a21oi_1 _23512_ (.A1(_08387_),
    .A2(_09857_),
    .Y(_09900_),
    .B1(_09893_));
 sg13g2_nand3_1 _23513_ (.B(_09885_),
    .C(_09899_),
    .A(net6550),
    .Y(_09901_));
 sg13g2_o21ai_1 _23514_ (.B1(_09901_),
    .Y(_09902_),
    .A1(net6551),
    .A2(_09853_));
 sg13g2_nand2_1 _23515_ (.Y(_09903_),
    .A(_01595_),
    .B(net6034));
 sg13g2_o21ai_1 _23516_ (.B1(_09903_),
    .Y(_09904_),
    .A1(net6034),
    .A2(net6026));
 sg13g2_nand2_1 _23517_ (.Y(_09905_),
    .A(_01594_),
    .B(net6040));
 sg13g2_o21ai_1 _23518_ (.B1(_09905_),
    .Y(_09906_),
    .A1(net6051),
    .A2(net6040));
 sg13g2_nor2b_1 _23519_ (.A(net7651),
    .B_N(net338),
    .Y(_09907_));
 sg13g2_a21oi_1 _23520_ (.A1(net317),
    .A2(net7651),
    .Y(_09908_),
    .B1(_09907_));
 sg13g2_nor2_1 _23521_ (.A(net7647),
    .B(_09908_),
    .Y(_09909_));
 sg13g2_a21oi_1 _23522_ (.A1(net325),
    .A2(net7476),
    .Y(_09910_),
    .B1(_09909_));
 sg13g2_a21oi_1 _23523_ (.A1(_01988_),
    .A2(net7651),
    .Y(_09911_),
    .B1(_09907_));
 sg13g2_nor2_1 _23524_ (.A(net7647),
    .B(_09911_),
    .Y(_09912_));
 sg13g2_a21oi_1 _23525_ (.A1(_01996_),
    .A2(net7476),
    .Y(_09913_),
    .B1(_09912_));
 sg13g2_nor2_1 _23526_ (.A(net7664),
    .B(_09913_),
    .Y(_09914_));
 sg13g2_a221oi_1 _23527_ (.B2(net334),
    .C1(_09914_),
    .B1(_09381_),
    .A1(_02004_),
    .Y(_09915_),
    .A2(_09379_));
 sg13g2_o21ai_1 _23528_ (.B1(_09915_),
    .Y(_09916_),
    .A1(_09372_),
    .A2(_09910_));
 sg13g2_nor2_1 _23529_ (.A(net6846),
    .B(_09735_),
    .Y(_09917_));
 sg13g2_a21oi_1 _23530_ (.A1(net6846),
    .A2(_09709_),
    .Y(_09918_),
    .B1(_09917_));
 sg13g2_nand2_1 _23531_ (.Y(_09919_),
    .A(net6802),
    .B(_09918_));
 sg13g2_o21ai_1 _23532_ (.B1(_09919_),
    .Y(_09920_),
    .A1(net6802),
    .A2(_09811_));
 sg13g2_nor2_1 _23533_ (.A(net6758),
    .B(_09920_),
    .Y(_09921_));
 sg13g2_nor3_1 _23534_ (.A(net6846),
    .B(_09741_),
    .C(_09744_),
    .Y(_09922_));
 sg13g2_a21oi_1 _23535_ (.A1(net6846),
    .A2(_09728_),
    .Y(_09923_),
    .B1(_09922_));
 sg13g2_nand3_1 _23536_ (.B(_09816_),
    .C(_09900_),
    .A(_09684_),
    .Y(_09924_));
 sg13g2_mux2_1 _23537_ (.A0(net7028),
    .A1(net7007),
    .S(net6965),
    .X(_09925_));
 sg13g2_mux2_1 _23538_ (.A0(_09509_),
    .A1(_09925_),
    .S(net6913),
    .X(_09926_));
 sg13g2_nor2_1 _23539_ (.A(_08641_),
    .B(net7077),
    .Y(_09927_));
 sg13g2_mux4_1 _23540_ (.S0(net6874),
    .A0(_09737_),
    .A1(_09739_),
    .A2(_09926_),
    .A3(_09865_),
    .S1(_09408_),
    .X(_09928_));
 sg13g2_nand2_1 _23541_ (.Y(_09929_),
    .A(net6802),
    .B(_09928_));
 sg13g2_o21ai_1 _23542_ (.B1(_09929_),
    .Y(_09930_),
    .A1(net6802),
    .A2(_09923_));
 sg13g2_a21oi_1 _23543_ (.A1(net6758),
    .A2(_09930_),
    .Y(_09931_),
    .B1(_09921_));
 sg13g2_nand2_1 _23544_ (.Y(_09932_),
    .A(net6954),
    .B(_09931_));
 sg13g2_nor2_1 _23545_ (.A(_09405_),
    .B(_09519_),
    .Y(_09933_));
 sg13g2_mux2_1 _23546_ (.A0(_09518_),
    .A1(_09701_),
    .S(_09747_),
    .X(_09934_));
 sg13g2_a21oi_1 _23547_ (.A1(net6758),
    .A2(_09934_),
    .Y(_09935_),
    .B1(_09933_));
 sg13g2_a21oi_1 _23548_ (.A1(net6961),
    .A2(_09935_),
    .Y(_09936_),
    .B1(_08205_));
 sg13g2_nand3_1 _23549_ (.B(net7028),
    .C(_09390_),
    .A(net6901),
    .Y(_09937_));
 sg13g2_o21ai_1 _23550_ (.B1(_09937_),
    .Y(_09938_),
    .A1(net7028),
    .A2(net6907));
 sg13g2_nand2_1 _23551_ (.Y(_09939_),
    .A(net7028),
    .B(net6880));
 sg13g2_a22oi_1 _23552_ (.Y(_09940_),
    .B1(_09939_),
    .B2(_10789_),
    .A2(_09938_),
    .A1(net6909));
 sg13g2_a221oi_1 _23553_ (.B2(_09936_),
    .C1(_09940_),
    .B1(_09932_),
    .A1(net6984),
    .Y(_09941_),
    .A2(net6640));
 sg13g2_a22oi_1 _23554_ (.Y(_09942_),
    .B1(net6867),
    .B2(_00136_),
    .A2(net6841),
    .A1(_00200_));
 sg13g2_a22oi_1 _23555_ (.Y(_09943_),
    .B1(net6867),
    .B2(_00141_),
    .A2(net6841),
    .A1(_00205_));
 sg13g2_inv_1 _23556_ (.Y(_09944_),
    .A(_09945_));
 sg13g2_nor2_1 _23557_ (.A(_09428_),
    .B(_09927_),
    .Y(_09945_));
 sg13g2_a22oi_1 _23558_ (.Y(_09946_),
    .B1(_09567_),
    .B2(_00334_),
    .A2(_09565_),
    .A1(_00346_));
 sg13g2_a22oi_1 _23559_ (.Y(_09947_),
    .B1(net6673),
    .B2(\cs_registers_i.debug_single_step_o ),
    .A2(net6679),
    .A1(_00422_));
 sg13g2_nand2_1 _23560_ (.Y(_09948_),
    .A(_09946_),
    .B(_09947_));
 sg13g2_a221oi_1 _23561_ (.B2(_00270_),
    .C1(_09948_),
    .B1(net6688),
    .A1(_00372_),
    .Y(_09949_),
    .A2(net6701));
 sg13g2_nor2_1 _23562_ (.A(_09546_),
    .B(_09562_),
    .Y(_09950_));
 sg13g2_a221oi_1 _23563_ (.B2(_00113_),
    .C1(_09950_),
    .B1(_09569_),
    .A1(_00302_),
    .Y(_09951_),
    .A2(net6695));
 sg13g2_a22oi_1 _23564_ (.Y(_09952_),
    .B1(net6675),
    .B2(_00497_),
    .A2(net6778),
    .A1(net373));
 sg13g2_nand3_1 _23565_ (.B(_09951_),
    .C(_09952_),
    .A(_09949_),
    .Y(_09953_));
 sg13g2_nand2b_1 _23566_ (.Y(_09954_),
    .B(net6712),
    .A_N(_09942_));
 sg13g2_o21ai_1 _23567_ (.B1(_09954_),
    .Y(_09955_),
    .A1(net6652),
    .A2(_09943_));
 sg13g2_a21oi_1 _23568_ (.A1(net6795),
    .A2(_09955_),
    .Y(_09956_),
    .B1(_09953_));
 sg13g2_nand2_1 _23569_ (.Y(_09957_),
    .A(_01634_),
    .B(_09671_));
 sg13g2_nand3_1 _23570_ (.B(_09956_),
    .C(_09957_),
    .A(net6549),
    .Y(_09958_));
 sg13g2_a21oi_1 _23571_ (.A1(_00100_),
    .A2(net7088),
    .Y(_09959_),
    .B1(_09958_));
 sg13g2_o21ai_1 _23572_ (.B1(_09959_),
    .Y(_09960_),
    .A1(net7382),
    .A2(_09941_));
 sg13g2_o21ai_1 _23573_ (.B1(_09960_),
    .Y(_09961_),
    .A1(net6552),
    .A2(_09916_));
 sg13g2_nand2_1 _23574_ (.Y(_09962_),
    .A(_01593_),
    .B(net6042));
 sg13g2_o21ai_1 _23575_ (.B1(_09962_),
    .Y(_09963_),
    .A1(net6042),
    .A2(net6020));
 sg13g2_mux2_1 _23576_ (.A0(_09792_),
    .A1(_09800_),
    .S(net6850),
    .X(_09964_));
 sg13g2_nor2_1 _23577_ (.A(net6803),
    .B(_09964_),
    .Y(_09965_));
 sg13g2_nor2_1 _23578_ (.A(net7006),
    .B(net6958),
    .Y(_09966_));
 sg13g2_a21oi_1 _23579_ (.A1(net7029),
    .A2(net6958),
    .Y(_09967_),
    .B1(_09966_));
 sg13g2_mux2_1 _23580_ (.A0(_09925_),
    .A1(_09967_),
    .S(net6913),
    .X(_09968_));
 sg13g2_mux2_1 _23581_ (.A0(_09510_),
    .A1(_09968_),
    .S(net6842),
    .X(_09969_));
 sg13g2_nand2_1 _23582_ (.Y(_09970_),
    .A(net6845),
    .B(_09799_));
 sg13g2_o21ai_1 _23583_ (.B1(_09970_),
    .Y(_09971_),
    .A1(net6845),
    .A2(_09969_));
 sg13g2_nand2b_1 _23584_ (.Y(_09972_),
    .B(net8001),
    .A_N(_01633_));
 sg13g2_a21oi_1 _23585_ (.A1(net6803),
    .A2(_09971_),
    .Y(_09973_),
    .B1(_09965_));
 sg13g2_nand2_1 _23586_ (.Y(_09974_),
    .A(net6757),
    .B(_09973_));
 sg13g2_nor2_1 _23587_ (.A(net6845),
    .B(_09795_),
    .Y(_09975_));
 sg13g2_a21oi_1 _23588_ (.A1(net6845),
    .A2(_09783_),
    .Y(_09976_),
    .B1(_09975_));
 sg13g2_nand2_1 _23589_ (.Y(_09977_),
    .A(net6800),
    .B(_09976_));
 sg13g2_o21ai_1 _23590_ (.B1(_09972_),
    .Y(_09978_),
    .A1(_01618_),
    .A2(net7480));
 sg13g2_o21ai_1 _23591_ (.B1(_09977_),
    .Y(_09979_),
    .A1(net6800),
    .A2(_09705_));
 sg13g2_o21ai_1 _23592_ (.B1(_09974_),
    .Y(_09980_),
    .A1(net6758),
    .A2(_09979_));
 sg13g2_nand2_1 _23593_ (.Y(_09981_),
    .A(_09416_),
    .B(_09747_));
 sg13g2_nand2_1 _23594_ (.Y(_09982_),
    .A(_09518_),
    .B(_09981_));
 sg13g2_o21ai_1 _23595_ (.B1(_09982_),
    .Y(_09983_),
    .A1(_09525_),
    .A2(_09981_));
 sg13g2_a21oi_1 _23596_ (.A1(net6758),
    .A2(_09983_),
    .Y(_09984_),
    .B1(_09933_));
 sg13g2_nand2_1 _23597_ (.Y(_09985_),
    .A(net6955),
    .B(_09980_));
 sg13g2_o21ai_1 _23598_ (.B1(_09985_),
    .Y(_09986_),
    .A1(net6955),
    .A2(_09984_));
 sg13g2_nand2_1 _23599_ (.Y(_09987_),
    .A(net7296),
    .B(_09986_));
 sg13g2_a22oi_1 _23600_ (.Y(_09988_),
    .B1(net6867),
    .B2(_00140_),
    .A2(net6841),
    .A1(_00204_));
 sg13g2_a22oi_1 _23601_ (.Y(_09989_),
    .B1(_09541_),
    .B2(_00125_),
    .A2(net6841),
    .A1(_00189_));
 sg13g2_and2_1 _23602_ (.A(net7029),
    .B(_09388_),
    .X(_09990_));
 sg13g2_nor3_1 _23603_ (.A(_09945_),
    .B(net7029),
    .C(_09389_),
    .Y(_09991_));
 sg13g2_o21ai_1 _23604_ (.B1(net6912),
    .Y(_09992_),
    .A1(_09990_),
    .A2(_09991_));
 sg13g2_o21ai_1 _23605_ (.B1(_09945_),
    .Y(_09993_),
    .A1(net7029),
    .A2(_09393_));
 sg13g2_and2_1 _23606_ (.A(_08222_),
    .B(net7365),
    .X(_09994_));
 sg13g2_o21ai_1 _23607_ (.B1(_01633_),
    .Y(_09995_),
    .A1(_08661_),
    .A2(_08753_));
 sg13g2_nand2_1 _23608_ (.Y(_09996_),
    .A(_09140_),
    .B(_09995_));
 sg13g2_a221oi_1 _23609_ (.B2(net6717),
    .C1(_09996_),
    .B1(_09994_),
    .A1(_09992_),
    .Y(_09997_),
    .A2(_09993_));
 sg13g2_nand2b_1 _23610_ (.Y(_09998_),
    .B(net6711),
    .A_N(_09989_));
 sg13g2_and2_1 _23611_ (.A(_00259_),
    .B(_09579_),
    .X(_09999_));
 sg13g2_a221oi_1 _23612_ (.B2(_00486_),
    .C1(_09999_),
    .B1(_09589_),
    .A1(_00323_),
    .Y(_10000_),
    .A2(_09583_));
 sg13g2_a22oi_1 _23613_ (.Y(_10001_),
    .B1(_09577_),
    .B2(_00291_),
    .A2(net6824),
    .A1(net362));
 sg13g2_a22oi_1 _23614_ (.Y(_10002_),
    .B1(_09586_),
    .B2(_00345_),
    .A2(_09575_),
    .A1(_00411_));
 sg13g2_a22oi_1 _23615_ (.Y(_10003_),
    .B1(_09675_),
    .B2(_06145_),
    .A2(_09582_),
    .A1(_00361_));
 sg13g2_nand4_1 _23616_ (.B(_10001_),
    .C(_10002_),
    .A(_10000_),
    .Y(_10004_),
    .D(_10003_));
 sg13g2_nand2b_1 _23617_ (.Y(_10005_),
    .B(net6707),
    .A_N(_09988_));
 sg13g2_a21oi_1 _23618_ (.A1(_09998_),
    .A2(_10005_),
    .Y(_10006_),
    .B1(_09538_));
 sg13g2_nor2_1 _23619_ (.A(_10004_),
    .B(_10006_),
    .Y(_10007_));
 sg13g2_mux4_1 _23620_ (.S0(net7918),
    .A0(_01486_),
    .A1(_01521_),
    .A2(_01557_),
    .A3(_01592_),
    .S1(net7830),
    .X(_10008_));
 sg13g2_nand4_1 _23621_ (.B(_09987_),
    .C(_09997_),
    .A(net6551),
    .Y(_10009_),
    .D(_10007_));
 sg13g2_nor2b_1 _23622_ (.A(net7655),
    .B_N(net327),
    .Y(_10010_));
 sg13g2_a21oi_1 _23623_ (.A1(net347),
    .A2(net7655),
    .Y(_10011_),
    .B1(_10010_));
 sg13g2_nor2_1 _23624_ (.A(net7644),
    .B(_10011_),
    .Y(_10012_));
 sg13g2_a21oi_1 _23625_ (.A1(net324),
    .A2(net7475),
    .Y(_10013_),
    .B1(_10012_));
 sg13g2_a21oi_1 _23626_ (.A1(_02011_),
    .A2(net7655),
    .Y(_10014_),
    .B1(_10010_));
 sg13g2_nor2_1 _23627_ (.A(net7645),
    .B(_10014_),
    .Y(_10015_));
 sg13g2_a21oi_1 _23628_ (.A1(_01995_),
    .A2(net7476),
    .Y(_10016_),
    .B1(_10015_));
 sg13g2_nor2_1 _23629_ (.A(net7664),
    .B(_10016_),
    .Y(_10017_));
 sg13g2_nand2_1 _23630_ (.Y(_10018_),
    .A(net7814),
    .B(_09150_));
 sg13g2_a221oi_1 _23631_ (.B2(net333),
    .C1(_10017_),
    .B1(_09381_),
    .A1(_02003_),
    .Y(_10019_),
    .A2(_09379_));
 sg13g2_nor2_1 _23632_ (.A(_10008_),
    .B(_10018_),
    .Y(_10020_));
 sg13g2_o21ai_1 _23633_ (.B1(_10019_),
    .Y(_10021_),
    .A1(_09372_),
    .A2(_10013_));
 sg13g2_o21ai_1 _23634_ (.B1(net6394),
    .Y(_10022_),
    .A1(net6552),
    .A2(_10021_));
 sg13g2_nand2_1 _23635_ (.Y(_10023_),
    .A(_01592_),
    .B(net6041));
 sg13g2_o21ai_1 _23636_ (.B1(_10023_),
    .Y(_10024_),
    .A1(net6041),
    .A2(net6106));
 sg13g2_nand2_1 _23637_ (.Y(_10025_),
    .A(_00078_),
    .B(_08739_));
 sg13g2_a21oi_1 _23638_ (.A1(_01632_),
    .A2(_09535_),
    .Y(_10026_),
    .B1(_08242_));
 sg13g2_nand2_1 _23639_ (.Y(_10027_),
    .A(_10025_),
    .B(_10026_));
 sg13g2_nor2_1 _23640_ (.A(net6848),
    .B(_09862_),
    .Y(_10028_));
 sg13g2_a21oi_1 _23641_ (.A1(net6848),
    .A2(_09874_),
    .Y(_10029_),
    .B1(_10028_));
 sg13g2_nand2_1 _23642_ (.Y(_10030_),
    .A(net6800),
    .B(_10029_));
 sg13g2_o21ai_1 _23643_ (.B1(_10030_),
    .Y(_10031_),
    .A1(net6801),
    .A2(_09649_));
 sg13g2_nor2_1 _23644_ (.A(net6756),
    .B(_10031_),
    .Y(_10032_));
 sg13g2_nand2_1 _23645_ (.Y(_10033_),
    .A(net6847),
    .B(_09866_));
 sg13g2_nor2_1 _23646_ (.A(_03812_),
    .B(net6958),
    .Y(_10034_));
 sg13g2_nor2_1 _23647_ (.A(net7072),
    .B(net6964),
    .Y(_10035_));
 sg13g2_nor3_1 _23648_ (.A(net6973),
    .B(_10034_),
    .C(_10035_),
    .Y(_10036_));
 sg13g2_a21oi_1 _23649_ (.A1(net6973),
    .A2(_09967_),
    .Y(_10037_),
    .B1(_10036_));
 sg13g2_nor2_1 _23650_ (.A(net6877),
    .B(_10037_),
    .Y(_10038_));
 sg13g2_a21oi_1 _23651_ (.A1(net6877),
    .A2(_09926_),
    .Y(_10039_),
    .B1(_10038_));
 sg13g2_o21ai_1 _23652_ (.B1(_10033_),
    .Y(_10040_),
    .A1(_09409_),
    .A2(_10039_));
 sg13g2_nor2_1 _23653_ (.A(net6850),
    .B(_09873_),
    .Y(_10041_));
 sg13g2_a21oi_1 _23654_ (.A1(net6848),
    .A2(_09868_),
    .Y(_10042_),
    .B1(_10041_));
 sg13g2_nand2_1 _23655_ (.Y(_10043_),
    .A(net6802),
    .B(_10040_));
 sg13g2_o21ai_1 _23656_ (.B1(_10043_),
    .Y(_10044_),
    .A1(net6802),
    .A2(_10042_));
 sg13g2_a21oi_1 _23657_ (.A1(net6756),
    .A2(_10044_),
    .Y(_10045_),
    .B1(_10032_));
 sg13g2_o21ai_1 _23658_ (.B1(_09410_),
    .Y(_10046_),
    .A1(net6953),
    .A2(_06800_));
 sg13g2_nand2b_1 _23659_ (.Y(_10047_),
    .B(_10046_),
    .A_N(_09413_));
 sg13g2_nor2_1 _23660_ (.A(_09405_),
    .B(_09518_),
    .Y(_10048_));
 sg13g2_o21ai_1 _23661_ (.B1(net6964),
    .Y(_10049_),
    .A1(_10047_),
    .A2(_10048_));
 sg13g2_nand2_1 _23662_ (.Y(_10050_),
    .A(net7294),
    .B(_10049_));
 sg13g2_a21oi_1 _23663_ (.A1(net6958),
    .A2(_10045_),
    .Y(_10051_),
    .B1(_10050_));
 sg13g2_and2_1 _23664_ (.A(net6982),
    .B(net6743),
    .X(_10052_));
 sg13g2_nand3_1 _23665_ (.B(net7072),
    .C(net6972),
    .A(net6977),
    .Y(_10053_));
 sg13g2_o21ai_1 _23666_ (.B1(_10053_),
    .Y(_10054_),
    .A1(net7072),
    .A2(net6907));
 sg13g2_nand2_1 _23667_ (.Y(_10055_),
    .A(net7072),
    .B(net6880));
 sg13g2_a22oi_1 _23668_ (.Y(_10056_),
    .B1(_10055_),
    .B2(net6913),
    .A2(_10054_),
    .A1(net6909));
 sg13g2_nor4_1 _23669_ (.A(net7378),
    .B(_10051_),
    .C(_10052_),
    .D(_10056_),
    .Y(_10057_));
 sg13g2_o21ai_1 _23670_ (.B1(_10057_),
    .Y(_10058_),
    .A1(_08014_),
    .A2(net6056));
 sg13g2_nand3_1 _23671_ (.B(_10027_),
    .C(_10058_),
    .A(_06770_),
    .Y(_10059_));
 sg13g2_a22oi_1 _23672_ (.Y(_10060_),
    .B1(_09541_),
    .B2(_00114_),
    .A2(net6837),
    .A1(_00178_));
 sg13g2_nand2b_1 _23673_ (.Y(_10061_),
    .B(net6711),
    .A_N(_10060_));
 sg13g2_a22oi_1 _23674_ (.Y(_10062_),
    .B1(net6868),
    .B2(_00139_),
    .A2(net6841),
    .A1(_00203_));
 sg13g2_nor4_1 _23675_ (.A(_08874_),
    .B(_06810_),
    .C(_06814_),
    .D(_09546_),
    .Y(_10063_));
 sg13g2_mux4_1 _23676_ (.S0(net7864),
    .A0(_01345_),
    .A1(_01381_),
    .A2(_01416_),
    .A3(_01451_),
    .S1(net7830),
    .X(_10064_));
 sg13g2_nor3_1 _23677_ (.A(net6900),
    .B(_09546_),
    .C(_09561_),
    .Y(_10065_));
 sg13g2_nor3_1 _23678_ (.A(net7814),
    .B(net7490),
    .C(_10064_),
    .Y(_10066_));
 sg13g2_a22oi_1 _23679_ (.Y(_10067_),
    .B1(_09583_),
    .B2(_00312_),
    .A2(net6824),
    .A1(net351));
 sg13g2_a22oi_1 _23680_ (.Y(_10068_),
    .B1(_09585_),
    .B2(_00112_),
    .A2(_09575_),
    .A1(_00400_));
 sg13g2_a22oi_1 _23681_ (.Y(_10069_),
    .B1(_09675_),
    .B2(_06149_),
    .A2(_09586_),
    .A1(_00344_));
 sg13g2_a22oi_1 _23682_ (.Y(_10070_),
    .B1(_09589_),
    .B2(_00475_),
    .A2(_09577_),
    .A1(_00280_));
 sg13g2_nand4_1 _23683_ (.B(_10068_),
    .C(_10069_),
    .A(_10067_),
    .Y(_10071_),
    .D(_10070_));
 sg13g2_nor4_1 _23684_ (.A(_08874_),
    .B(_06810_),
    .C(_06814_),
    .D(_09590_),
    .Y(_10072_));
 sg13g2_and2_1 _23685_ (.A(_00350_),
    .B(_09582_),
    .X(_10073_));
 sg13g2_nand2b_1 _23686_ (.Y(_10074_),
    .B(net6707),
    .A_N(_10062_));
 sg13g2_a21oi_1 _23687_ (.A1(_10061_),
    .A2(_10074_),
    .Y(_10075_),
    .B1(_09538_));
 sg13g2_nor4_1 _23688_ (.A(_10071_),
    .B(_10072_),
    .C(_10073_),
    .D(_10075_),
    .Y(_10076_));
 sg13g2_nand3_1 _23689_ (.B(_10059_),
    .C(_10076_),
    .A(net6551),
    .Y(_10077_));
 sg13g2_nor2b_1 _23690_ (.A(net7650),
    .B_N(net316),
    .Y(_10078_));
 sg13g2_a21oi_1 _23691_ (.A1(_02010_),
    .A2(net7649),
    .Y(_10079_),
    .B1(_10078_));
 sg13g2_nor2_1 _23692_ (.A(net7642),
    .B(_10079_),
    .Y(_10080_));
 sg13g2_a21oi_1 _23693_ (.A1(_01994_),
    .A2(_09366_),
    .Y(_10081_),
    .B1(_10080_));
 sg13g2_a21oi_1 _23694_ (.A1(net346),
    .A2(net7649),
    .Y(_10082_),
    .B1(_10078_));
 sg13g2_nor2_1 _23695_ (.A(net7642),
    .B(_10082_),
    .Y(_10083_));
 sg13g2_a21oi_1 _23696_ (.A1(net323),
    .A2(_09366_),
    .Y(_10084_),
    .B1(_10083_));
 sg13g2_nor2_1 _23697_ (.A(_09372_),
    .B(_10084_),
    .Y(_10085_));
 sg13g2_a221oi_1 _23698_ (.B2(net332),
    .C1(_10085_),
    .B1(_09381_),
    .A1(_02002_),
    .Y(_10086_),
    .A2(_09379_));
 sg13g2_o21ai_1 _23699_ (.B1(_10086_),
    .Y(_10087_),
    .A1(_00007_),
    .A2(_10081_));
 sg13g2_o21ai_1 _23700_ (.B1(_10077_),
    .Y(_10088_),
    .A1(_09364_),
    .A2(_10087_));
 sg13g2_nand2_1 _23701_ (.Y(_10089_),
    .A(_01591_),
    .B(net6038));
 sg13g2_o21ai_1 _23702_ (.B1(_10089_),
    .Y(_10090_),
    .A1(net6038),
    .A2(net5867));
 sg13g2_nor2_1 _23703_ (.A(_01915_),
    .B(_09373_),
    .Y(_10091_));
 sg13g2_nand2_1 _23704_ (.Y(_10092_),
    .A(_08510_),
    .B(_01888_));
 sg13g2_nand4_1 _23705_ (.B(net6466),
    .C(_09679_),
    .A(net7669),
    .Y(_10093_),
    .D(_10091_));
 sg13g2_nor2_1 _23706_ (.A(_09607_),
    .B(_10092_),
    .Y(_10094_));
 sg13g2_nand2_1 _23707_ (.Y(_10095_),
    .A(net7474),
    .B(_10094_));
 sg13g2_nand2_1 _23708_ (.Y(_10096_),
    .A(_01590_),
    .B(net6387));
 sg13g2_mux4_1 _23709_ (.S0(net7656),
    .A0(net345),
    .A1(net322),
    .A2(net331),
    .A3(net340),
    .S1(_01987_),
    .X(_10097_));
 sg13g2_and3_1 _23710_ (.X(_10098_),
    .A(_01981_),
    .B(\load_store_unit_i.data_sign_ext_q ),
    .C(_10097_));
 sg13g2_mux4_1 _23711_ (.S0(net7656),
    .A0(net322),
    .A1(net331),
    .A2(net340),
    .A3(net345),
    .S1(net7648),
    .X(_10099_));
 sg13g2_a21o_1 _23712_ (.A2(_10099_),
    .A1(net7661),
    .B1(_10098_),
    .X(_10100_));
 sg13g2_a21oi_1 _23713_ (.A1(\load_store_unit_i.data_sign_ext_q ),
    .A2(_10100_),
    .Y(_10101_),
    .B1(net6552));
 sg13g2_inv_1 _23714_ (.Y(_10102_),
    .A(_10103_));
 sg13g2_mux4_1 _23715_ (.S0(net7648),
    .A0(net340),
    .A1(net322),
    .A2(net345),
    .A3(net331),
    .S1(net7651),
    .X(_10103_));
 sg13g2_o21ai_1 _23716_ (.B1(_10101_),
    .Y(_10104_),
    .A1(net7664),
    .A2(_10102_));
 sg13g2_nor2_1 _23717_ (.A(_03812_),
    .B(net6905),
    .Y(_10105_));
 sg13g2_nor3_1 _23718_ (.A(_03611_),
    .B(_03811_),
    .C(_09389_),
    .Y(_10106_));
 sg13g2_o21ai_1 _23719_ (.B1(net6912),
    .Y(_10107_),
    .A1(_10105_),
    .A2(_10106_));
 sg13g2_o21ai_1 _23720_ (.B1(_03611_),
    .Y(_10108_),
    .A1(_03811_),
    .A2(_09393_));
 sg13g2_a221oi_1 _23721_ (.B2(_10108_),
    .C1(net7378),
    .B1(_10107_),
    .A1(net6982),
    .Y(_10109_),
    .A2(net6567));
 sg13g2_nand2_1 _23722_ (.Y(_10110_),
    .A(net6964),
    .B(_10045_));
 sg13g2_o21ai_1 _23723_ (.B1(net6958),
    .Y(_10111_),
    .A1(_10047_),
    .A2(_10048_));
 sg13g2_nand3_1 _23724_ (.B(_10110_),
    .C(_10111_),
    .A(net7294),
    .Y(_10112_));
 sg13g2_a22oi_1 _23725_ (.Y(_10113_),
    .B1(_10109_),
    .B2(_10112_),
    .A2(_08716_),
    .A1(net7379));
 sg13g2_a22oi_1 _23726_ (.Y(_10114_),
    .B1(net6862),
    .B2(_00138_),
    .A2(net6832),
    .A1(_00202_));
 sg13g2_nand2b_1 _23727_ (.Y(_10115_),
    .B(net6709),
    .A_N(_10114_));
 sg13g2_a22oi_1 _23728_ (.Y(_10116_),
    .B1(net6862),
    .B2(_00173_),
    .A2(net6832),
    .A1(_00237_));
 sg13g2_o21ai_1 _23729_ (.B1(_10115_),
    .Y(_10117_),
    .A1(_06865_),
    .A2(_10116_));
 sg13g2_a22oi_1 _23730_ (.Y(_10118_),
    .B1(net6690),
    .B2(_00336_),
    .A2(net6696),
    .A1(_00304_));
 sg13g2_inv_1 _23731_ (.Y(_10119_),
    .A(_10118_));
 sg13g2_a221oi_1 _23732_ (.B2(_00528_),
    .C1(_10119_),
    .B1(net6672),
    .A1(_00424_),
    .Y(_10120_),
    .A2(net6679));
 sg13g2_a22oi_1 _23733_ (.Y(_10121_),
    .B1(net6689),
    .B2(_00272_),
    .A2(net6702),
    .A1(_00374_));
 sg13g2_a221oi_1 _23734_ (.B2(_00499_),
    .C1(net6685),
    .B1(net6676),
    .A1(_00349_),
    .Y(_10122_),
    .A2(_09565_));
 sg13g2_nand2_1 _23735_ (.Y(_10123_),
    .A(net375),
    .B(net6778));
 sg13g2_nand4_1 _23736_ (.B(_10121_),
    .C(_10122_),
    .A(_10120_),
    .Y(_10124_),
    .D(_10123_));
 sg13g2_a21oi_1 _23737_ (.A1(_09539_),
    .A2(_10117_),
    .Y(_10125_),
    .B1(_10124_));
 sg13g2_nand2_1 _23738_ (.Y(_10126_),
    .A(net6549),
    .B(_10125_));
 sg13g2_o21ai_1 _23739_ (.B1(_10104_),
    .Y(_10127_),
    .A1(_10113_),
    .A2(_10126_));
 sg13g2_nand3_1 _23740_ (.B(net7081),
    .C(net6385),
    .A(net5970),
    .Y(_10128_));
 sg13g2_nand2_1 _23741_ (.Y(_10129_),
    .A(net6017),
    .B(_10128_));
 sg13g2_and2_1 _23742_ (.A(net7084),
    .B(net6385),
    .X(_10130_));
 sg13g2_mux4_1 _23743_ (.S0(net7918),
    .A0(_01205_),
    .A1(_01240_),
    .A2(_01275_),
    .A3(_01310_),
    .S1(net7830),
    .X(_10131_));
 sg13g2_a21oi_1 _23744_ (.A1(_00102_),
    .A2(_10130_),
    .Y(_10132_),
    .B1(_10129_));
 sg13g2_o21ai_1 _23745_ (.B1(_10096_),
    .Y(_10133_),
    .A1(net6387),
    .A2(net5863));
 sg13g2_nand2_1 _23746_ (.Y(_10134_),
    .A(_01589_),
    .B(net6392));
 sg13g2_nor2_1 _23747_ (.A(net6955),
    .B(_09980_),
    .Y(_10135_));
 sg13g2_a21oi_1 _23748_ (.A1(net6955),
    .A2(_09984_),
    .Y(_10136_),
    .B1(_10135_));
 sg13g2_nand2_1 _23749_ (.Y(_10137_),
    .A(net7293),
    .B(_10136_));
 sg13g2_a22oi_1 _23750_ (.Y(_10138_),
    .B1(net6862),
    .B2(_00137_),
    .A2(net6832),
    .A1(_00201_));
 sg13g2_nand2b_1 _23751_ (.Y(_10139_),
    .B(net6709),
    .A_N(_10138_));
 sg13g2_a22oi_1 _23752_ (.Y(_10140_),
    .B1(net6862),
    .B2(_00172_),
    .A2(net6832),
    .A1(_00236_));
 sg13g2_o21ai_1 _23753_ (.B1(_10139_),
    .Y(_10141_),
    .A1(_06865_),
    .A2(_10140_));
 sg13g2_a21oi_1 _23754_ (.A1(_00303_),
    .A2(net6696),
    .Y(_10142_),
    .B1(_09661_));
 sg13g2_a22oi_1 _23755_ (.Y(_10143_),
    .B1(net6680),
    .B2(_00423_),
    .A2(net6691),
    .A1(_00335_));
 sg13g2_a22oi_1 _23756_ (.Y(_10144_),
    .B1(net6674),
    .B2(_00498_),
    .A2(net6778),
    .A1(net374));
 sg13g2_nand3_1 _23757_ (.B(_10143_),
    .C(_10144_),
    .A(_10142_),
    .Y(_10145_));
 sg13g2_a221oi_1 _23758_ (.B2(_00527_),
    .C1(_10145_),
    .B1(net6671),
    .A1(_00373_),
    .Y(_10146_),
    .A2(net6699));
 sg13g2_or2_1 _23759_ (.X(_10147_),
    .B(_09950_),
    .A(_09569_));
 sg13g2_a21oi_1 _23760_ (.A1(_00387_),
    .A2(net6705),
    .Y(_10148_),
    .B1(_10147_));
 sg13g2_a22oi_1 _23761_ (.Y(_10149_),
    .B1(net6686),
    .B2(_00271_),
    .A2(net6704),
    .A1(net424));
 sg13g2_nand3_1 _23762_ (.B(_10148_),
    .C(_10149_),
    .A(_10146_),
    .Y(_10150_));
 sg13g2_a21oi_1 _23763_ (.A1(_09539_),
    .A2(_10141_),
    .Y(_10151_),
    .B1(_10150_));
 sg13g2_nand3b_1 _23764_ (.B(net7006),
    .C(net6970),
    .Y(_10152_),
    .A_N(_03539_));
 sg13g2_o21ai_1 _23765_ (.B1(_10152_),
    .Y(_10153_),
    .A1(net7006),
    .A2(net6904));
 sg13g2_nand2_1 _23766_ (.Y(_10154_),
    .A(net7006),
    .B(net6878));
 sg13g2_a22oi_1 _23767_ (.Y(_10155_),
    .B1(_10154_),
    .B2(_03539_),
    .A2(_10153_),
    .A1(net6910));
 sg13g2_a21oi_1 _23768_ (.A1(_01665_),
    .A2(net7288),
    .Y(_10156_),
    .B1(_10155_));
 sg13g2_a21oi_1 _23769_ (.A1(net6570),
    .A2(net6902),
    .Y(_10157_),
    .B1(net6547));
 sg13g2_nand4_1 _23770_ (.B(_10151_),
    .C(_10156_),
    .A(_10137_),
    .Y(_10158_),
    .D(_10157_));
 sg13g2_a221oi_1 _23771_ (.B2(net6057),
    .C1(_10158_),
    .B1(net7081),
    .A1(_00101_),
    .Y(_10159_),
    .A2(net7084));
 sg13g2_inv_1 _23772_ (.Y(_10160_),
    .A(_10161_));
 sg13g2_mux4_1 _23773_ (.S0(net7645),
    .A0(net339),
    .A1(net321),
    .A2(net344),
    .A3(net330),
    .S1(net7653),
    .X(_10161_));
 sg13g2_o21ai_1 _23774_ (.B1(net6463),
    .Y(_10162_),
    .A1(net7662),
    .A2(_10160_));
 sg13g2_nand2b_1 _23775_ (.Y(_10163_),
    .B(net6384),
    .A_N(net6392));
 sg13g2_mux4_1 _23776_ (.S0(net7918),
    .A0(_01064_),
    .A1(_01099_),
    .A2(_01134_),
    .A3(_01169_),
    .S1(net7830),
    .X(_10164_));
 sg13g2_inv_1 _23777_ (.Y(_10165_),
    .A(\id_stage_i.controller_i.instr_fetch_err_i ));
 sg13g2_o21ai_1 _23778_ (.B1(_10134_),
    .Y(_10166_),
    .A1(net5858),
    .A2(_10163_));
 sg13g2_nand2_1 _23779_ (.Y(_10167_),
    .A(_01588_),
    .B(net6050));
 sg13g2_o21ai_1 _23780_ (.B1(_10167_),
    .Y(_10168_),
    .A1(net6050),
    .A2(net6022));
 sg13g2_nand2_1 _23781_ (.Y(_10169_),
    .A(_01587_),
    .B(net6386));
 sg13g2_nand3b_1 _23782_ (.B(net7007),
    .C(net6970),
    .Y(_10170_),
    .A_N(_03474_));
 sg13g2_o21ai_1 _23783_ (.B1(_10170_),
    .Y(_10171_),
    .A1(net7007),
    .A2(net6904));
 sg13g2_nand2_1 _23784_ (.Y(_10172_),
    .A(net7007),
    .B(net6878));
 sg13g2_a22oi_1 _23785_ (.Y(_10173_),
    .B1(_10172_),
    .B2(_03474_),
    .A2(_10171_),
    .A1(net6910));
 sg13g2_and2_1 _23786_ (.A(net6954),
    .B(_09935_),
    .X(_10174_));
 sg13g2_a21oi_1 _23787_ (.A1(net6963),
    .A2(_09931_),
    .Y(_10175_),
    .B1(_10174_));
 sg13g2_a221oi_1 _23788_ (.B2(net7295),
    .C1(_10173_),
    .B1(_10175_),
    .A1(net6983),
    .Y(_10176_),
    .A2(net6571));
 sg13g2_a21oi_1 _23789_ (.A1(net7923),
    .A2(_01664_),
    .Y(_10177_),
    .B1(net7367));
 sg13g2_a21o_1 _23790_ (.A2(_10176_),
    .A1(net7367),
    .B1(_10177_),
    .X(_10178_));
 sg13g2_nor2_1 _23791_ (.A(net7815),
    .B(net7835),
    .Y(_10179_));
 sg13g2_a22oi_1 _23792_ (.Y(_10180_),
    .B1(net6704),
    .B2(net423),
    .A2(net6705),
    .A1(_00386_));
 sg13g2_nand2_1 _23793_ (.Y(_10181_),
    .A(_00371_),
    .B(net6699));
 sg13g2_or2_1 _23794_ (.X(_10182_),
    .B(_01893_),
    .A(_01894_));
 sg13g2_a21oi_1 _23795_ (.A1(_00301_),
    .A2(net6696),
    .Y(_10183_),
    .B1(net6683));
 sg13g2_a22oi_1 _23796_ (.Y(_10184_),
    .B1(net6680),
    .B2(_00421_),
    .A2(net6691),
    .A1(_00333_));
 sg13g2_a22oi_1 _23797_ (.Y(_10185_),
    .B1(net6676),
    .B2(_00496_),
    .A2(net6780),
    .A1(net372));
 sg13g2_nand3_1 _23798_ (.B(_10184_),
    .C(_10185_),
    .A(_10183_),
    .Y(_10186_));
 sg13g2_a221oi_1 _23799_ (.B2(_00526_),
    .C1(_10186_),
    .B1(net6671),
    .A1(_00269_),
    .Y(_10187_),
    .A2(net6686));
 sg13g2_nand3_1 _23800_ (.B(_10181_),
    .C(_10187_),
    .A(_10180_),
    .Y(_10188_));
 sg13g2_nor2b_1 _23801_ (.A(net7815),
    .B_N(net7835),
    .Y(_10189_));
 sg13g2_a22oi_1 _23802_ (.Y(_10190_),
    .B1(net6862),
    .B2(_00171_),
    .A2(net6832),
    .A1(_00235_));
 sg13g2_nand2b_1 _23803_ (.Y(_10191_),
    .B(_01893_),
    .A_N(_01894_));
 sg13g2_a22oi_1 _23804_ (.Y(_10192_),
    .B1(net6862),
    .B2(_00135_),
    .A2(net6837),
    .A1(_00199_));
 sg13g2_nand2b_1 _23805_ (.Y(_10193_),
    .B(net6713),
    .A_N(_10192_));
 sg13g2_o21ai_1 _23806_ (.B1(_10193_),
    .Y(_10194_),
    .A1(_06865_),
    .A2(_10190_));
 sg13g2_a21oi_1 _23807_ (.A1(_09539_),
    .A2(_10194_),
    .Y(_10195_),
    .B1(_10188_));
 sg13g2_nand2_1 _23808_ (.Y(_10196_),
    .A(net6058),
    .B(_08742_));
 sg13g2_nand4_1 _23809_ (.B(_10178_),
    .C(_10195_),
    .A(net6548),
    .Y(_10197_),
    .D(_10196_));
 sg13g2_mux2_1 _23810_ (.A0(_10131_),
    .A1(_10164_),
    .S(net7485),
    .X(_10198_));
 sg13g2_nor2_1 _23811_ (.A(net7500),
    .B(_10198_),
    .Y(_10199_));
 sg13g2_nor3_1 _23812_ (.A(_10020_),
    .B(_10066_),
    .C(_10199_),
    .Y(_10200_));
 sg13g2_a21oi_1 _23813_ (.A1(_00099_),
    .A2(net7088),
    .Y(_10201_),
    .B1(_10197_));
 sg13g2_mux4_1 _23814_ (.S0(net7641),
    .A0(net337),
    .A1(net320),
    .A2(net343),
    .A3(net329),
    .S1(net7649),
    .X(_10202_));
 sg13g2_nand2_1 _23815_ (.Y(_10203_),
    .A(net7628),
    .B(_10202_));
 sg13g2_a21o_1 _23816_ (.A2(_10203_),
    .A1(net6465),
    .B1(net5852),
    .X(_10204_));
 sg13g2_o21ai_1 _23817_ (.B1(_10169_),
    .Y(_10205_),
    .A1(net6018),
    .A2(net5808));
 sg13g2_nand2_1 _23818_ (.Y(_10206_),
    .A(_01586_),
    .B(net6392));
 sg13g2_inv_1 _23819_ (.Y(_10207_),
    .A(_10208_));
 sg13g2_mux4_1 _23820_ (.S0(net7646),
    .A0(net336),
    .A1(net319),
    .A2(net342),
    .A3(net328),
    .S1(net7653),
    .X(_10208_));
 sg13g2_o21ai_1 _23821_ (.B1(net6464),
    .Y(_10209_),
    .A1(net7662),
    .A2(_10207_));
 sg13g2_nand2_1 _23822_ (.Y(_10210_),
    .A(net6956),
    .B(_09531_));
 sg13g2_o21ai_1 _23823_ (.B1(_10210_),
    .Y(_10211_),
    .A1(net6954),
    .A2(_09517_));
 sg13g2_nand3_1 _23824_ (.B(_03796_),
    .C(net6971),
    .A(_03406_),
    .Y(_10212_));
 sg13g2_o21ai_1 _23825_ (.B1(_10212_),
    .Y(_10213_),
    .A1(_03796_),
    .A2(_09387_));
 sg13g2_a21oi_1 _23826_ (.A1(_03796_),
    .A2(net6879),
    .Y(_10214_),
    .B1(_03406_));
 sg13g2_inv_1 _23827_ (.Y(_10215_),
    .A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ));
 sg13g2_a21oi_1 _23828_ (.A1(net6912),
    .A2(_10213_),
    .Y(_10216_),
    .B1(_10214_));
 sg13g2_a221oi_1 _23829_ (.B2(net7296),
    .C1(_10216_),
    .B1(_10211_),
    .A1(net6573),
    .Y(_10217_),
    .A2(_09994_));
 sg13g2_a22oi_1 _23830_ (.Y(_10218_),
    .B1(net6862),
    .B2(_00134_),
    .A2(net6837),
    .A1(_00198_));
 sg13g2_nand2b_1 _23831_ (.Y(_10219_),
    .B(net6709),
    .A_N(_10218_));
 sg13g2_a22oi_1 _23832_ (.Y(_10220_),
    .B1(net6862),
    .B2(_00170_),
    .A2(net6837),
    .A1(_00234_));
 sg13g2_o21ai_1 _23833_ (.B1(_10219_),
    .Y(_10221_),
    .A1(_06865_),
    .A2(_10220_));
 sg13g2_a22oi_1 _23834_ (.Y(_10222_),
    .B1(net6671),
    .B2(_00525_),
    .A2(net6705),
    .A1(_00385_));
 sg13g2_nand2_1 _23835_ (.Y(_10223_),
    .A(net422),
    .B(net6704));
 sg13g2_a21oi_1 _23836_ (.A1(_00420_),
    .A2(net6680),
    .Y(_10224_),
    .B1(net6683));
 sg13g2_a22oi_1 _23837_ (.Y(_10225_),
    .B1(net6691),
    .B2(_00332_),
    .A2(net6696),
    .A1(_00300_));
 sg13g2_a22oi_1 _23838_ (.Y(_10226_),
    .B1(net6676),
    .B2(_00495_),
    .A2(net6780),
    .A1(net371));
 sg13g2_nand3_1 _23839_ (.B(_10225_),
    .C(_10226_),
    .A(_10224_),
    .Y(_10227_));
 sg13g2_a221oi_1 _23840_ (.B2(_00268_),
    .C1(_10227_),
    .B1(net6686),
    .A1(_00370_),
    .Y(_10228_),
    .A2(net6699));
 sg13g2_nand3_1 _23841_ (.B(_10223_),
    .C(_10228_),
    .A(_10222_),
    .Y(_10229_));
 sg13g2_a21o_1 _23842_ (.A2(_10221_),
    .A1(_09539_),
    .B1(_10229_),
    .X(_10230_));
 sg13g2_a21oi_1 _23843_ (.A1(_01663_),
    .A2(net7288),
    .Y(_10231_),
    .B1(_10230_));
 sg13g2_nand3_1 _23844_ (.B(_10217_),
    .C(_10231_),
    .A(net6548),
    .Y(_10232_));
 sg13g2_and3_1 _23845_ (.X(_10233_),
    .A(net6397),
    .B(net7081),
    .C(_10209_));
 sg13g2_and2_1 _23846_ (.A(net7084),
    .B(_10209_),
    .X(_10234_));
 sg13g2_mux4_1 _23847_ (.S0(net7863),
    .A0(_00789_),
    .A1(_00821_),
    .A2(_00853_),
    .A3(_00888_),
    .S1(net7832),
    .X(_10235_));
 sg13g2_a221oi_1 _23848_ (.B2(_00098_),
    .C1(_10233_),
    .B1(_10234_),
    .A1(_10209_),
    .Y(_10236_),
    .A2(_10232_));
 sg13g2_o21ai_1 _23849_ (.B1(_10206_),
    .Y(_10237_),
    .A1(net6392),
    .A2(net5849));
 sg13g2_nand2_1 _23850_ (.Y(_10238_),
    .A(_01585_),
    .B(net6390));
 sg13g2_inv_1 _23851_ (.Y(_10239_),
    .A(_10240_));
 sg13g2_mux4_1 _23852_ (.S0(net7646),
    .A0(net335),
    .A1(net318),
    .A2(net341),
    .A3(net326),
    .S1(net7653),
    .X(_10240_));
 sg13g2_o21ai_1 _23853_ (.B1(_10101_),
    .Y(_10241_),
    .A1(net7662),
    .A2(_10239_));
 sg13g2_nand3b_1 _23854_ (.B(net7008),
    .C(net6970),
    .Y(_10242_),
    .A_N(_03328_));
 sg13g2_o21ai_1 _23855_ (.B1(_10242_),
    .Y(_10243_),
    .A1(net7008),
    .A2(net6905));
 sg13g2_nand2_1 _23856_ (.Y(_10244_),
    .A(net7008),
    .B(net6879));
 sg13g2_a22oi_1 _23857_ (.Y(_10245_),
    .B1(_10244_),
    .B2(_03328_),
    .A2(_10243_),
    .A1(net6911));
 sg13g2_a21oi_1 _23858_ (.A1(net6984),
    .A2(net6575),
    .Y(_10246_),
    .B1(_10245_));
 sg13g2_nor2_1 _23859_ (.A(net6954),
    .B(_09880_),
    .Y(_10247_));
 sg13g2_o21ai_1 _23860_ (.B1(net7294),
    .Y(_10248_),
    .A1(net6964),
    .A2(_09881_));
 sg13g2_o21ai_1 _23861_ (.B1(_10246_),
    .Y(_10249_),
    .A1(_10247_),
    .A2(_10248_));
 sg13g2_nand2_1 _23862_ (.Y(_10250_),
    .A(net7367),
    .B(_10249_));
 sg13g2_a22oi_1 _23863_ (.Y(_10251_),
    .B1(net6704),
    .B2(net421),
    .A2(net6705),
    .A1(_00384_));
 sg13g2_nand2_1 _23864_ (.Y(_10252_),
    .A(_00369_),
    .B(net6700));
 sg13g2_a21oi_1 _23865_ (.A1(_00299_),
    .A2(net6697),
    .Y(_10253_),
    .B1(net6682));
 sg13g2_a22oi_1 _23866_ (.Y(_10254_),
    .B1(net6681),
    .B2(_00419_),
    .A2(net6694),
    .A1(_00331_));
 sg13g2_a22oi_1 _23867_ (.Y(_10255_),
    .B1(net6677),
    .B2(_00494_),
    .A2(net6781),
    .A1(net370));
 sg13g2_nand3_1 _23868_ (.B(_10254_),
    .C(_10255_),
    .A(_10253_),
    .Y(_10256_));
 sg13g2_a221oi_1 _23869_ (.B2(_00524_),
    .C1(_10256_),
    .B1(net6670),
    .A1(_00267_),
    .Y(_10257_),
    .A2(net6687));
 sg13g2_nand3_1 _23870_ (.B(_10252_),
    .C(_10257_),
    .A(_10251_),
    .Y(_10258_));
 sg13g2_a22oi_1 _23871_ (.Y(_10259_),
    .B1(net6868),
    .B2(_00168_),
    .A2(net6833),
    .A1(_00232_));
 sg13g2_a22oi_1 _23872_ (.Y(_10260_),
    .B1(net6868),
    .B2(_00133_),
    .A2(net6833),
    .A1(_00197_));
 sg13g2_nand2b_1 _23873_ (.Y(_10261_),
    .B(net6713),
    .A_N(_10260_));
 sg13g2_o21ai_1 _23874_ (.B1(_10261_),
    .Y(_10262_),
    .A1(_06865_),
    .A2(_10259_));
 sg13g2_a21oi_1 _23875_ (.A1(_09539_),
    .A2(_10262_),
    .Y(_10263_),
    .B1(_10258_));
 sg13g2_nand2_1 _23876_ (.Y(_10264_),
    .A(_01662_),
    .B(net7289));
 sg13g2_nand4_1 _23877_ (.B(_10250_),
    .C(_10263_),
    .A(net6548),
    .Y(_10265_),
    .D(_10264_));
 sg13g2_and2_1 _23878_ (.A(net7081),
    .B(_10241_),
    .X(_10266_));
 sg13g2_and3_1 _23879_ (.X(_10267_),
    .A(_00097_),
    .B(net7084),
    .C(_10241_));
 sg13g2_mux4_1 _23880_ (.S0(net7863),
    .A0(_00923_),
    .A1(_00958_),
    .A2(_00993_),
    .A3(_01029_),
    .S1(net7832),
    .X(_10268_));
 sg13g2_a221oi_1 _23881_ (.B2(net6398),
    .C1(_10267_),
    .B1(_10266_),
    .A1(_10241_),
    .Y(_10269_),
    .A2(_10265_));
 sg13g2_o21ai_1 _23882_ (.B1(_10238_),
    .Y(_10270_),
    .A1(net6390),
    .A2(net5800));
 sg13g2_nand2_1 _23883_ (.Y(_10271_),
    .A(_01584_),
    .B(net6386));
 sg13g2_nor2_1 _23884_ (.A(net6963),
    .B(_09933_),
    .Y(_10272_));
 sg13g2_inv_1 _23885_ (.Y(_10273_),
    .A(_10272_));
 sg13g2_a22oi_1 _23886_ (.Y(_10274_),
    .B1(_09812_),
    .B2(_10272_),
    .A2(_09805_),
    .A1(net6962));
 sg13g2_nand2_1 _23887_ (.Y(_10275_),
    .A(net7293),
    .B(_10274_));
 sg13g2_a22oi_1 _23888_ (.Y(_10276_),
    .B1(net6864),
    .B2(_00132_),
    .A2(net6834),
    .A1(_00196_));
 sg13g2_nand2b_1 _23889_ (.Y(_10277_),
    .B(net6708),
    .A_N(_10276_));
 sg13g2_a22oi_1 _23890_ (.Y(_10278_),
    .B1(net6863),
    .B2(_00167_),
    .A2(net6833),
    .A1(_00231_));
 sg13g2_nand2b_1 _23891_ (.Y(_10279_),
    .B(net7814),
    .A_N(_10268_));
 sg13g2_o21ai_1 _23892_ (.B1(_10277_),
    .Y(_10280_),
    .A1(net6650),
    .A2(_10278_));
 sg13g2_a22oi_1 _23893_ (.Y(_10281_),
    .B1(net6686),
    .B2(_00266_),
    .A2(net6706),
    .A1(_00383_));
 sg13g2_nand2_1 _23894_ (.Y(_10282_),
    .A(net420),
    .B(net6704));
 sg13g2_a21oi_1 _23895_ (.A1(_00298_),
    .A2(net6697),
    .Y(_10283_),
    .B1(net6682));
 sg13g2_a22oi_1 _23896_ (.Y(_10284_),
    .B1(net6681),
    .B2(_00418_),
    .A2(net6694),
    .A1(_00330_));
 sg13g2_a22oi_1 _23897_ (.Y(_10285_),
    .B1(net6677),
    .B2(_00493_),
    .A2(net6781),
    .A1(net369));
 sg13g2_nand3_1 _23898_ (.B(_10284_),
    .C(_10285_),
    .A(_10283_),
    .Y(_10286_));
 sg13g2_o21ai_1 _23899_ (.B1(_10279_),
    .Y(_10287_),
    .A1(net7814),
    .A2(_10235_));
 sg13g2_a221oi_1 _23900_ (.B2(_00523_),
    .C1(_10286_),
    .B1(net6672),
    .A1(_00368_),
    .Y(_10288_),
    .A2(net6699));
 sg13g2_nand3_1 _23901_ (.B(_10282_),
    .C(_10288_),
    .A(_10281_),
    .Y(_10289_));
 sg13g2_a21oi_1 _23902_ (.A1(net6797),
    .A2(_10280_),
    .Y(_10290_),
    .B1(_10289_));
 sg13g2_nor2_1 _23903_ (.A(_03785_),
    .B(net6906),
    .Y(_10291_));
 sg13g2_nor3_1 _23904_ (.A(_03257_),
    .B(_03784_),
    .C(_09389_),
    .Y(_10292_));
 sg13g2_o21ai_1 _23905_ (.B1(net6908),
    .Y(_10293_),
    .A1(_10291_),
    .A2(_10292_));
 sg13g2_o21ai_1 _23906_ (.B1(_03257_),
    .Y(_10294_),
    .A1(_03784_),
    .A2(_09393_));
 sg13g2_a22oi_1 _23907_ (.Y(_10295_),
    .B1(_10293_),
    .B2(_10294_),
    .A2(net7288),
    .A1(_01661_));
 sg13g2_a21oi_1 _23908_ (.A1(net6576),
    .A2(net6902),
    .Y(_10296_),
    .B1(net6547));
 sg13g2_nand4_1 _23909_ (.B(_10290_),
    .C(_10295_),
    .A(_10275_),
    .Y(_10297_),
    .D(_10296_));
 sg13g2_a21o_1 _23910_ (.A2(_08742_),
    .A1(net6399),
    .B1(_10297_),
    .X(_10298_));
 sg13g2_mux2_1 _23911_ (.A0(_00661_),
    .A1(_00693_),
    .S(net7860),
    .X(_10299_));
 sg13g2_nor2_1 _23912_ (.A(net7510),
    .B(_10299_),
    .Y(_10300_));
 sg13g2_a21oi_1 _23913_ (.A1(net5924),
    .A2(net7087),
    .Y(_10301_),
    .B1(_10298_));
 sg13g2_nor2b_1 _23914_ (.A(net7651),
    .B_N(net317),
    .Y(_10302_));
 sg13g2_a21oi_1 _23915_ (.A1(net325),
    .A2(net7651),
    .Y(_10303_),
    .B1(_10302_));
 sg13g2_nand2_1 _23916_ (.Y(_10304_),
    .A(net7644),
    .B(_10303_));
 sg13g2_mux2_1 _23917_ (.A0(net334),
    .A1(net338),
    .S(net7655),
    .X(_10305_));
 sg13g2_o21ai_1 _23918_ (.B1(_10304_),
    .Y(_10306_),
    .A1(net7644),
    .A2(_10305_));
 sg13g2_o21ai_1 _23919_ (.B1(net6464),
    .Y(_10307_),
    .A1(net7663),
    .A2(_10306_));
 sg13g2_nand2b_1 _23920_ (.Y(_10308_),
    .B(_10307_),
    .A_N(net5846));
 sg13g2_o21ai_1 _23921_ (.B1(_10271_),
    .Y(_10309_),
    .A1(net6018),
    .A2(net5797));
 sg13g2_nand2_1 _23922_ (.Y(_10310_),
    .A(_01583_),
    .B(net6393));
 sg13g2_a22oi_1 _23923_ (.Y(_10311_),
    .B1(_10272_),
    .B2(_09706_),
    .A2(_09750_),
    .A1(net6962));
 sg13g2_nand2_1 _23924_ (.Y(_10312_),
    .A(net7293),
    .B(_10311_));
 sg13g2_a22oi_1 _23925_ (.Y(_10313_),
    .B1(net6864),
    .B2(_00131_),
    .A2(net6835),
    .A1(_00195_));
 sg13g2_nand2b_1 _23926_ (.Y(_10314_),
    .B(net6708),
    .A_N(_10313_));
 sg13g2_a22oi_1 _23927_ (.Y(_10315_),
    .B1(net6863),
    .B2(_00166_),
    .A2(net6833),
    .A1(_00230_));
 sg13g2_o21ai_1 _23928_ (.B1(_10314_),
    .Y(_10316_),
    .A1(net6650),
    .A2(_10315_));
 sg13g2_a22oi_1 _23929_ (.Y(_10317_),
    .B1(net6686),
    .B2(_00265_),
    .A2(net6706),
    .A1(_00399_));
 sg13g2_nand2_1 _23930_ (.Y(_10318_),
    .A(net433),
    .B(net6703));
 sg13g2_a21oi_1 _23931_ (.A1(_00297_),
    .A2(net6697),
    .Y(_10319_),
    .B1(net6682));
 sg13g2_mux2_1 _23932_ (.A0(_00725_),
    .A1(_00757_),
    .S(net7860),
    .X(_10320_));
 sg13g2_a22oi_1 _23933_ (.Y(_10321_),
    .B1(net6680),
    .B2(_00417_),
    .A2(net6694),
    .A1(_00329_));
 sg13g2_a22oi_1 _23934_ (.Y(_10322_),
    .B1(net6677),
    .B2(_00492_),
    .A2(net6781),
    .A1(net368));
 sg13g2_nand3_1 _23935_ (.B(_10321_),
    .C(_10322_),
    .A(_10319_),
    .Y(_10323_));
 sg13g2_nor2_1 _23936_ (.A(_09004_),
    .B(_10320_),
    .Y(_10324_));
 sg13g2_a221oi_1 _23937_ (.B2(_00522_),
    .C1(_10323_),
    .B1(net6672),
    .A1(_00367_),
    .Y(_10325_),
    .A2(net6699));
 sg13g2_nand3_1 _23938_ (.B(_10318_),
    .C(_10325_),
    .A(_10317_),
    .Y(_10326_));
 sg13g2_a21oi_1 _23939_ (.A1(net6797),
    .A2(_10316_),
    .Y(_10327_),
    .B1(_10326_));
 sg13g2_nor2_1 _23940_ (.A(_03780_),
    .B(net6906),
    .Y(_10328_));
 sg13g2_nor3_1 _23941_ (.A(_03193_),
    .B(net7009),
    .C(_09389_),
    .Y(_10329_));
 sg13g2_o21ai_1 _23942_ (.B1(net6910),
    .Y(_10330_),
    .A1(_10328_),
    .A2(_10329_));
 sg13g2_o21ai_1 _23943_ (.B1(_03193_),
    .Y(_10331_),
    .A1(net7009),
    .A2(_09393_));
 sg13g2_a22oi_1 _23944_ (.Y(_10332_),
    .B1(_10330_),
    .B2(_10331_),
    .A2(net7288),
    .A1(_01659_));
 sg13g2_a21oi_1 _23945_ (.A1(net6579),
    .A2(net6902),
    .Y(_10333_),
    .B1(net6547));
 sg13g2_nand4_1 _23946_ (.B(_10327_),
    .C(_10332_),
    .A(_10312_),
    .Y(_10334_),
    .D(_10333_));
 sg13g2_a21o_1 _23947_ (.A2(_08742_),
    .A1(net6400),
    .B1(_10334_),
    .X(_10335_));
 sg13g2_mux2_1 _23948_ (.A0(_01225_),
    .A1(_01577_),
    .S(net7860),
    .X(_10336_));
 sg13g2_a21oi_1 _23949_ (.A1(_00095_),
    .A2(net7084),
    .Y(_10337_),
    .B1(_10335_));
 sg13g2_a221oi_1 _23950_ (.B2(net7834),
    .C1(_01894_),
    .B1(_10336_),
    .A1(_00873_),
    .Y(_10338_),
    .A2(_08988_));
 sg13g2_inv_1 _23951_ (.Y(_10339_),
    .A(_10340_));
 sg13g2_mux4_1 _23952_ (.S0(net7645),
    .A0(net333),
    .A1(net347),
    .A2(net327),
    .A3(net324),
    .S1(net7652),
    .X(_10340_));
 sg13g2_o21ai_1 _23953_ (.B1(net6463),
    .Y(_10341_),
    .A1(net7662),
    .A2(_10339_));
 sg13g2_nand2b_1 _23954_ (.Y(_10342_),
    .B(net6379),
    .A_N(net6393));
 sg13g2_o21ai_1 _23955_ (.B1(_10310_),
    .Y(_10343_),
    .A1(net5919),
    .A2(_10342_));
 sg13g2_or3_1 _23956_ (.A(_10300_),
    .B(_10324_),
    .C(_10338_),
    .X(_10344_));
 sg13g2_nand2_1 _23957_ (.Y(_10345_),
    .A(_01582_),
    .B(net6386));
 sg13g2_a21oi_1 _23958_ (.A1(_09650_),
    .A2(_10272_),
    .Y(_10346_),
    .B1(_08205_));
 sg13g2_o21ai_1 _23959_ (.B1(_10346_),
    .Y(_10347_),
    .A1(net6955),
    .A2(_09641_));
 sg13g2_a22oi_1 _23960_ (.Y(_10348_),
    .B1(net6703),
    .B2(net432),
    .A2(net6706),
    .A1(_00398_));
 sg13g2_nand2_1 _23961_ (.Y(_10349_),
    .A(_00366_),
    .B(net6700));
 sg13g2_a21oi_1 _23962_ (.A1(_00296_),
    .A2(net6695),
    .Y(_10350_),
    .B1(net6684));
 sg13g2_a22oi_1 _23963_ (.Y(_10351_),
    .B1(_10344_),
    .B2(net7530),
    .A2(_10287_),
    .A1(net7546));
 sg13g2_a22oi_1 _23964_ (.Y(_10352_),
    .B1(net6681),
    .B2(_00416_),
    .A2(net6693),
    .A1(_00328_));
 sg13g2_a22oi_1 _23965_ (.Y(_10353_),
    .B1(net6677),
    .B2(_00491_),
    .A2(net6781),
    .A1(net367));
 sg13g2_nand3_1 _23966_ (.B(_10352_),
    .C(_10353_),
    .A(_10350_),
    .Y(_10354_));
 sg13g2_a221oi_1 _23967_ (.B2(_00521_),
    .C1(_10354_),
    .B1(net6670),
    .A1(_00264_),
    .Y(_10355_),
    .A2(net6686));
 sg13g2_nand3_1 _23968_ (.B(_10349_),
    .C(_10355_),
    .A(_10348_),
    .Y(_10356_));
 sg13g2_a22oi_1 _23969_ (.Y(_10357_),
    .B1(net6863),
    .B2(_00165_),
    .A2(net6833),
    .A1(_00229_));
 sg13g2_a22oi_1 _23970_ (.Y(_10358_),
    .B1(net6864),
    .B2(_00130_),
    .A2(net6835),
    .A1(_00194_));
 sg13g2_nand2b_1 _23971_ (.Y(_10359_),
    .B(net6713),
    .A_N(_10358_));
 sg13g2_o21ai_1 _23972_ (.B1(_10359_),
    .Y(_10360_),
    .A1(net6650),
    .A2(_10357_));
 sg13g2_a21oi_1 _23973_ (.A1(net6797),
    .A2(_10360_),
    .Y(_10361_),
    .B1(_10356_));
 sg13g2_nand3b_1 _23974_ (.B(net7010),
    .C(net6970),
    .Y(_10362_),
    .A_N(net7030));
 sg13g2_o21ai_1 _23975_ (.B1(_10362_),
    .Y(_10363_),
    .A1(net7010),
    .A2(net6904));
 sg13g2_nand2_1 _23976_ (.Y(_10364_),
    .A(net7010),
    .B(net6878));
 sg13g2_a22oi_1 _23977_ (.Y(_10365_),
    .B1(_10364_),
    .B2(net7030),
    .A2(_10363_),
    .A1(net6910));
 sg13g2_a21oi_1 _23978_ (.A1(_01658_),
    .A2(net7288),
    .Y(_10366_),
    .B1(_10365_));
 sg13g2_a221oi_1 _23979_ (.B2(net6582),
    .C1(net6547),
    .B1(net6902),
    .A1(net6478),
    .Y(_10367_),
    .A2(net7082));
 sg13g2_nand4_1 _23980_ (.B(_10361_),
    .C(_10366_),
    .A(_10347_),
    .Y(_10368_),
    .D(_10367_));
 sg13g2_a21oi_1 _23981_ (.A1(_00094_),
    .A2(net7088),
    .Y(_10369_),
    .B1(_10368_));
 sg13g2_nand2_1 _23982_ (.Y(_10370_),
    .A(_10200_),
    .B(_10351_));
 sg13g2_mux4_1 _23983_ (.S0(net7642),
    .A0(net332),
    .A1(net346),
    .A2(net316),
    .A3(net323),
    .S1(net7649),
    .X(_10371_));
 sg13g2_nand2_1 _23984_ (.Y(_10372_),
    .A(net7628),
    .B(_10371_));
 sg13g2_a21o_1 _23985_ (.A2(_10372_),
    .A1(net6465),
    .B1(net5845),
    .X(_10373_));
 sg13g2_o21ai_1 _23986_ (.B1(_10345_),
    .Y(_10374_),
    .A1(net6018),
    .A2(net5789));
 sg13g2_nand2_1 _23987_ (.Y(_10375_),
    .A(_01581_),
    .B(net6387));
 sg13g2_a221oi_1 _23988_ (.B2(net8007),
    .C1(_09978_),
    .B1(_10370_),
    .A1(net7354),
    .Y(_10376_),
    .A2(net7077));
 sg13g2_nand3b_1 _23989_ (.B(_03769_),
    .C(net6970),
    .Y(_10377_),
    .A_N(_03054_));
 sg13g2_o21ai_1 _23990_ (.B1(_10377_),
    .Y(_10378_),
    .A1(_03769_),
    .A2(net6904));
 sg13g2_nand2_1 _23991_ (.Y(_10379_),
    .A(_03769_),
    .B(net6878));
 sg13g2_a22oi_1 _23992_ (.Y(_10380_),
    .B1(_10379_),
    .B2(_03054_),
    .A2(_10378_),
    .A1(net6910));
 sg13g2_nor2_1 _23993_ (.A(net6754),
    .B(_10029_),
    .Y(_10381_));
 sg13g2_nor2_1 _23994_ (.A(_09933_),
    .B(_10381_),
    .Y(_10382_));
 sg13g2_nor2_1 _23995_ (.A(net6756),
    .B(_09649_),
    .Y(_10383_));
 sg13g2_a21oi_1 _23996_ (.A1(_09405_),
    .A2(_10042_),
    .Y(_10384_),
    .B1(_10383_));
 sg13g2_nor2_1 _23997_ (.A(net6799),
    .B(_10382_),
    .Y(_10385_));
 sg13g2_a21oi_1 _23998_ (.A1(net6799),
    .A2(_10384_),
    .Y(_10386_),
    .B1(_10385_));
 sg13g2_nor2_1 _23999_ (.A(_09402_),
    .B(_09631_),
    .Y(_10387_));
 sg13g2_a21oi_1 _24000_ (.A1(_09402_),
    .A2(_09635_),
    .Y(_10388_),
    .B1(_10387_));
 sg13g2_nor2_1 _24001_ (.A(_09406_),
    .B(_10388_),
    .Y(_10389_));
 sg13g2_inv_1 _24002_ (.Y(_10390_),
    .A(_10389_));
 sg13g2_a22oi_1 _24003_ (.Y(_10391_),
    .B1(_10390_),
    .B2(_10272_),
    .A2(_10386_),
    .A1(net6964));
 sg13g2_a221oi_1 _24004_ (.B2(net7295),
    .C1(_10380_),
    .B1(_10391_),
    .A1(net6983),
    .Y(_10392_),
    .A2(net6603));
 sg13g2_a22oi_1 _24005_ (.Y(_10393_),
    .B1(net6687),
    .B2(_00263_),
    .A2(_09558_),
    .A1(_00397_));
 sg13g2_nand2_1 _24006_ (.Y(_10394_),
    .A(_00365_),
    .B(net6700));
 sg13g2_a21oi_1 _24007_ (.A1(_00295_),
    .A2(net6695),
    .Y(_10395_),
    .B1(net6684));
 sg13g2_a22oi_1 _24008_ (.Y(_10396_),
    .B1(net6681),
    .B2(_00415_),
    .A2(net6693),
    .A1(_00327_));
 sg13g2_a22oi_1 _24009_ (.Y(_10397_),
    .B1(net6677),
    .B2(_00490_),
    .A2(net6781),
    .A1(net366));
 sg13g2_nand3_1 _24010_ (.B(_10396_),
    .C(_10397_),
    .A(_10395_),
    .Y(_10398_));
 sg13g2_a221oi_1 _24011_ (.B2(_00520_),
    .C1(_10398_),
    .B1(net6670),
    .A1(net431),
    .Y(_10399_),
    .A2(net6703));
 sg13g2_nand3_1 _24012_ (.B(_10394_),
    .C(_10399_),
    .A(_10393_),
    .Y(_10400_));
 sg13g2_a22oi_1 _24013_ (.Y(_10401_),
    .B1(net6863),
    .B2(_00164_),
    .A2(net6833),
    .A1(_00228_));
 sg13g2_a22oi_1 _24014_ (.Y(_10402_),
    .B1(net6864),
    .B2(_00129_),
    .A2(net6835),
    .A1(_00193_));
 sg13g2_nand2b_1 _24015_ (.Y(_10403_),
    .B(net6713),
    .A_N(_10402_));
 sg13g2_o21ai_1 _24016_ (.B1(_10403_),
    .Y(_10404_),
    .A1(net6650),
    .A2(_10401_));
 sg13g2_mux2_1 _24017_ (.A0(_08254_),
    .A1(net6981),
    .S(_09945_),
    .X(_10405_));
 sg13g2_a21oi_1 _24018_ (.A1(net6797),
    .A2(_10404_),
    .Y(_10406_),
    .B1(_10400_));
 sg13g2_nand2_1 _24019_ (.Y(_10407_),
    .A(net7978),
    .B(net7289));
 sg13g2_nand3_1 _24020_ (.B(_10406_),
    .C(_10407_),
    .A(net6548),
    .Y(_10408_));
 sg13g2_a21oi_1 _24021_ (.A1(net6557),
    .A2(_08742_),
    .Y(_10409_),
    .B1(_10408_));
 sg13g2_o21ai_1 _24022_ (.B1(_10409_),
    .Y(_10410_),
    .A1(net7382),
    .A2(_10392_));
 sg13g2_a21oi_1 _24023_ (.A1(_00093_),
    .A2(net7084),
    .Y(_10411_),
    .B1(_10410_));
 sg13g2_inv_1 _24024_ (.Y(_10412_),
    .A(_10413_));
 sg13g2_mux4_1 _24025_ (.S0(net7656),
    .A0(net331),
    .A1(_02009_),
    .A2(net345),
    .A3(net322),
    .S1(net7648),
    .X(_10413_));
 sg13g2_o21ai_1 _24026_ (.B1(_10405_),
    .Y(_10414_),
    .A1(net7364),
    .A2(_10376_));
 sg13g2_o21ai_1 _24027_ (.B1(net6464),
    .Y(_10415_),
    .A1(net7663),
    .A2(_10412_));
 sg13g2_nand2b_1 _24028_ (.Y(_10416_),
    .B(net6373),
    .A_N(net6387));
 sg13g2_inv_1 _24029_ (.Y(_10417_),
    .A(_01862_));
 sg13g2_o21ai_1 _24030_ (.B1(_10375_),
    .Y(_10418_),
    .A1(net5914),
    .A2(_10416_));
 sg13g2_nand2_1 _24031_ (.Y(_10419_),
    .A(_01580_),
    .B(net6386));
 sg13g2_nor2_1 _24032_ (.A(net6753),
    .B(_09976_),
    .Y(_10420_));
 sg13g2_or3_1 _24033_ (.A(net6800),
    .B(_09933_),
    .C(_10420_),
    .X(_10421_));
 sg13g2_mux2_1 _24034_ (.A0(_09705_),
    .A1(_09964_),
    .S(net6757),
    .X(_10422_));
 sg13g2_o21ai_1 _24035_ (.B1(_10421_),
    .Y(_10423_),
    .A1(net6798),
    .A2(_10422_));
 sg13g2_a21oi_1 _24036_ (.A1(net6756),
    .A2(_09719_),
    .Y(_10424_),
    .B1(_10048_));
 sg13g2_nand2_1 _24037_ (.Y(_10425_),
    .A(net6957),
    .B(_10424_));
 sg13g2_o21ai_1 _24038_ (.B1(_10425_),
    .Y(_10426_),
    .A1(net6957),
    .A2(_10423_));
 sg13g2_a22oi_1 _24039_ (.Y(_10427_),
    .B1(net6864),
    .B2(_00128_),
    .A2(net6835),
    .A1(_00192_));
 sg13g2_nand2b_1 _24040_ (.Y(_10428_),
    .B(net6708),
    .A_N(_10427_));
 sg13g2_a22oi_1 _24041_ (.Y(_10429_),
    .B1(net6863),
    .B2(_00163_),
    .A2(net6833),
    .A1(_00227_));
 sg13g2_o21ai_1 _24042_ (.B1(_10428_),
    .Y(_10430_),
    .A1(net6650),
    .A2(_10429_));
 sg13g2_a22oi_1 _24043_ (.Y(_10431_),
    .B1(net6703),
    .B2(net430),
    .A2(_09558_),
    .A1(_00396_));
 sg13g2_nand2_1 _24044_ (.Y(_10432_),
    .A(_00364_),
    .B(net6700));
 sg13g2_a21oi_1 _24045_ (.A1(_00294_),
    .A2(net6695),
    .Y(_10433_),
    .B1(net6684));
 sg13g2_mux4_1 _24046_ (.S0(net7777),
    .A0(_00790_),
    .A1(_00822_),
    .A2(_00854_),
    .A3(_00889_),
    .S1(net7726),
    .X(_10434_));
 sg13g2_a22oi_1 _24047_ (.Y(_10435_),
    .B1(net6681),
    .B2(_00414_),
    .A2(net6694),
    .A1(_00326_));
 sg13g2_a22oi_1 _24048_ (.Y(_10436_),
    .B1(net6677),
    .B2(_00489_),
    .A2(net6781),
    .A1(net365));
 sg13g2_nand3_1 _24049_ (.B(_10435_),
    .C(_10436_),
    .A(_10433_),
    .Y(_10437_));
 sg13g2_nand2_1 _24050_ (.Y(_10438_),
    .A(_08255_),
    .B(_10434_));
 sg13g2_a221oi_1 _24051_ (.B2(_00519_),
    .C1(_10437_),
    .B1(net6670),
    .A1(_00262_),
    .Y(_10439_),
    .A2(net6688));
 sg13g2_nand3_1 _24052_ (.B(_10432_),
    .C(_10439_),
    .A(_10431_),
    .Y(_10440_));
 sg13g2_a21oi_1 _24053_ (.A1(net6797),
    .A2(_10430_),
    .Y(_10441_),
    .B1(_10440_));
 sg13g2_nand2_1 _24054_ (.Y(_10442_),
    .A(_02987_),
    .B(_03764_));
 sg13g2_nor2_1 _24055_ (.A(_02987_),
    .B(_03764_),
    .Y(_10443_));
 sg13g2_o21ai_1 _24056_ (.B1(net6910),
    .Y(_10444_),
    .A1(_09388_),
    .A2(_10443_));
 sg13g2_nor3_1 _24057_ (.A(_02987_),
    .B(_03764_),
    .C(net6970),
    .Y(_10445_));
 sg13g2_a221oi_1 _24058_ (.B2(_10444_),
    .C1(_10445_),
    .B1(_10442_),
    .A1(_01656_),
    .Y(_10446_),
    .A2(net7288));
 sg13g2_nand3_1 _24059_ (.B(_10441_),
    .C(_10446_),
    .A(net6550),
    .Y(_10447_));
 sg13g2_a221oi_1 _24060_ (.B2(net7293),
    .C1(_10447_),
    .B1(_10426_),
    .A1(net6605),
    .Y(_10448_),
    .A2(net6902));
 sg13g2_and2_1 _24061_ (.A(_08305_),
    .B(_08313_),
    .X(_10449_));
 sg13g2_nand3_1 _24062_ (.B(_08871_),
    .C(_10448_),
    .A(_08863_),
    .Y(_10450_));
 sg13g2_nand2_1 _24063_ (.Y(_10451_),
    .A(net7643),
    .B(_09690_));
 sg13g2_mux2_1 _24064_ (.A0(net330),
    .A1(_02008_),
    .S(net7652),
    .X(_10452_));
 sg13g2_o21ai_1 _24065_ (.B1(_10451_),
    .Y(_10453_),
    .A1(net7643),
    .A2(_10452_));
 sg13g2_mux2_1 _24066_ (.A0(_01588_),
    .A1(_00758_),
    .S(net7715),
    .X(_10454_));
 sg13g2_o21ai_1 _24067_ (.B1(net6464),
    .Y(_10455_),
    .A1(net7663),
    .A2(_10453_));
 sg13g2_nand2_1 _24068_ (.Y(_10456_),
    .A(net5844),
    .B(_10455_));
 sg13g2_o21ai_1 _24069_ (.B1(_10419_),
    .Y(_10457_),
    .A1(net6018),
    .A2(net5778));
 sg13g2_nand2_1 _24070_ (.Y(_10458_),
    .A(_01579_),
    .B(net6387));
 sg13g2_a21oi_1 _24071_ (.A1(net6756),
    .A2(_09789_),
    .Y(_10459_),
    .B1(_10048_));
 sg13g2_mux4_1 _24072_ (.S0(net6802),
    .A0(_09519_),
    .A1(_09810_),
    .A2(_09918_),
    .A3(_09923_),
    .S1(net6758),
    .X(_10460_));
 sg13g2_nand2_1 _24073_ (.Y(_10461_),
    .A(net6956),
    .B(_10459_));
 sg13g2_o21ai_1 _24074_ (.B1(_10461_),
    .Y(_10462_),
    .A1(net6956),
    .A2(_10460_));
 sg13g2_and2_1 _24075_ (.A(_08305_),
    .B(_08307_),
    .X(_10463_));
 sg13g2_nor3_1 _24076_ (.A(_02920_),
    .B(_03759_),
    .C(_09389_),
    .Y(_10464_));
 sg13g2_inv_1 _24077_ (.Y(_10465_),
    .A(_10463_));
 sg13g2_a21o_1 _24078_ (.A2(_09388_),
    .A1(_03759_),
    .B1(_10464_),
    .X(_10466_));
 sg13g2_nand2_1 _24079_ (.Y(_10467_),
    .A(_03760_),
    .B(net6879));
 sg13g2_a22oi_1 _24080_ (.Y(_10468_),
    .B1(_10467_),
    .B2(_02920_),
    .A2(_10466_),
    .A1(net6911));
 sg13g2_a221oi_1 _24081_ (.B2(net7295),
    .C1(_10468_),
    .B1(_10462_),
    .A1(net6983),
    .Y(_10469_),
    .A2(net6584));
 sg13g2_a21oi_1 _24082_ (.A1(net7923),
    .A2(net7979),
    .Y(_10470_),
    .B1(net7367));
 sg13g2_a21o_1 _24083_ (.A2(_10469_),
    .A1(net7367),
    .B1(_10470_),
    .X(_10471_));
 sg13g2_a22oi_1 _24084_ (.Y(_10472_),
    .B1(_09547_),
    .B2(\cs_registers_i.csr_mstatus_tw_o ),
    .A2(net6779),
    .A1(net364));
 sg13g2_a21oi_1 _24085_ (.A1(_00293_),
    .A2(net6695),
    .Y(_10473_),
    .B1(net6684));
 sg13g2_a22oi_1 _24086_ (.Y(_10474_),
    .B1(net6681),
    .B2(_00413_),
    .A2(net6693),
    .A1(_00325_));
 sg13g2_nand3_1 _24087_ (.B(_10473_),
    .C(_10474_),
    .A(_10472_),
    .Y(_10475_));
 sg13g2_a221oi_1 _24088_ (.B2(_00488_),
    .C1(_10475_),
    .B1(net6674),
    .A1(_00395_),
    .Y(_10476_),
    .A2(_09558_));
 sg13g2_a21oi_1 _24089_ (.A1(_08288_),
    .A2(_10454_),
    .Y(_10477_),
    .B1(net7691));
 sg13g2_a22oi_1 _24090_ (.Y(_10478_),
    .B1(net6670),
    .B2(_00518_),
    .A2(net6689),
    .A1(_00261_));
 sg13g2_a22oi_1 _24091_ (.Y(_10479_),
    .B1(net6700),
    .B2(_00363_),
    .A2(net6703),
    .A1(net429));
 sg13g2_nand3_1 _24092_ (.B(_10478_),
    .C(_10479_),
    .A(_10476_),
    .Y(_10480_));
 sg13g2_a22oi_1 _24093_ (.Y(_10481_),
    .B1(net6863),
    .B2(_00162_),
    .A2(net6835),
    .A1(_00226_));
 sg13g2_a22oi_1 _24094_ (.Y(_10482_),
    .B1(net6864),
    .B2(_00127_),
    .A2(net6834),
    .A1(_00191_));
 sg13g2_nand2b_1 _24095_ (.Y(_10483_),
    .B(net6713),
    .A_N(_10482_));
 sg13g2_o21ai_1 _24096_ (.B1(_10483_),
    .Y(_10484_),
    .A1(net6649),
    .A2(_10481_));
 sg13g2_a21oi_1 _24097_ (.A1(net6797),
    .A2(_10484_),
    .Y(_10485_),
    .B1(_10480_));
 sg13g2_a21oi_1 _24098_ (.A1(_00107_),
    .A2(net7082),
    .Y(_10486_),
    .B1(net6547));
 sg13g2_nand3_1 _24099_ (.B(_10485_),
    .C(_10486_),
    .A(_10471_),
    .Y(_10487_));
 sg13g2_a21oi_1 _24100_ (.A1(_00091_),
    .A2(net7087),
    .Y(_10488_),
    .B1(_10487_));
 sg13g2_nand2_1 _24101_ (.Y(_10489_),
    .A(net7641),
    .B(_09836_));
 sg13g2_mux2_1 _24102_ (.A0(net329),
    .A1(_02007_),
    .S(_01986_),
    .X(_10490_));
 sg13g2_o21ai_1 _24103_ (.B1(_10489_),
    .Y(_10491_),
    .A1(net7641),
    .A2(_10490_));
 sg13g2_a22oi_1 _24104_ (.Y(_10492_),
    .B1(_10463_),
    .B2(_00884_),
    .A2(_10449_),
    .A1(_01236_));
 sg13g2_o21ai_1 _24105_ (.B1(net6465),
    .Y(_10493_),
    .A1(_00007_),
    .A2(_10491_));
 sg13g2_nand2b_1 _24106_ (.Y(_10494_),
    .B(net6366),
    .A_N(net6387));
 sg13g2_o21ai_1 _24107_ (.B1(_10458_),
    .Y(_10495_),
    .A1(net5910),
    .A2(_10494_));
 sg13g2_a21oi_1 _24108_ (.A1(net6756),
    .A2(_09488_),
    .Y(_10496_),
    .B1(_10048_));
 sg13g2_nand2_1 _24109_ (.Y(_10497_),
    .A(net6799),
    .B(_09456_));
 sg13g2_o21ai_1 _24110_ (.B1(_10497_),
    .Y(_10498_),
    .A1(net6799),
    .A2(_10496_));
 sg13g2_nor2_1 _24111_ (.A(net6800),
    .B(_09530_),
    .Y(_10499_));
 sg13g2_a21oi_1 _24112_ (.A1(net6800),
    .A2(_09864_),
    .Y(_10500_),
    .B1(_10499_));
 sg13g2_nor2_1 _24113_ (.A(_09406_),
    .B(_10500_),
    .Y(_10501_));
 sg13g2_inv_1 _24114_ (.Y(_10502_),
    .A(_10501_));
 sg13g2_a22oi_1 _24115_ (.Y(_10503_),
    .B1(_10502_),
    .B2(_10272_),
    .A2(_10498_),
    .A1(net6962));
 sg13g2_nand2_1 _24116_ (.Y(_10504_),
    .A(net7293),
    .B(_10503_));
 sg13g2_a22oi_1 _24117_ (.Y(_10505_),
    .B1(net6865),
    .B2(_00126_),
    .A2(net6835),
    .A1(_00190_));
 sg13g2_nand2b_1 _24118_ (.Y(_10506_),
    .B(net6709),
    .A_N(_10505_));
 sg13g2_a22oi_1 _24119_ (.Y(_10507_),
    .B1(net6865),
    .B2(_00161_),
    .A2(net6835),
    .A1(_00225_));
 sg13g2_o21ai_1 _24120_ (.B1(_10506_),
    .Y(_10508_),
    .A1(net6649),
    .A2(_10507_));
 sg13g2_a22oi_1 _24121_ (.Y(_10509_),
    .B1(_09567_),
    .B2(_00324_),
    .A2(_09566_),
    .A1(_00292_));
 sg13g2_nand2_1 _24122_ (.Y(_10510_),
    .A(_00412_),
    .B(_09570_));
 sg13g2_a22oi_1 _24123_ (.Y(_10511_),
    .B1(net6677),
    .B2(_00487_),
    .A2(_06886_),
    .A1(net363));
 sg13g2_nand3_1 _24124_ (.B(_10510_),
    .C(_10511_),
    .A(_10509_),
    .Y(_10512_));
 sg13g2_a221oi_1 _24125_ (.B2(_00517_),
    .C1(_10512_),
    .B1(net6672),
    .A1(_00394_),
    .Y(_10513_),
    .A2(net6706));
 sg13g2_a21oi_1 _24126_ (.A1(net428),
    .A2(net6704),
    .Y(_10514_),
    .B1(_10147_));
 sg13g2_a22oi_1 _24127_ (.Y(_10515_),
    .B1(net6689),
    .B2(_00260_),
    .A2(net6702),
    .A1(_00362_));
 sg13g2_nand3_1 _24128_ (.B(_10514_),
    .C(_10515_),
    .A(_10513_),
    .Y(_10516_));
 sg13g2_a21oi_1 _24129_ (.A1(net6797),
    .A2(_10508_),
    .Y(_10517_),
    .B1(_10516_));
 sg13g2_nor2_1 _24130_ (.A(_03755_),
    .B(net6906),
    .Y(_10518_));
 sg13g2_nor3_1 _24131_ (.A(_02853_),
    .B(_03754_),
    .C(_09389_),
    .Y(_10519_));
 sg13g2_o21ai_1 _24132_ (.B1(net6910),
    .Y(_10520_),
    .A1(_10518_),
    .A2(_10519_));
 sg13g2_o21ai_1 _24133_ (.B1(_02853_),
    .Y(_10521_),
    .A1(_03754_),
    .A2(_09393_));
 sg13g2_a22oi_1 _24134_ (.Y(_10522_),
    .B1(_10520_),
    .B2(_10521_),
    .A2(net7288),
    .A1(net7980));
 sg13g2_mux4_1 _24135_ (.S0(net7778),
    .A0(_00924_),
    .A1(_00959_),
    .A2(_00995_),
    .A3(_01030_),
    .S1(net7728),
    .X(_10523_));
 sg13g2_a221oi_1 _24136_ (.B2(net6586),
    .C1(net6547),
    .B1(net6902),
    .A1(net6620),
    .Y(_10524_),
    .A2(net7082));
 sg13g2_nand4_1 _24137_ (.B(_10517_),
    .C(_10522_),
    .A(_10504_),
    .Y(_10525_),
    .D(_10524_));
 sg13g2_mux2_1 _24138_ (.A0(_00662_),
    .A1(_00694_),
    .S(net7776),
    .X(_10526_));
 sg13g2_a21oi_1 _24139_ (.A1(net5954),
    .A2(net7088),
    .Y(_10527_),
    .B1(_10525_));
 sg13g2_nand2_1 _24140_ (.Y(_10528_),
    .A(net7643),
    .B(_09849_));
 sg13g2_mux2_1 _24141_ (.A0(net328),
    .A1(_02006_),
    .S(net7652),
    .X(_10529_));
 sg13g2_o21ai_1 _24142_ (.B1(_10528_),
    .Y(_10530_),
    .A1(net7643),
    .A2(_10529_));
 sg13g2_o21ai_1 _24143_ (.B1(net6463),
    .Y(_10531_),
    .A1(net7663),
    .A2(_10530_));
 sg13g2_nor2b_1 _24144_ (.A(net5906),
    .B_N(_10531_),
    .Y(_10532_));
 sg13g2_mux2_1 _24145_ (.A0(net5839),
    .A1(_01578_),
    .S(_10095_),
    .X(_10533_));
 sg13g2_nand2_1 _24146_ (.Y(_10534_),
    .A(_01577_),
    .B(net6050));
 sg13g2_o21ai_1 _24147_ (.B1(_10534_),
    .Y(_10535_),
    .A1(net6050),
    .A2(net6108));
 sg13g2_nand2_1 _24148_ (.Y(_10536_),
    .A(_01576_),
    .B(_10093_));
 sg13g2_nand3_1 _24149_ (.B(net7012),
    .C(net6970),
    .A(_02780_),
    .Y(_10537_));
 sg13g2_o21ai_1 _24150_ (.B1(_10537_),
    .Y(_10538_),
    .A1(net7012),
    .A2(net6904));
 sg13g2_a21oi_1 _24151_ (.A1(net7012),
    .A2(net6878),
    .Y(_10539_),
    .B1(_02780_));
 sg13g2_a21oi_1 _24152_ (.A1(net6911),
    .A2(_10538_),
    .Y(_10540_),
    .B1(_10539_));
 sg13g2_nor2_1 _24153_ (.A(net6754),
    .B(_09864_),
    .Y(_10541_));
 sg13g2_nor3_1 _24154_ (.A(net6799),
    .B(_10048_),
    .C(_10541_),
    .Y(_10542_));
 sg13g2_a21oi_1 _24155_ (.A1(net6799),
    .A2(_09878_),
    .Y(_10543_),
    .B1(_10542_));
 sg13g2_a21oi_1 _24156_ (.A1(net6798),
    .A2(_09432_),
    .Y(_10544_),
    .B1(net6755));
 sg13g2_o21ai_1 _24157_ (.B1(_10544_),
    .Y(_10545_),
    .A1(_09403_),
    .A2(_09489_));
 sg13g2_a22oi_1 _24158_ (.Y(_10546_),
    .B1(_10545_),
    .B2(_10272_),
    .A2(_10543_),
    .A1(net6963));
 sg13g2_a221oi_1 _24159_ (.B2(net7293),
    .C1(_10540_),
    .B1(_10546_),
    .A1(net6983),
    .Y(_10547_),
    .A2(net6607));
 sg13g2_or2_1 _24160_ (.X(_10548_),
    .B(_10547_),
    .A(net7382));
 sg13g2_a22oi_1 _24161_ (.Y(_10549_),
    .B1(net6865),
    .B2(_00124_),
    .A2(net6834),
    .A1(_00188_));
 sg13g2_nand2b_1 _24162_ (.Y(_10550_),
    .B(net6708),
    .A_N(_10549_));
 sg13g2_a22oi_1 _24163_ (.Y(_10551_),
    .B1(net6865),
    .B2(_00160_),
    .A2(net6834),
    .A1(_00224_));
 sg13g2_o21ai_1 _24164_ (.B1(_10550_),
    .Y(_10552_),
    .A1(net6649),
    .A2(_10551_));
 sg13g2_a22oi_1 _24165_ (.Y(_10553_),
    .B1(net6671),
    .B2(_00516_),
    .A2(net6705),
    .A1(_00393_));
 sg13g2_nand2_1 _24166_ (.Y(_10554_),
    .A(_00360_),
    .B(net6699));
 sg13g2_a21oi_1 _24167_ (.A1(_00410_),
    .A2(_09570_),
    .Y(_10555_),
    .B1(net6683));
 sg13g2_a22oi_1 _24168_ (.Y(_10556_),
    .B1(_09567_),
    .B2(_00322_),
    .A2(_09566_),
    .A1(_00290_));
 sg13g2_a22oi_1 _24169_ (.Y(_10557_),
    .B1(net6677),
    .B2(_00485_),
    .A2(_06886_),
    .A1(net361));
 sg13g2_a22oi_1 _24170_ (.Y(_10558_),
    .B1(_10526_),
    .B2(net7518),
    .A2(net7594),
    .A1(_00726_));
 sg13g2_nand3_1 _24171_ (.B(_10556_),
    .C(_10557_),
    .A(_10555_),
    .Y(_10559_));
 sg13g2_a221oi_1 _24172_ (.B2(_00258_),
    .C1(_10559_),
    .B1(net6687),
    .A1(net427),
    .Y(_10560_),
    .A2(_09560_));
 sg13g2_nand3_1 _24173_ (.B(_10554_),
    .C(_10560_),
    .A(_10553_),
    .Y(_10561_));
 sg13g2_a21oi_1 _24174_ (.A1(net6795),
    .A2(_10552_),
    .Y(_10562_),
    .B1(_10561_));
 sg13g2_nand2_1 _24175_ (.Y(_10563_),
    .A(_01653_),
    .B(net7289));
 sg13g2_nand4_1 _24176_ (.B(_10548_),
    .C(_10562_),
    .A(net6548),
    .Y(_10564_),
    .D(_10563_));
 sg13g2_a21o_1 _24177_ (.A2(_08742_),
    .A1(net6635),
    .B1(_10564_),
    .X(_10565_));
 sg13g2_o21ai_1 _24178_ (.B1(net7714),
    .Y(_10566_),
    .A1(net7533),
    .A2(_10523_));
 sg13g2_a21oi_1 _24179_ (.A1(net5955),
    .A2(net7087),
    .Y(_10567_),
    .B1(_10565_));
 sg13g2_nand2_1 _24180_ (.Y(_10568_),
    .A(net7643),
    .B(_09374_));
 sg13g2_mux2_1 _24181_ (.A0(net326),
    .A1(_02005_),
    .S(net7652),
    .X(_10569_));
 sg13g2_o21ai_1 _24182_ (.B1(_10568_),
    .Y(_10570_),
    .A1(net7643),
    .A2(_10569_));
 sg13g2_o21ai_1 _24183_ (.B1(net6463),
    .Y(_10571_),
    .A1(net7663),
    .A2(_10570_));
 sg13g2_nand2b_1 _24184_ (.Y(_10572_),
    .B(_10571_),
    .A_N(net5905));
 sg13g2_o21ai_1 _24185_ (.B1(_10536_),
    .Y(_10573_),
    .A1(net6018),
    .A2(net5837));
 sg13g2_nand2_1 _24186_ (.Y(_10574_),
    .A(_01575_),
    .B(net6386));
 sg13g2_a21o_1 _24187_ (.A2(_10558_),
    .A1(net7533),
    .B1(_10566_),
    .X(_10575_));
 sg13g2_nand3_1 _24188_ (.B(net7013),
    .C(net6970),
    .A(_02715_),
    .Y(_10576_));
 sg13g2_o21ai_1 _24189_ (.B1(_10576_),
    .Y(_10577_),
    .A1(net7013),
    .A2(net6904));
 sg13g2_a21oi_1 _24190_ (.A1(net7013),
    .A2(net6878),
    .Y(_10578_),
    .B1(_02715_));
 sg13g2_a21oi_1 _24191_ (.A1(net6911),
    .A2(_10577_),
    .Y(_10579_),
    .B1(_10578_));
 sg13g2_a21oi_1 _24192_ (.A1(net6983),
    .A2(net6608),
    .Y(_10580_),
    .B1(_10579_));
 sg13g2_nand4_1 _24193_ (.B(_10477_),
    .C(_10492_),
    .A(_10438_),
    .Y(_10581_),
    .D(_10575_));
 sg13g2_nand3_1 _24194_ (.B(_01652_),
    .C(net7382),
    .A(net7923),
    .Y(_10582_));
 sg13g2_o21ai_1 _24195_ (.B1(_10582_),
    .Y(_10583_),
    .A1(net7382),
    .A2(_10580_));
 sg13g2_and2_1 _24196_ (.A(net6803),
    .B(_09796_),
    .X(_10584_));
 sg13g2_a21oi_1 _24197_ (.A1(net6798),
    .A2(_09785_),
    .Y(_10585_),
    .B1(_10584_));
 sg13g2_nand2_1 _24198_ (.Y(_10586_),
    .A(net6753),
    .B(_09934_));
 sg13g2_o21ai_1 _24199_ (.B1(_10586_),
    .Y(_10587_),
    .A1(net6753),
    .A2(_10585_));
 sg13g2_nor2_1 _24200_ (.A(net6754),
    .B(_09920_),
    .Y(_10588_));
 sg13g2_nor2_1 _24201_ (.A(_10273_),
    .B(_10588_),
    .Y(_10589_));
 sg13g2_nor2_1 _24202_ (.A(_08205_),
    .B(_10589_),
    .Y(_10590_));
 sg13g2_o21ai_1 _24203_ (.B1(_10590_),
    .Y(_10591_),
    .A1(net6955),
    .A2(_10587_));
 sg13g2_a22oi_1 _24204_ (.Y(_10592_),
    .B1(net6704),
    .B2(net426),
    .A2(net6705),
    .A1(_00392_));
 sg13g2_nand2_1 _24205_ (.Y(_10593_),
    .A(_00359_),
    .B(net6699));
 sg13g2_a21oi_1 _24206_ (.A1(_00289_),
    .A2(net6696),
    .Y(_10594_),
    .B1(net6683));
 sg13g2_a22oi_1 _24207_ (.Y(_10595_),
    .B1(net6680),
    .B2(_00409_),
    .A2(net6691),
    .A1(_00321_));
 sg13g2_a22oi_1 _24208_ (.Y(_10596_),
    .B1(net6676),
    .B2(_00484_),
    .A2(net6780),
    .A1(net360));
 sg13g2_nand3_1 _24209_ (.B(_10595_),
    .C(_10596_),
    .A(_10594_),
    .Y(_10597_));
 sg13g2_a221oi_1 _24210_ (.B2(_00515_),
    .C1(_10597_),
    .B1(net6671),
    .A1(_00257_),
    .Y(_10598_),
    .A2(net6686));
 sg13g2_nand3_1 _24211_ (.B(_10593_),
    .C(_10598_),
    .A(_10592_),
    .Y(_10599_));
 sg13g2_a22oi_1 _24212_ (.Y(_10600_),
    .B1(net6865),
    .B2(_00159_),
    .A2(net6834),
    .A1(_00223_));
 sg13g2_a22oi_1 _24213_ (.Y(_10601_),
    .B1(net6866),
    .B2(_00123_),
    .A2(net6836),
    .A1(_00187_));
 sg13g2_nand2b_1 _24214_ (.Y(_10602_),
    .B(net6713),
    .A_N(_10601_));
 sg13g2_o21ai_1 _24215_ (.B1(_10602_),
    .Y(_10603_),
    .A1(net6649),
    .A2(_10600_));
 sg13g2_a21oi_1 _24216_ (.A1(net6795),
    .A2(_10603_),
    .Y(_10604_),
    .B1(_10599_));
 sg13g2_nand2_1 _24217_ (.Y(_10605_),
    .A(_00100_),
    .B(net7082));
 sg13g2_nand4_1 _24218_ (.B(_10591_),
    .C(_10604_),
    .A(net6550),
    .Y(_10606_),
    .D(_10605_));
 sg13g2_or2_1 _24219_ (.X(_10607_),
    .B(_10606_),
    .A(_10583_));
 sg13g2_mux4_1 _24220_ (.S0(net7777),
    .A0(_01065_),
    .A1(_01100_),
    .A2(_01135_),
    .A3(_01171_),
    .S1(net7728),
    .X(_10608_));
 sg13g2_a21oi_1 _24221_ (.A1(net5969),
    .A2(net7088),
    .Y(_10609_),
    .B1(_10607_));
 sg13g2_nand2_1 _24222_ (.Y(_10610_),
    .A(net7647),
    .B(_09908_));
 sg13g2_mux2_1 _24223_ (.A0(net325),
    .A1(_02004_),
    .S(net7651),
    .X(_10611_));
 sg13g2_nand2b_1 _24224_ (.Y(_10612_),
    .B(net7433),
    .A_N(_10608_));
 sg13g2_o21ai_1 _24225_ (.B1(_10610_),
    .Y(_10613_),
    .A1(net7647),
    .A2(_10611_));
 sg13g2_o21ai_1 _24226_ (.B1(net6464),
    .Y(_10614_),
    .A1(net7663),
    .A2(_10613_));
 sg13g2_nand2b_1 _24227_ (.Y(_10615_),
    .B(_10614_),
    .A_N(net5932));
 sg13g2_o21ai_1 _24228_ (.B1(_10574_),
    .Y(_10616_),
    .A1(net6018),
    .A2(net5900));
 sg13g2_nand2_1 _24229_ (.Y(_10617_),
    .A(_01574_),
    .B(net6386));
 sg13g2_nand3_1 _24230_ (.B(net7014),
    .C(net6971),
    .A(_02653_),
    .Y(_10618_));
 sg13g2_o21ai_1 _24231_ (.B1(_10618_),
    .Y(_10619_),
    .A1(net7014),
    .A2(net6904));
 sg13g2_a21oi_1 _24232_ (.A1(net7014),
    .A2(net6878),
    .Y(_10620_),
    .B1(_02653_));
 sg13g2_a21oi_1 _24233_ (.A1(net6910),
    .A2(_10619_),
    .Y(_10621_),
    .B1(_10620_));
 sg13g2_a21oi_1 _24234_ (.A1(net6983),
    .A2(net6609),
    .Y(_10622_),
    .B1(_10621_));
 sg13g2_mux2_1 _24235_ (.A0(_09714_),
    .A1(_09736_),
    .S(_09402_),
    .X(_10623_));
 sg13g2_mux2_1 _24236_ (.A0(_09983_),
    .A1(_10623_),
    .S(net6757),
    .X(_10624_));
 sg13g2_nor2_1 _24237_ (.A(net6954),
    .B(_10624_),
    .Y(_10625_));
 sg13g2_nor2_1 _24238_ (.A(_09406_),
    .B(_09979_),
    .Y(_10626_));
 sg13g2_o21ai_1 _24239_ (.B1(net7293),
    .Y(_10627_),
    .A1(_10273_),
    .A2(_10626_));
 sg13g2_o21ai_1 _24240_ (.B1(_10622_),
    .Y(_10628_),
    .A1(_10625_),
    .A2(_10627_));
 sg13g2_a22oi_1 _24241_ (.Y(_10629_),
    .B1(net6866),
    .B2(_00122_),
    .A2(net6836),
    .A1(_00186_));
 sg13g2_nand2b_1 _24242_ (.Y(_10630_),
    .B(net6708),
    .A_N(_10629_));
 sg13g2_a22oi_1 _24243_ (.Y(_10631_),
    .B1(net6866),
    .B2(_00157_),
    .A2(net6836),
    .A1(_00221_));
 sg13g2_o21ai_1 _24244_ (.B1(_10630_),
    .Y(_10632_),
    .A1(net6649),
    .A2(_10631_));
 sg13g2_a22oi_1 _24245_ (.Y(_10633_),
    .B1(net6676),
    .B2(_00483_),
    .A2(net6780),
    .A1(net359));
 sg13g2_a21oi_1 _24246_ (.A1(_00288_),
    .A2(net6698),
    .Y(_10634_),
    .B1(net6683));
 sg13g2_a22oi_1 _24247_ (.Y(_10635_),
    .B1(net6680),
    .B2(_00408_),
    .A2(_09567_),
    .A1(_00320_));
 sg13g2_nand3_1 _24248_ (.B(_10634_),
    .C(_10635_),
    .A(_10633_),
    .Y(_10636_));
 sg13g2_a221oi_1 _24249_ (.B2(_00514_),
    .C1(_10636_),
    .B1(net6672),
    .A1(_00472_),
    .Y(_10637_),
    .A2(_09547_));
 sg13g2_a22oi_1 _24250_ (.Y(_10638_),
    .B1(net6699),
    .B2(_00358_),
    .A2(net6704),
    .A1(net425));
 sg13g2_a22oi_1 _24251_ (.Y(_10639_),
    .B1(net6686),
    .B2(_00256_),
    .A2(net6705),
    .A1(_00391_));
 sg13g2_nand3_1 _24252_ (.B(_10638_),
    .C(_10639_),
    .A(_10637_),
    .Y(_10640_));
 sg13g2_a21oi_1 _24253_ (.A1(net6795),
    .A2(_10632_),
    .Y(_10641_),
    .B1(_10640_));
 sg13g2_nand2_1 _24254_ (.Y(_10642_),
    .A(_01651_),
    .B(net7288));
 sg13g2_nand3_1 _24255_ (.B(_10641_),
    .C(_10642_),
    .A(net6548),
    .Y(_10643_));
 sg13g2_a221oi_1 _24256_ (.B2(net7367),
    .C1(_10643_),
    .B1(_10628_),
    .A1(_00089_),
    .Y(_10644_),
    .A2(net7082));
 sg13g2_mux4_1 _24257_ (.S0(net7777),
    .A0(_01206_),
    .A1(_01241_),
    .A2(_01276_),
    .A3(_01311_),
    .S1(net7728),
    .X(_10645_));
 sg13g2_or2_1 _24258_ (.X(_10646_),
    .B(_10645_),
    .A(net7587));
 sg13g2_nand2_1 _24259_ (.Y(_10647_),
    .A(_08926_),
    .B(_10644_));
 sg13g2_nand2_1 _24260_ (.Y(_10648_),
    .A(net7644),
    .B(_10011_));
 sg13g2_mux2_1 _24261_ (.A0(net324),
    .A1(_02003_),
    .S(net7655),
    .X(_10649_));
 sg13g2_o21ai_1 _24262_ (.B1(_10648_),
    .Y(_10650_),
    .A1(net7643),
    .A2(_10649_));
 sg13g2_o21ai_1 _24263_ (.B1(net6464),
    .Y(_10651_),
    .A1(net7663),
    .A2(_10650_));
 sg13g2_nand2_1 _24264_ (.Y(_10652_),
    .A(net5931),
    .B(_10651_));
 sg13g2_o21ai_1 _24265_ (.B1(_10617_),
    .Y(_10653_),
    .A1(net6018),
    .A2(net5895));
 sg13g2_nand2_1 _24266_ (.Y(_10654_),
    .A(_01573_),
    .B(net6388));
 sg13g2_nand2_1 _24267_ (.Y(_10655_),
    .A(net7642),
    .B(_10082_));
 sg13g2_mux2_1 _24268_ (.A0(net323),
    .A1(_02002_),
    .S(net7649),
    .X(_10656_));
 sg13g2_o21ai_1 _24269_ (.B1(_10655_),
    .Y(_10657_),
    .A1(net7642),
    .A2(_10656_));
 sg13g2_o21ai_1 _24270_ (.B1(net6465),
    .Y(_10658_),
    .A1(_00007_),
    .A2(_10657_));
 sg13g2_nand2_1 _24271_ (.Y(_10659_),
    .A(net6982),
    .B(net6610));
 sg13g2_mux2_1 _24272_ (.A0(_01417_),
    .A1(_01452_),
    .S(net7778),
    .X(_10660_));
 sg13g2_nand3_1 _24273_ (.B(net7015),
    .C(net6971),
    .A(_02586_),
    .Y(_10661_));
 sg13g2_o21ai_1 _24274_ (.B1(_10661_),
    .Y(_10662_),
    .A1(net7015),
    .A2(net6905));
 sg13g2_a21oi_1 _24275_ (.A1(net7015),
    .A2(net6879),
    .Y(_10663_),
    .B1(_02586_));
 sg13g2_a21oi_1 _24276_ (.A1(net6912),
    .A2(_10662_),
    .Y(_10664_),
    .B1(_10663_));
 sg13g2_nor3_1 _24277_ (.A(net7585),
    .B(_08464_),
    .C(_10660_),
    .Y(_10665_));
 sg13g2_a22oi_1 _24278_ (.Y(_10666_),
    .B1(net6866),
    .B2(_00121_),
    .A2(net6836),
    .A1(_00185_));
 sg13g2_nand2b_1 _24279_ (.Y(_10667_),
    .B(net6708),
    .A_N(_10666_));
 sg13g2_a22oi_1 _24280_ (.Y(_10668_),
    .B1(net6866),
    .B2(_00156_),
    .A2(net6836),
    .A1(_00220_));
 sg13g2_o21ai_1 _24281_ (.B1(_10667_),
    .Y(_10669_),
    .A1(net6649),
    .A2(_10668_));
 sg13g2_a22oi_1 _24282_ (.Y(_10670_),
    .B1(_09556_),
    .B2(net419),
    .A2(_09551_),
    .A1(_00482_));
 sg13g2_or2_1 _24283_ (.X(_10671_),
    .B(_10670_),
    .A(_09559_));
 sg13g2_a21oi_1 _24284_ (.A1(_00319_),
    .A2(net6694),
    .Y(_10672_),
    .B1(net6682));
 sg13g2_a22oi_1 _24285_ (.Y(_10673_),
    .B1(net6681),
    .B2(_00407_),
    .A2(_09566_),
    .A1(_00287_));
 sg13g2_nand2_1 _24286_ (.Y(_10674_),
    .A(_10672_),
    .B(_10673_));
 sg13g2_a21oi_1 _24287_ (.A1(net358),
    .A2(net6779),
    .Y(_10675_),
    .B1(_10674_));
 sg13g2_a22oi_1 _24288_ (.Y(_10676_),
    .B1(net6687),
    .B2(_00255_),
    .A2(net6706),
    .A1(_00382_));
 sg13g2_a22oi_1 _24289_ (.Y(_10677_),
    .B1(_10065_),
    .B2(_00513_),
    .A2(net6702),
    .A1(_00357_));
 sg13g2_nand4_1 _24290_ (.B(_10675_),
    .C(_10676_),
    .A(_10671_),
    .Y(_10678_),
    .D(_10677_));
 sg13g2_a21oi_1 _24291_ (.A1(net6796),
    .A2(_10669_),
    .Y(_10679_),
    .B1(_10678_));
 sg13g2_nor2b_1 _24292_ (.A(_10664_),
    .B_N(_10679_),
    .Y(_10680_));
 sg13g2_mux2_1 _24293_ (.A0(_01347_),
    .A1(_01382_),
    .S(net7778),
    .X(_10681_));
 sg13g2_nor3_1 _24294_ (.A(net7585),
    .B(_08503_),
    .C(_10681_),
    .Y(_10682_));
 sg13g2_a21o_1 _24295_ (.A2(_10680_),
    .A1(_10659_),
    .B1(net7378),
    .X(_10683_));
 sg13g2_nor2_1 _24296_ (.A(_09405_),
    .B(_10047_),
    .Y(_10684_));
 sg13g2_mux2_1 _24297_ (.A0(_09630_),
    .A1(_09635_),
    .S(_09403_),
    .X(_10685_));
 sg13g2_a21oi_1 _24298_ (.A1(net6756),
    .A2(_10685_),
    .Y(_10686_),
    .B1(_10684_));
 sg13g2_nand2_1 _24299_ (.Y(_10687_),
    .A(net6964),
    .B(_10686_));
 sg13g2_o21ai_1 _24300_ (.B1(_10272_),
    .Y(_10688_),
    .A1(_09406_),
    .A2(_10031_));
 sg13g2_nand3_1 _24301_ (.B(_10687_),
    .C(_10688_),
    .A(net7294),
    .Y(_10689_));
 sg13g2_and3_1 _24302_ (.X(_10690_),
    .A(_00078_),
    .B(_08708_),
    .C(_08721_));
 sg13g2_a221oi_1 _24303_ (.B2(_00085_),
    .C1(_10690_),
    .B1(_08709_),
    .A1(_01650_),
    .Y(_10691_),
    .A2(_08661_));
 sg13g2_nand3_1 _24304_ (.B(_10689_),
    .C(net5967),
    .A(_10683_),
    .Y(_10692_));
 sg13g2_o21ai_1 _24305_ (.B1(_10658_),
    .Y(_10693_),
    .A1(_09365_),
    .A2(net5930));
 sg13g2_o21ai_1 _24306_ (.B1(_10654_),
    .Y(_10694_),
    .A1(net6388),
    .A2(net5891));
 sg13g2_o21ai_1 _24307_ (.B1(net6961),
    .Y(_10695_),
    .A1(_09406_),
    .A2(_10031_));
 sg13g2_nand2_1 _24308_ (.Y(_10696_),
    .A(net6954),
    .B(_10686_));
 sg13g2_nand3_1 _24309_ (.B(_10695_),
    .C(_10696_),
    .A(net7294),
    .Y(_10697_));
 sg13g2_and2_1 _24310_ (.A(net6612),
    .B(net6902),
    .X(_10698_));
 sg13g2_nand2_1 _24311_ (.Y(_10699_),
    .A(_02535_),
    .B(_03730_));
 sg13g2_mux2_1 _24312_ (.A0(_01487_),
    .A1(_01523_),
    .S(net7778),
    .X(_10700_));
 sg13g2_nor3_1 _24313_ (.A(net7585),
    .B(_08485_),
    .C(_10700_),
    .Y(_10701_));
 sg13g2_a22oi_1 _24314_ (.Y(_10702_),
    .B1(net6866),
    .B2(_00155_),
    .A2(net6836),
    .A1(_00219_));
 sg13g2_a22oi_1 _24315_ (.Y(_10703_),
    .B1(net6866),
    .B2(_00120_),
    .A2(net6836),
    .A1(_00184_));
 sg13g2_mux4_1 _24316_ (.S0(net7648),
    .A0(net322),
    .A1(_02009_),
    .A2(_02001_),
    .A3(net345),
    .S1(net7656),
    .X(_10704_));
 sg13g2_a21oi_1 _24317_ (.A1(_06077_),
    .A2(_10704_),
    .Y(_10705_),
    .B1(_10100_));
 sg13g2_and2_1 _24318_ (.A(_09365_),
    .B(_10705_),
    .X(_10706_));
 sg13g2_mux2_1 _24319_ (.A0(net6971),
    .A1(_09388_),
    .S(_10699_),
    .X(_10707_));
 sg13g2_o21ai_1 _24320_ (.B1(net7365),
    .Y(_10708_),
    .A1(_02535_),
    .A2(_03730_));
 sg13g2_a21o_1 _24321_ (.A2(_10707_),
    .A1(net6912),
    .B1(_10708_),
    .X(_10709_));
 sg13g2_a221oi_1 _24322_ (.B2(_08956_),
    .C1(_10698_),
    .B1(_08708_),
    .A1(_01648_),
    .Y(_10710_),
    .A2(_08661_));
 sg13g2_nand2b_1 _24323_ (.Y(_10711_),
    .B(net6710),
    .A_N(_10703_));
 sg13g2_mux2_1 _24324_ (.A0(_01558_),
    .A1(_01593_),
    .S(net7778),
    .X(_10712_));
 sg13g2_nor2_1 _24325_ (.A(net7553),
    .B(_10712_),
    .Y(_10713_));
 sg13g2_a22oi_1 _24326_ (.Y(_10714_),
    .B1(_09583_),
    .B2(_00318_),
    .A2(net6824),
    .A1(net357));
 sg13g2_a22oi_1 _24327_ (.Y(_10715_),
    .B1(_10072_),
    .B2(_00512_),
    .A2(_09579_),
    .A1(_00254_));
 sg13g2_a22oi_1 _24328_ (.Y(_10716_),
    .B1(_09675_),
    .B2(\cs_registers_i.debug_ebreakm_o ),
    .A2(_09575_),
    .A1(_00406_));
 sg13g2_a22oi_1 _24329_ (.Y(_10717_),
    .B1(_09589_),
    .B2(_00481_),
    .A2(_09577_),
    .A1(_00286_));
 sg13g2_nand4_1 _24330_ (.B(_10715_),
    .C(_10716_),
    .A(_10714_),
    .Y(_10718_),
    .D(_10717_));
 sg13g2_and2_1 _24331_ (.A(_00356_),
    .B(_09582_),
    .X(_10719_));
 sg13g2_nand2b_1 _24332_ (.Y(_10720_),
    .B(net6707),
    .A_N(_10702_));
 sg13g2_a21oi_1 _24333_ (.A1(_10711_),
    .A2(_10720_),
    .Y(_10721_),
    .B1(_09538_));
 sg13g2_nor4_1 _24334_ (.A(_09585_),
    .B(_10718_),
    .C(_10719_),
    .D(_10721_),
    .Y(_10722_));
 sg13g2_and4_1 _24335_ (.A(_10697_),
    .B(_10709_),
    .C(net5887),
    .D(_10722_),
    .X(_10723_));
 sg13g2_a21oi_1 _24336_ (.A1(net6551),
    .A2(_10723_),
    .Y(_10724_),
    .B1(_10706_));
 sg13g2_mux2_1 _24337_ (.A0(net5775),
    .A1(_01572_),
    .S(net6387),
    .X(_10725_));
 sg13g2_nand2_1 _24338_ (.Y(_10726_),
    .A(_01571_),
    .B(net6388));
 sg13g2_a22oi_1 _24339_ (.Y(_10727_),
    .B1(_09614_),
    .B2(net330),
    .A2(net7475),
    .A1(net339));
 sg13g2_nand2b_1 _24340_ (.Y(_10728_),
    .B(net7661),
    .A_N(_10727_));
 sg13g2_a22oi_1 _24341_ (.Y(_10729_),
    .B1(_09616_),
    .B2(net321),
    .A2(_09377_),
    .A1(net344));
 sg13g2_or2_1 _24342_ (.X(_10730_),
    .B(_10729_),
    .A(_09378_));
 sg13g2_a22oi_1 _24343_ (.Y(_10731_),
    .B1(_09614_),
    .B2(_02000_),
    .A2(net7475),
    .A1(_02008_));
 sg13g2_or2_1 _24344_ (.X(_10732_),
    .B(_10731_),
    .A(net7664));
 sg13g2_nor4_1 _24345_ (.A(_10665_),
    .B(_10682_),
    .C(_10701_),
    .D(_10713_),
    .Y(_10733_));
 sg13g2_nor2_1 _24346_ (.A(net6552),
    .B(_10098_),
    .Y(_10734_));
 sg13g2_nand4_1 _24347_ (.B(_10730_),
    .C(_10732_),
    .A(_10728_),
    .Y(_10735_),
    .D(_10734_));
 sg13g2_mux2_1 _24348_ (.A0(_10624_),
    .A1(_10626_),
    .S(net6963),
    .X(_10736_));
 sg13g2_nand3_1 _24349_ (.B(net7016),
    .C(net6971),
    .A(_02477_),
    .Y(_10737_));
 sg13g2_o21ai_1 _24350_ (.B1(_10737_),
    .Y(_10738_),
    .A1(net7016),
    .A2(net6905));
 sg13g2_a21oi_1 _24351_ (.A1(net7016),
    .A2(net6879),
    .Y(_10739_),
    .B1(_02477_));
 sg13g2_a21oi_1 _24352_ (.A1(net6911),
    .A2(_10738_),
    .Y(_10740_),
    .B1(_10739_));
 sg13g2_a221oi_1 _24353_ (.B2(net7296),
    .C1(_10740_),
    .B1(_10736_),
    .A1(_08222_),
    .Y(_10741_),
    .A2(net6614));
 sg13g2_or2_1 _24354_ (.X(_10742_),
    .B(_10741_),
    .A(net7382));
 sg13g2_and2_1 _24355_ (.A(_00511_),
    .B(_10065_),
    .X(_10743_));
 sg13g2_a221oi_1 _24356_ (.B2(_00253_),
    .C1(_10743_),
    .B1(_09568_),
    .A1(_00355_),
    .Y(_10744_),
    .A2(_09563_));
 sg13g2_a21oi_1 _24357_ (.A1(_00317_),
    .A2(net6692),
    .Y(_10745_),
    .B1(net6685));
 sg13g2_a22oi_1 _24358_ (.Y(_10746_),
    .B1(net6681),
    .B2(_00405_),
    .A2(net6697),
    .A1(_00285_));
 sg13g2_a22oi_1 _24359_ (.Y(_10747_),
    .B1(net6674),
    .B2(_00480_),
    .A2(net6778),
    .A1(net356));
 sg13g2_nand4_1 _24360_ (.B(_10745_),
    .C(_10746_),
    .A(_10744_),
    .Y(_10748_),
    .D(_10747_));
 sg13g2_a22oi_1 _24361_ (.Y(_10749_),
    .B1(net6869),
    .B2(_00154_),
    .A2(net6839),
    .A1(_00218_));
 sg13g2_and4_1 _24362_ (.A(_10581_),
    .B(_10612_),
    .C(_10646_),
    .D(_10733_),
    .X(_10750_));
 sg13g2_a22oi_1 _24363_ (.Y(_10751_),
    .B1(net6866),
    .B2(_00119_),
    .A2(net6836),
    .A1(_00183_));
 sg13g2_nand2b_1 _24364_ (.Y(_10752_),
    .B(net6713),
    .A_N(_10751_));
 sg13g2_o21ai_1 _24365_ (.B1(_10752_),
    .Y(_10753_),
    .A1(net6651),
    .A2(_10749_));
 sg13g2_a21o_1 _24366_ (.A2(_10753_),
    .A1(net6796),
    .B1(_10748_),
    .X(_10754_));
 sg13g2_a21oi_1 _24367_ (.A1(_01647_),
    .A2(_09671_),
    .Y(_10755_),
    .B1(_10754_));
 sg13g2_nor2_1 _24368_ (.A(_08641_),
    .B(_10750_),
    .Y(_10756_));
 sg13g2_nand4_1 _24369_ (.B(net6550),
    .C(_10742_),
    .A(_08971_),
    .Y(_10757_),
    .D(_10755_));
 sg13g2_nand2_1 _24370_ (.Y(_10758_),
    .A(_10735_),
    .B(_10757_));
 sg13g2_o21ai_1 _24371_ (.B1(_10726_),
    .Y(_10759_),
    .A1(net6388),
    .A2(net5882));
 sg13g2_nand2_1 _24372_ (.Y(_10760_),
    .A(_01570_),
    .B(net6390));
 sg13g2_mux4_1 _24373_ (.S0(net7649),
    .A0(net320),
    .A1(net329),
    .A2(net337),
    .A3(net343),
    .S1(net7642),
    .X(_10761_));
 sg13g2_mux4_1 _24374_ (.S0(net7641),
    .A0(net320),
    .A1(_02007_),
    .A2(_01999_),
    .A3(net343),
    .S1(net7649),
    .X(_10762_));
 sg13g2_a22oi_1 _24375_ (.Y(_10763_),
    .B1(_10762_),
    .B2(net7628),
    .A2(_10761_),
    .A1(_01982_));
 sg13g2_mux2_1 _24376_ (.A0(_10587_),
    .A1(_10588_),
    .S(net6962),
    .X(_10764_));
 sg13g2_nand3_1 _24377_ (.B(net7017),
    .C(net6971),
    .A(_02401_),
    .Y(_10765_));
 sg13g2_o21ai_1 _24378_ (.B1(_10765_),
    .Y(_10766_),
    .A1(net7017),
    .A2(net6904));
 sg13g2_a21oi_1 _24379_ (.A1(net7017),
    .A2(net6878),
    .Y(_10767_),
    .B1(_02401_));
 sg13g2_a21oi_1 _24380_ (.A1(net6911),
    .A2(_10766_),
    .Y(_10768_),
    .B1(_10767_));
 sg13g2_a221oi_1 _24381_ (.B2(net7295),
    .C1(_10768_),
    .B1(_10764_),
    .A1(net6984),
    .Y(_10769_),
    .A2(net6599));
 sg13g2_or2_1 _24382_ (.X(_10770_),
    .B(_10769_),
    .A(net7382));
 sg13g2_a22oi_1 _24383_ (.Y(_10771_),
    .B1(net6690),
    .B2(_00316_),
    .A2(net6696),
    .A1(_00284_));
 sg13g2_inv_1 _24384_ (.Y(_10772_),
    .A(_10771_));
 sg13g2_o21ai_1 _24385_ (.B1(_08851_),
    .Y(_10773_),
    .A1(\id_stage_i.controller_i.instr_is_compressed_i ),
    .A2(_09363_));
 sg13g2_a221oi_1 _24386_ (.B2(_00510_),
    .C1(_10772_),
    .B1(net6672),
    .A1(_00404_),
    .Y(_10774_),
    .A2(net6679));
 sg13g2_a22oi_1 _24387_ (.Y(_10775_),
    .B1(_09568_),
    .B2(_00252_),
    .A2(_09563_),
    .A1(_00354_));
 sg13g2_a221oi_1 _24388_ (.B2(_00245_),
    .C1(net6685),
    .B1(net6673),
    .A1(_00479_),
    .Y(_10776_),
    .A2(net6674));
 sg13g2_nand2_1 _24389_ (.Y(_10777_),
    .A(net355),
    .B(net6777));
 sg13g2_nand4_1 _24390_ (.B(_10775_),
    .C(_10776_),
    .A(_10774_),
    .Y(_10778_),
    .D(_10777_));
 sg13g2_a22oi_1 _24391_ (.Y(_10779_),
    .B1(net6870),
    .B2(_00153_),
    .A2(net6839),
    .A1(_00217_));
 sg13g2_a22oi_1 _24392_ (.Y(_10780_),
    .B1(net6869),
    .B2(_00118_),
    .A2(net6838),
    .A1(_00182_));
 sg13g2_nand2b_1 _24393_ (.Y(_10781_),
    .B(net6712),
    .A_N(_10780_));
 sg13g2_o21ai_1 _24394_ (.B1(_10781_),
    .Y(_10782_),
    .A1(net6652),
    .A2(_10779_));
 sg13g2_a21oi_1 _24395_ (.A1(net6795),
    .A2(_10782_),
    .Y(_10783_),
    .B1(_10778_));
 sg13g2_nand2_1 _24396_ (.Y(_10784_),
    .A(_01646_),
    .B(_09671_));
 sg13g2_nand4_1 _24397_ (.B(_10770_),
    .C(_10783_),
    .A(net6550),
    .Y(_10785_),
    .D(_10784_));
 sg13g2_a21oi_1 _24398_ (.A1(net6058),
    .A2(net7088),
    .Y(_10786_),
    .B1(_10785_));
 sg13g2_a221oi_1 _24399_ (.B2(_01917_),
    .C1(_10773_),
    .B1(_09397_),
    .A1(net7699),
    .Y(_10787_),
    .A2(_08800_));
 sg13g2_nor2_1 _24400_ (.A(_10756_),
    .B(_10787_),
    .Y(_10788_));
 sg13g2_or2_1 _24401_ (.X(_10789_),
    .B(_10787_),
    .A(_10756_));
 sg13g2_a21o_1 _24402_ (.A2(_10763_),
    .A1(_10734_),
    .B1(_10786_),
    .X(_10790_));
 sg13g2_o21ai_1 _24403_ (.B1(_10760_),
    .Y(_10791_),
    .A1(net6390),
    .A2(net5928));
 sg13g2_nand2_1 _24404_ (.Y(_10792_),
    .A(_01569_),
    .B(net6390));
 sg13g2_mux4_1 _24405_ (.S0(net7653),
    .A0(net319),
    .A1(net328),
    .A2(net336),
    .A3(net342),
    .S1(net7646),
    .X(_10793_));
 sg13g2_mux4_1 _24406_ (.S0(net7646),
    .A0(net319),
    .A1(_02006_),
    .A2(_01998_),
    .A3(net342),
    .S1(net7653),
    .X(_10794_));
 sg13g2_a22oi_1 _24407_ (.Y(_10795_),
    .B1(_10794_),
    .B2(_06077_),
    .A2(_10793_),
    .A1(net7661));
 sg13g2_or2_1 _24408_ (.X(_10796_),
    .B(_10545_),
    .A(net6956));
 sg13g2_o21ai_1 _24409_ (.B1(_10796_),
    .Y(_10797_),
    .A1(net6963),
    .A2(_10543_));
 sg13g2_nand3_1 _24410_ (.B(net7018),
    .C(net6971),
    .A(_02326_),
    .Y(_10798_));
 sg13g2_o21ai_1 _24411_ (.B1(_10798_),
    .Y(_10799_),
    .A1(net7018),
    .A2(net6905));
 sg13g2_a21oi_1 _24412_ (.A1(net7018),
    .A2(net6879),
    .Y(_10800_),
    .B1(_02326_));
 sg13g2_a21oi_1 _24413_ (.A1(net6911),
    .A2(_10799_),
    .Y(_10801_),
    .B1(_10800_));
 sg13g2_a221oi_1 _24414_ (.B2(net7296),
    .C1(_10801_),
    .B1(_10797_),
    .A1(_08222_),
    .Y(_10802_),
    .A2(net6602));
 sg13g2_a21oi_1 _24415_ (.A1(net7923),
    .A2(_01645_),
    .Y(_10803_),
    .B1(net7368));
 sg13g2_a21o_1 _24416_ (.A2(_10802_),
    .A1(net7368),
    .B1(_10803_),
    .X(_10804_));
 sg13g2_a22oi_1 _24417_ (.Y(_10805_),
    .B1(net6676),
    .B2(_00478_),
    .A2(_09547_),
    .A1(_00474_));
 sg13g2_a22oi_1 _24418_ (.Y(_10806_),
    .B1(_09570_),
    .B2(_00403_),
    .A2(net6698),
    .A1(_00283_));
 sg13g2_a22oi_1 _24419_ (.Y(_10807_),
    .B1(net6673),
    .B2(\cs_registers_i.debug_ebreaku_o ),
    .A2(net6691),
    .A1(_00315_));
 sg13g2_mux2_1 _24420_ (.A0(_01236_),
    .A1(_01588_),
    .S(net7867),
    .X(_10808_));
 sg13g2_a22oi_1 _24421_ (.Y(_10809_),
    .B1(net6671),
    .B2(_00509_),
    .A2(net6778),
    .A1(net354));
 sg13g2_nand4_1 _24422_ (.B(_10806_),
    .C(_10807_),
    .A(_10805_),
    .Y(_10810_),
    .D(_10809_));
 sg13g2_a221oi_1 _24423_ (.B2(_00251_),
    .C1(_10147_),
    .B1(_09568_),
    .A1(_00353_),
    .Y(_10811_),
    .A2(_09563_));
 sg13g2_nand2b_1 _24424_ (.Y(_10812_),
    .B(_10811_),
    .A_N(_10810_));
 sg13g2_a22oi_1 _24425_ (.Y(_10813_),
    .B1(net6869),
    .B2(_00152_),
    .A2(net6838),
    .A1(_00216_));
 sg13g2_a22oi_1 _24426_ (.Y(_10814_),
    .B1(net6870),
    .B2(_00117_),
    .A2(net6838),
    .A1(_00181_));
 sg13g2_nand2b_1 _24427_ (.Y(_10815_),
    .B(net6712),
    .A_N(_10814_));
 sg13g2_o21ai_1 _24428_ (.B1(_10815_),
    .Y(_10816_),
    .A1(net6651),
    .A2(_10813_));
 sg13g2_a21oi_1 _24429_ (.A1(net6795),
    .A2(_10816_),
    .Y(_10817_),
    .B1(_10812_));
 sg13g2_nand2_1 _24430_ (.Y(_10818_),
    .A(_01645_),
    .B(net7082));
 sg13g2_nand4_1 _24431_ (.B(_10804_),
    .C(_10817_),
    .A(net6548),
    .Y(_10819_),
    .D(_10818_));
 sg13g2_a21oi_1 _24432_ (.A1(_00081_),
    .A2(net7087),
    .Y(_10820_),
    .B1(_10819_));
 sg13g2_a221oi_1 _24433_ (.B2(net7833),
    .C1(net7816),
    .B1(_10808_),
    .A1(_00884_),
    .Y(_10821_),
    .A2(net7527));
 sg13g2_a21o_1 _24434_ (.A2(_10795_),
    .A1(_10734_),
    .B1(net6016),
    .X(_10822_));
 sg13g2_o21ai_1 _24435_ (.B1(_10792_),
    .Y(_10823_),
    .A1(net6390),
    .A2(net5966));
 sg13g2_nand2_1 _24436_ (.Y(_10824_),
    .A(_01568_),
    .B(net6389));
 sg13g2_o21ai_1 _24437_ (.B1(net7293),
    .Y(_10825_),
    .A1(net6957),
    .A2(_10501_));
 sg13g2_mux2_1 _24438_ (.A0(_00662_),
    .A1(_00694_),
    .S(net7867),
    .X(_10826_));
 sg13g2_a21oi_1 _24439_ (.A1(net6957),
    .A2(_10498_),
    .Y(_10827_),
    .B1(_10825_));
 sg13g2_nand3_1 _24440_ (.B(net7019),
    .C(net6972),
    .A(net7031),
    .Y(_10828_));
 sg13g2_o21ai_1 _24441_ (.B1(_10828_),
    .Y(_10829_),
    .A1(net7019),
    .A2(net6906));
 sg13g2_a21oi_1 _24442_ (.A1(net7019),
    .A2(net6880),
    .Y(_10830_),
    .B1(net7032));
 sg13g2_nor2_1 _24443_ (.A(net7509),
    .B(_10826_),
    .Y(_10831_));
 sg13g2_a21oi_1 _24444_ (.A1(net6908),
    .A2(_10829_),
    .Y(_10832_),
    .B1(_10830_));
 sg13g2_a21o_1 _24445_ (.A2(net6621),
    .A1(net6984),
    .B1(_10832_),
    .X(_10833_));
 sg13g2_o21ai_1 _24446_ (.B1(net7365),
    .Y(_10834_),
    .A1(_10827_),
    .A2(_10833_));
 sg13g2_a22oi_1 _24447_ (.Y(_10835_),
    .B1(net6870),
    .B2(_00116_),
    .A2(net6838),
    .A1(_00180_));
 sg13g2_nand2b_1 _24448_ (.Y(_10836_),
    .B(net6710),
    .A_N(_10835_));
 sg13g2_a22oi_1 _24449_ (.Y(_10837_),
    .B1(net6869),
    .B2(_00151_),
    .A2(net6838),
    .A1(_00215_));
 sg13g2_o21ai_1 _24450_ (.B1(_10836_),
    .Y(_10838_),
    .A1(net6651),
    .A2(_10837_));
 sg13g2_a22oi_1 _24451_ (.Y(_10839_),
    .B1(_09661_),
    .B2(_00244_),
    .A2(net6698),
    .A1(_00282_));
 sg13g2_inv_1 _24452_ (.Y(_10840_),
    .A(_10839_));
 sg13g2_a221oi_1 _24453_ (.B2(_00250_),
    .C1(_10840_),
    .B1(net6687),
    .A1(_00314_),
    .Y(_10841_),
    .A2(net6691));
 sg13g2_a221oi_1 _24454_ (.B2(_00402_),
    .C1(net6685),
    .B1(net6678),
    .A1(_00473_),
    .Y(_10842_),
    .A2(_09547_));
 sg13g2_a22oi_1 _24455_ (.Y(_10843_),
    .B1(net6674),
    .B2(_00477_),
    .A2(net6778),
    .A1(net353));
 sg13g2_a22oi_1 _24456_ (.Y(_10844_),
    .B1(net6700),
    .B2(_00352_),
    .A2(net6706),
    .A1(_00388_));
 sg13g2_a22oi_1 _24457_ (.Y(_10845_),
    .B1(_10065_),
    .B2(_00508_),
    .A2(_09560_),
    .A1(net418));
 sg13g2_and2_1 _24458_ (.A(_10844_),
    .B(_10845_),
    .X(_10846_));
 sg13g2_nand4_1 _24459_ (.B(_10842_),
    .C(_10843_),
    .A(_10841_),
    .Y(_10847_),
    .D(_10846_));
 sg13g2_a21oi_1 _24460_ (.A1(net6796),
    .A2(_10838_),
    .Y(_10848_),
    .B1(_10847_));
 sg13g2_nand2_1 _24461_ (.Y(_10849_),
    .A(_01644_),
    .B(_09671_));
 sg13g2_nand4_1 _24462_ (.B(_10834_),
    .C(_10848_),
    .A(net6550),
    .Y(_10850_),
    .D(_10849_));
 sg13g2_mux2_1 _24463_ (.A0(_00726_),
    .A1(_00758_),
    .S(net7867),
    .X(_10851_));
 sg13g2_a21oi_1 _24464_ (.A1(_00080_),
    .A2(net7087),
    .Y(_10852_),
    .B1(_10850_));
 sg13g2_mux4_1 _24465_ (.S0(net7653),
    .A0(net318),
    .A1(net326),
    .A2(net335),
    .A3(net341),
    .S1(net7646),
    .X(_10853_));
 sg13g2_mux4_1 _24466_ (.S0(net7645),
    .A0(net318),
    .A1(_02005_),
    .A2(_01997_),
    .A3(net341),
    .S1(net7653),
    .X(_10854_));
 sg13g2_a22oi_1 _24467_ (.Y(_10855_),
    .B1(_10854_),
    .B2(_06077_),
    .A2(_10853_),
    .A1(net7661));
 sg13g2_o21ai_1 _24468_ (.B1(net7530),
    .Y(_10856_),
    .A1(net7521),
    .A2(_10851_));
 sg13g2_a21o_1 _24469_ (.A2(_10855_),
    .A1(_10734_),
    .B1(net6103),
    .X(_10857_));
 sg13g2_nor3_1 _24470_ (.A(_10821_),
    .B(_10831_),
    .C(_10856_),
    .Y(_10858_));
 sg13g2_o21ai_1 _24471_ (.B1(_10824_),
    .Y(_10859_),
    .A1(net6389),
    .A2(net6012));
 sg13g2_nand2_1 _24472_ (.Y(_10860_),
    .A(_01567_),
    .B(net6386));
 sg13g2_o21ai_1 _24473_ (.B1(net7385),
    .Y(_10861_),
    .A1(net7482),
    .A2(_01643_));
 sg13g2_nor2_1 _24474_ (.A(_09024_),
    .B(_10861_),
    .Y(_10862_));
 sg13g2_and2_1 _24475_ (.A(_00507_),
    .B(_10065_),
    .X(_10863_));
 sg13g2_a221oi_1 _24476_ (.B2(_00249_),
    .C1(_10863_),
    .B1(_09568_),
    .A1(_00351_),
    .Y(_10864_),
    .A2(_09563_));
 sg13g2_a21oi_1 _24477_ (.A1(_00281_),
    .A2(net6698),
    .Y(_10865_),
    .B1(net6685));
 sg13g2_a22oi_1 _24478_ (.Y(_10866_),
    .B1(_09570_),
    .B2(_00401_),
    .A2(net6690),
    .A1(_00313_));
 sg13g2_a22oi_1 _24479_ (.Y(_10867_),
    .B1(net6674),
    .B2(_00476_),
    .A2(net6777),
    .A1(net352));
 sg13g2_nand4_1 _24480_ (.B(_10865_),
    .C(_10866_),
    .A(_10864_),
    .Y(_10868_),
    .D(_10867_));
 sg13g2_a22oi_1 _24481_ (.Y(_10869_),
    .B1(net6869),
    .B2(_00150_),
    .A2(net6838),
    .A1(_00214_));
 sg13g2_a22oi_1 _24482_ (.Y(_10870_),
    .B1(net6870),
    .B2(_00115_),
    .A2(net6838),
    .A1(_00179_));
 sg13g2_nand2b_1 _24483_ (.Y(_10871_),
    .B(net6712),
    .A_N(_10870_));
 sg13g2_o21ai_1 _24484_ (.B1(_10871_),
    .Y(_10872_),
    .A1(net6651),
    .A2(_10869_));
 sg13g2_a21oi_1 _24485_ (.A1(net6796),
    .A2(_10872_),
    .Y(_10873_),
    .B1(_10868_));
 sg13g2_nand2_1 _24486_ (.Y(_10874_),
    .A(net6961),
    .B(_10459_));
 sg13g2_o21ai_1 _24487_ (.B1(_10874_),
    .Y(_10875_),
    .A1(net6961),
    .A2(_10460_));
 sg13g2_nand3_1 _24488_ (.B(net7020),
    .C(net6909),
    .A(_02172_),
    .Y(_10876_));
 sg13g2_nand2b_1 _24489_ (.Y(_10877_),
    .B(net7033),
    .A_N(net7020));
 sg13g2_nand3_1 _24490_ (.B(_10876_),
    .C(_10877_),
    .A(net6880),
    .Y(_10878_));
 sg13g2_nand3_1 _24491_ (.B(net7020),
    .C(_09389_),
    .A(_02172_),
    .Y(_10879_));
 sg13g2_nand2_1 _24492_ (.Y(_10880_),
    .A(_10878_),
    .B(_10879_));
 sg13g2_a21oi_1 _24493_ (.A1(net7294),
    .A2(_10875_),
    .Y(_10881_),
    .B1(_10880_));
 sg13g2_a21oi_1 _24494_ (.A1(net6622),
    .A2(_09994_),
    .Y(_10882_),
    .B1(_09365_));
 sg13g2_nand3_1 _24495_ (.B(_10881_),
    .C(_10882_),
    .A(_10873_),
    .Y(_10883_));
 sg13g2_mux2_1 _24496_ (.A0(_01276_),
    .A1(_01311_),
    .S(net7863),
    .X(_10884_));
 sg13g2_nor2_1 _24497_ (.A(net7524),
    .B(_10884_),
    .Y(_10885_));
 sg13g2_nand2_1 _24498_ (.Y(_10886_),
    .A(net7644),
    .B(_10305_));
 sg13g2_o21ai_1 _24499_ (.B1(_10886_),
    .Y(_10887_),
    .A1(net7648),
    .A2(_10303_));
 sg13g2_mux2_1 _24500_ (.A0(_01065_),
    .A1(_01100_),
    .S(net7863),
    .X(_10888_));
 sg13g2_mux4_1 _24501_ (.S0(net7647),
    .A0(net317),
    .A1(_02004_),
    .A2(_01996_),
    .A3(net338),
    .S1(net7651),
    .X(_10889_));
 sg13g2_a221oi_1 _24502_ (.B2(_06077_),
    .C1(_10098_),
    .B1(_10889_),
    .A1(net7661),
    .Y(_10890_),
    .A2(_10887_));
 sg13g2_nor2_1 _24503_ (.A(_10182_),
    .B(_10888_),
    .Y(_10891_));
 sg13g2_nand2_1 _24504_ (.Y(_10892_),
    .A(_09365_),
    .B(_10890_));
 sg13g2_o21ai_1 _24505_ (.B1(_10892_),
    .Y(_10893_),
    .A1(_10862_),
    .A2(_10883_));
 sg13g2_o21ai_1 _24506_ (.B1(_10860_),
    .Y(_10894_),
    .A1(_10095_),
    .A2(net5958));
 sg13g2_nand2_1 _24507_ (.Y(_10895_),
    .A(_01566_),
    .B(net6043));
 sg13g2_o21ai_1 _24508_ (.B1(_10895_),
    .Y(_10896_),
    .A1(net6043),
    .A2(net5864));
 sg13g2_nand2_1 _24509_ (.Y(_10897_),
    .A(_01565_),
    .B(net6389));
 sg13g2_nand2_1 _24510_ (.Y(_10898_),
    .A(net6962),
    .B(_10424_));
 sg13g2_o21ai_1 _24511_ (.B1(_10898_),
    .Y(_10899_),
    .A1(net6962),
    .A2(_10423_));
 sg13g2_nand3b_1 _24512_ (.B(net7021),
    .C(_09390_),
    .Y(_10900_),
    .A_N(_02105_));
 sg13g2_o21ai_1 _24513_ (.B1(_10900_),
    .Y(_10901_),
    .A1(net7021),
    .A2(_09387_));
 sg13g2_nand2_1 _24514_ (.Y(_10902_),
    .A(net7021),
    .B(net6880));
 sg13g2_a22oi_1 _24515_ (.Y(_10903_),
    .B1(_10902_),
    .B2(_02105_),
    .A2(_10901_),
    .A1(net6909));
 sg13g2_a221oi_1 _24516_ (.B2(net7296),
    .C1(_10903_),
    .B1(_10899_),
    .A1(net6984),
    .Y(_10904_),
    .A2(net6625));
 sg13g2_or2_1 _24517_ (.X(_10905_),
    .B(_10904_),
    .A(net7379));
 sg13g2_and2_1 _24518_ (.A(_00530_),
    .B(_10065_),
    .X(_10906_));
 sg13g2_a221oi_1 _24519_ (.B2(_00279_),
    .C1(_10906_),
    .B1(net6689),
    .A1(_00381_),
    .Y(_10907_),
    .A2(net6702));
 sg13g2_a21oi_1 _24520_ (.A1(_00343_),
    .A2(net6690),
    .Y(_10908_),
    .B1(net6685));
 sg13g2_a22oi_1 _24521_ (.Y(_10909_),
    .B1(_09570_),
    .B2(_00431_),
    .A2(net6696),
    .A1(_00311_));
 sg13g2_a22oi_1 _24522_ (.Y(_10910_),
    .B1(net6674),
    .B2(_00506_),
    .A2(net6778),
    .A1(net382));
 sg13g2_nand4_1 _24523_ (.B(_10908_),
    .C(_10909_),
    .A(_10907_),
    .Y(_10911_),
    .D(_10910_));
 sg13g2_a22oi_1 _24524_ (.Y(_10912_),
    .B1(net6869),
    .B2(_00149_),
    .A2(net6839),
    .A1(_00213_));
 sg13g2_a22oi_1 _24525_ (.Y(_10913_),
    .B1(net6869),
    .B2(_00177_),
    .A2(net6838),
    .A1(_00241_));
 sg13g2_nand2b_1 _24526_ (.Y(_10914_),
    .B(net6712),
    .A_N(_10913_));
 sg13g2_o21ai_1 _24527_ (.B1(_10914_),
    .Y(_10915_),
    .A1(net6651),
    .A2(_10912_));
 sg13g2_mux2_1 _24528_ (.A0(_01135_),
    .A1(_01171_),
    .S(net7863),
    .X(_10916_));
 sg13g2_a21oi_1 _24529_ (.A1(net6796),
    .A2(_10915_),
    .Y(_10917_),
    .B1(_10911_));
 sg13g2_nand2_1 _24530_ (.Y(_10918_),
    .A(_01642_),
    .B(_09671_));
 sg13g2_nand4_1 _24531_ (.B(_10905_),
    .C(_10917_),
    .A(net6549),
    .Y(_10919_),
    .D(_10918_));
 sg13g2_nor2_1 _24532_ (.A(net7456),
    .B(_10916_),
    .Y(_10920_));
 sg13g2_a21oi_1 _24533_ (.A1(_00111_),
    .A2(net7087),
    .Y(_10921_),
    .B1(_10919_));
 sg13g2_a22oi_1 _24534_ (.Y(_10922_),
    .B1(_09614_),
    .B2(_01995_),
    .A2(net7476),
    .A1(_02003_));
 sg13g2_nor2_1 _24535_ (.A(net7664),
    .B(_10922_),
    .Y(_10923_));
 sg13g2_a22oi_1 _24536_ (.Y(_10924_),
    .B1(_09616_),
    .B2(net347),
    .A2(_09377_),
    .A1(net327));
 sg13g2_nor2_1 _24537_ (.A(_09378_),
    .B(_10924_),
    .Y(_10925_));
 sg13g2_a22oi_1 _24538_ (.Y(_10926_),
    .B1(_09614_),
    .B2(net324),
    .A2(net7475),
    .A1(net333));
 sg13g2_nor2b_1 _24539_ (.A(_10926_),
    .B_N(net7661),
    .Y(_10927_));
 sg13g2_nor3_1 _24540_ (.A(_10923_),
    .B(_10925_),
    .C(_10927_),
    .Y(_10928_));
 sg13g2_a21o_1 _24541_ (.A2(_10928_),
    .A1(_10734_),
    .B1(net6102),
    .X(_10929_));
 sg13g2_o21ai_1 _24542_ (.B1(_10897_),
    .Y(_10930_),
    .A1(net6389),
    .A2(net6009));
 sg13g2_nand2_1 _24543_ (.Y(_10931_),
    .A(_01564_),
    .B(net6388));
 sg13g2_nor2_1 _24544_ (.A(_03695_),
    .B(net6906),
    .Y(_10932_));
 sg13g2_nor3_1 _24545_ (.A(_02032_),
    .B(net7022),
    .C(_09389_),
    .Y(_10933_));
 sg13g2_o21ai_1 _24546_ (.B1(net6908),
    .Y(_10934_),
    .A1(_10932_),
    .A2(_10933_));
 sg13g2_o21ai_1 _24547_ (.B1(_02032_),
    .Y(_10935_),
    .A1(net7022),
    .A2(_09393_));
 sg13g2_a221oi_1 _24548_ (.B2(_10935_),
    .C1(net7378),
    .B1(_10934_),
    .A1(net6982),
    .Y(_10936_),
    .A2(net6626));
 sg13g2_o21ai_1 _24549_ (.B1(net7294),
    .Y(_10937_),
    .A1(net6954),
    .A2(_10389_));
 sg13g2_a21o_1 _24550_ (.A2(_10386_),
    .A1(net6954),
    .B1(_10937_),
    .X(_10938_));
 sg13g2_mux2_1 _24551_ (.A0(_01206_),
    .A1(_01241_),
    .S(net7863),
    .X(_10939_));
 sg13g2_a221oi_1 _24552_ (.B2(_01641_),
    .C1(net7370),
    .B1(_09535_),
    .A1(_00110_),
    .Y(_10940_),
    .A2(_08739_));
 sg13g2_a21oi_1 _24553_ (.A1(_10936_),
    .A2(_10938_),
    .Y(_10941_),
    .B1(_10940_));
 sg13g2_a22oi_1 _24554_ (.Y(_10942_),
    .B1(net6870),
    .B2(_00176_),
    .A2(net6839),
    .A1(_00240_));
 sg13g2_a22oi_1 _24555_ (.Y(_10943_),
    .B1(net6870),
    .B2(_00148_),
    .A2(net6839),
    .A1(_00212_));
 sg13g2_o21ai_1 _24556_ (.B1(net7502),
    .Y(_10944_),
    .A1(net7504),
    .A2(_10939_));
 sg13g2_nor4_1 _24557_ (.A(_10885_),
    .B(_10891_),
    .C(_10920_),
    .D(_10944_),
    .Y(_10945_));
 sg13g2_a21o_1 _24558_ (.A2(_10065_),
    .A1(_00529_),
    .B1(_10147_),
    .X(_10946_));
 sg13g2_a221oi_1 _24559_ (.B2(_00278_),
    .C1(_10946_),
    .B1(_09568_),
    .A1(_00380_),
    .Y(_10947_),
    .A2(_09563_));
 sg13g2_a22oi_1 _24560_ (.Y(_10948_),
    .B1(net6678),
    .B2(_00430_),
    .A2(net6692),
    .A1(_00342_));
 sg13g2_a22oi_1 _24561_ (.Y(_10949_),
    .B1(net6673),
    .B2(_00248_),
    .A2(net6698),
    .A1(_00310_));
 sg13g2_a22oi_1 _24562_ (.Y(_10950_),
    .B1(net6674),
    .B2(_00505_),
    .A2(net6777),
    .A1(net381));
 sg13g2_nand4_1 _24563_ (.B(_10948_),
    .C(_10949_),
    .A(_10947_),
    .Y(_10951_),
    .D(_10950_));
 sg13g2_nand2b_1 _24564_ (.Y(_10952_),
    .B(net6712),
    .A_N(_10942_));
 sg13g2_o21ai_1 _24565_ (.B1(_10952_),
    .Y(_10953_),
    .A1(net6651),
    .A2(_10943_));
 sg13g2_a21oi_1 _24566_ (.A1(net6796),
    .A2(_10953_),
    .Y(_10954_),
    .B1(_10951_));
 sg13g2_mux2_1 _24567_ (.A0(_00854_),
    .A1(_00889_),
    .S(net7866),
    .X(_10955_));
 sg13g2_nand2_1 _24568_ (.Y(_10956_),
    .A(net6551),
    .B(_10954_));
 sg13g2_nand3_1 _24569_ (.B(_10189_),
    .C(_10955_),
    .A(net7546),
    .Y(_10957_));
 sg13g2_mux4_1 _24570_ (.S0(net7650),
    .A0(net346),
    .A1(net323),
    .A2(net332),
    .A3(net316),
    .S1(_01987_),
    .X(_10958_));
 sg13g2_mux4_1 _24571_ (.S0(net7642),
    .A0(net346),
    .A1(_02002_),
    .A2(_01994_),
    .A3(net316),
    .S1(net7649),
    .X(_10959_));
 sg13g2_a22oi_1 _24572_ (.Y(_10960_),
    .B1(_10959_),
    .B2(net7628),
    .A2(_10958_),
    .A1(_01982_));
 sg13g2_nand2_1 _24573_ (.Y(_10961_),
    .A(_10734_),
    .B(_10960_));
 sg13g2_o21ai_1 _24574_ (.B1(_10961_),
    .Y(_10962_),
    .A1(_10941_),
    .A2(_10956_));
 sg13g2_o21ai_1 _24575_ (.B1(_10931_),
    .Y(_10963_),
    .A1(net6388),
    .A2(net6002));
 sg13g2_nand2_1 _24576_ (.Y(_10964_),
    .A(_01563_),
    .B(net6391));
 sg13g2_o21ai_1 _24577_ (.B1(_10964_),
    .Y(_10965_),
    .A1(net6119),
    .A2(net6391));
 sg13g2_nand2_1 _24578_ (.Y(_10966_),
    .A(_01562_),
    .B(net6389));
 sg13g2_o21ai_1 _24579_ (.B1(_10966_),
    .Y(_10967_),
    .A1(net6030),
    .A2(net6389));
 sg13g2_nand2_1 _24580_ (.Y(_10968_),
    .A(_01561_),
    .B(net6391));
 sg13g2_o21ai_1 _24581_ (.B1(_10968_),
    .Y(_10969_),
    .A1(net6113),
    .A2(net6391));
 sg13g2_mux2_1 _24582_ (.A0(_00790_),
    .A1(_00822_),
    .S(net7866),
    .X(_10970_));
 sg13g2_nand2_1 _24583_ (.Y(_10971_),
    .A(_01560_),
    .B(net6391));
 sg13g2_o21ai_1 _24584_ (.B1(_10971_),
    .Y(_10972_),
    .A1(net6026),
    .A2(net6391));
 sg13g2_nand2_1 _24585_ (.Y(_10973_),
    .A(_01559_),
    .B(net6388));
 sg13g2_nand3_1 _24586_ (.B(_10179_),
    .C(_10970_),
    .A(net7546),
    .Y(_10974_));
 sg13g2_o21ai_1 _24587_ (.B1(_10973_),
    .Y(_10975_),
    .A1(net6054),
    .A2(net6388));
 sg13g2_nand2_1 _24588_ (.Y(_10976_),
    .A(_01558_),
    .B(net6393));
 sg13g2_o21ai_1 _24589_ (.B1(_10976_),
    .Y(_10977_),
    .A1(net6020),
    .A2(net6393));
 sg13g2_nand2_1 _24590_ (.Y(_10978_),
    .A(_01557_),
    .B(net6389));
 sg13g2_o21ai_1 _24591_ (.B1(_10978_),
    .Y(_10979_),
    .A1(net6106),
    .A2(net6389));
 sg13g2_and4_1 _24592_ (.A(net7806),
    .B(_01895_),
    .C(net7812),
    .D(_01893_),
    .X(_10980_));
 sg13g2_nand2_1 _24593_ (.Y(_10981_),
    .A(_01556_),
    .B(net6386));
 sg13g2_nand4_1 _24594_ (.B(net7808),
    .C(net7812),
    .A(net7806),
    .Y(_10982_),
    .D(_01893_));
 sg13g2_o21ai_1 _24595_ (.B1(_10981_),
    .Y(_10983_),
    .A1(net5867),
    .A2(net6018));
 sg13g2_nand4_1 _24596_ (.B(_06619_),
    .C(_06621_),
    .A(net7670),
    .Y(_10984_),
    .D(_09604_));
 sg13g2_nor2_1 _24597_ (.A(_06622_),
    .B(_09607_),
    .Y(_10985_));
 sg13g2_nand2_1 _24598_ (.Y(_10986_),
    .A(_06619_),
    .B(_10985_));
 sg13g2_nand2_1 _24599_ (.Y(_10987_),
    .A(_01555_),
    .B(net6361));
 sg13g2_o21ai_1 _24600_ (.B1(_10987_),
    .Y(_10988_),
    .A1(net8286),
    .A2(net6361));
 sg13g2_or4_1 _24601_ (.A(net7670),
    .B(net6467),
    .C(_09680_),
    .D(_09682_),
    .X(_10989_));
 sg13g2_nor2_1 _24602_ (.A(net7668),
    .B(_09603_),
    .Y(_10990_));
 sg13g2_nor3_1 _24603_ (.A(net7668),
    .B(_09603_),
    .C(_09682_),
    .Y(_10991_));
 sg13g2_nand2_1 _24604_ (.Y(_10992_),
    .A(net7474),
    .B(net6346));
 sg13g2_nand2_1 _24605_ (.Y(_10993_),
    .A(_01554_),
    .B(net6348));
 sg13g2_o21ai_1 _24606_ (.B1(_10993_),
    .Y(_10994_),
    .A1(net5863),
    .A2(net6348));
 sg13g2_nand2_1 _24607_ (.Y(_10995_),
    .A(_01553_),
    .B(net6348));
 sg13g2_nand2b_1 _24608_ (.Y(_10996_),
    .B(net6381),
    .A_N(net6351));
 sg13g2_o21ai_1 _24609_ (.B1(_10995_),
    .Y(_10997_),
    .A1(net5855),
    .A2(_10996_));
 sg13g2_mux2_1 _24610_ (.A0(_01558_),
    .A1(_01593_),
    .S(net7866),
    .X(_10998_));
 sg13g2_nand2_1 _24611_ (.Y(_10999_),
    .A(_01552_),
    .B(net6352));
 sg13g2_o21ai_1 _24612_ (.B1(_10999_),
    .Y(_11000_),
    .A1(net5808),
    .A2(net6101));
 sg13g2_nand2_1 _24613_ (.Y(_11001_),
    .A(_01551_),
    .B(net6349));
 sg13g2_nand2_1 _24614_ (.Y(_11002_),
    .A(_10980_),
    .B(_10998_));
 sg13g2_o21ai_1 _24615_ (.B1(_11001_),
    .Y(_11003_),
    .A1(net5850),
    .A2(net6351));
 sg13g2_nand2_1 _24616_ (.Y(_11004_),
    .A(_01550_),
    .B(net6350));
 sg13g2_o21ai_1 _24617_ (.B1(_11004_),
    .Y(_11005_),
    .A1(net5802),
    .A2(net6350));
 sg13g2_nand2_1 _24618_ (.Y(_11006_),
    .A(_01549_),
    .B(net6352));
 sg13g2_o21ai_1 _24619_ (.B1(_11006_),
    .Y(_11007_),
    .A1(net5795),
    .A2(_10992_));
 sg13g2_nand2_1 _24620_ (.Y(_11008_),
    .A(_01548_),
    .B(_10989_));
 sg13g2_nand2b_1 _24621_ (.Y(_11009_),
    .B(net6379),
    .A_N(_10989_));
 sg13g2_o21ai_1 _24622_ (.B1(_11008_),
    .Y(_11010_),
    .A1(net5917),
    .A2(_11009_));
 sg13g2_nand2_1 _24623_ (.Y(_11011_),
    .A(_01547_),
    .B(net6352));
 sg13g2_o21ai_1 _24624_ (.B1(_11011_),
    .Y(_11012_),
    .A1(net5791),
    .A2(net6101));
 sg13g2_nand2_1 _24625_ (.Y(_11013_),
    .A(_01546_),
    .B(net6347));
 sg13g2_nand2b_1 _24626_ (.Y(_11014_),
    .B(net6374),
    .A_N(net6347));
 sg13g2_o21ai_1 _24627_ (.B1(_11013_),
    .Y(_11015_),
    .A1(net5912),
    .A2(_11014_));
 sg13g2_nand2_1 _24628_ (.Y(_11016_),
    .A(_01545_),
    .B(net6352));
 sg13g2_mux2_1 _24629_ (.A0(_01487_),
    .A1(_01523_),
    .S(net7866),
    .X(_11017_));
 sg13g2_o21ai_1 _24630_ (.B1(_11016_),
    .Y(_11018_),
    .A1(net5778),
    .A2(_10992_));
 sg13g2_nand2_1 _24631_ (.Y(_11019_),
    .A(_01544_),
    .B(net6362));
 sg13g2_nand2b_1 _24632_ (.Y(_11020_),
    .B(net6382),
    .A_N(net6362));
 sg13g2_o21ai_1 _24633_ (.B1(_11019_),
    .Y(_11021_),
    .A1(net5854),
    .A2(_11020_));
 sg13g2_nand3_1 _24634_ (.B(_09150_),
    .C(_11017_),
    .A(net7515),
    .Y(_11022_));
 sg13g2_nand2_1 _24635_ (.Y(_11023_),
    .A(_01543_),
    .B(net6347));
 sg13g2_nand2b_1 _24636_ (.Y(_11024_),
    .B(net6366),
    .A_N(net6347));
 sg13g2_o21ai_1 _24637_ (.B1(_11023_),
    .Y(_11025_),
    .A1(net5910),
    .A2(_11024_));
 sg13g2_mux2_1 _24638_ (.A0(net5840),
    .A1(_01542_),
    .S(_10992_),
    .X(_11026_));
 sg13g2_nand2_1 _24639_ (.Y(_11027_),
    .A(_01541_),
    .B(net6355));
 sg13g2_o21ai_1 _24640_ (.B1(_11027_),
    .Y(_11028_),
    .A1(net5834),
    .A2(_10992_));
 sg13g2_nand2_1 _24641_ (.Y(_11029_),
    .A(_01540_),
    .B(net6352));
 sg13g2_o21ai_1 _24642_ (.B1(_11029_),
    .Y(_11030_),
    .A1(net5900),
    .A2(net6101));
 sg13g2_nand2_1 _24643_ (.Y(_11031_),
    .A(_01539_),
    .B(net6352));
 sg13g2_o21ai_1 _24644_ (.B1(_11031_),
    .Y(_11032_),
    .A1(net5895),
    .A2(net6101));
 sg13g2_nand2_1 _24645_ (.Y(_11033_),
    .A(_01538_),
    .B(net6353));
 sg13g2_o21ai_1 _24646_ (.B1(_11033_),
    .Y(_11034_),
    .A1(net5891),
    .A2(net6353));
 sg13g2_mux2_1 _24647_ (.A0(net5775),
    .A1(_01537_),
    .S(net6347),
    .X(_11035_));
 sg13g2_nand2_1 _24648_ (.Y(_11036_),
    .A(_01536_),
    .B(net6355));
 sg13g2_o21ai_1 _24649_ (.B1(_11036_),
    .Y(_11037_),
    .A1(net5882),
    .A2(net6353));
 sg13g2_nand2_1 _24650_ (.Y(_11038_),
    .A(_01535_),
    .B(net6351));
 sg13g2_o21ai_1 _24651_ (.B1(_11038_),
    .Y(_11039_),
    .A1(net5927),
    .A2(net6351));
 sg13g2_mux2_1 _24652_ (.A0(_01347_),
    .A1(_01382_),
    .S(net7866),
    .X(_11040_));
 sg13g2_nand2_1 _24653_ (.Y(_11041_),
    .A(_01534_),
    .B(net6350));
 sg13g2_o21ai_1 _24654_ (.B1(_11041_),
    .Y(_11042_),
    .A1(net5966),
    .A2(net6350));
 sg13g2_nand2_1 _24655_ (.Y(_11043_),
    .A(_01533_),
    .B(net6363));
 sg13g2_o21ai_1 _24656_ (.B1(_11043_),
    .Y(_11044_),
    .A1(net5804),
    .A2(net6000));
 sg13g2_nand3_1 _24657_ (.B(_10179_),
    .C(_11040_),
    .A(net7497),
    .Y(_11045_));
 sg13g2_nand2_1 _24658_ (.Y(_11046_),
    .A(_01532_),
    .B(net6354));
 sg13g2_o21ai_1 _24659_ (.B1(_11046_),
    .Y(_11047_),
    .A1(net6012),
    .A2(net6354));
 sg13g2_nand2_1 _24660_ (.Y(_11048_),
    .A(_01531_),
    .B(net6352));
 sg13g2_o21ai_1 _24661_ (.B1(_11048_),
    .Y(_11049_),
    .A1(net5958),
    .A2(_10992_));
 sg13g2_nand2_1 _24662_ (.Y(_11050_),
    .A(_01530_),
    .B(net6350));
 sg13g2_o21ai_1 _24663_ (.B1(_11050_),
    .Y(_11051_),
    .A1(net6009),
    .A2(net6350));
 sg13g2_nand2_1 _24664_ (.Y(_11052_),
    .A(_01529_),
    .B(net6354));
 sg13g2_o21ai_1 _24665_ (.B1(_11052_),
    .Y(_11053_),
    .A1(net6004),
    .A2(net6354));
 sg13g2_nand2_1 _24666_ (.Y(_11054_),
    .A(_01528_),
    .B(net6349));
 sg13g2_o21ai_1 _24667_ (.B1(_11054_),
    .Y(_11055_),
    .A1(net6118),
    .A2(net6349));
 sg13g2_nand2_1 _24668_ (.Y(_11056_),
    .A(_01527_),
    .B(net6350));
 sg13g2_o21ai_1 _24669_ (.B1(_11056_),
    .Y(_11057_),
    .A1(net6031),
    .A2(net6350));
 sg13g2_nand2_1 _24670_ (.Y(_11058_),
    .A(_01526_),
    .B(net6349));
 sg13g2_o21ai_1 _24671_ (.B1(_11058_),
    .Y(_11059_),
    .A1(net6113),
    .A2(net6349));
 sg13g2_mux2_1 _24672_ (.A0(_01417_),
    .A1(_01452_),
    .S(net7866),
    .X(_11060_));
 sg13g2_nand2_1 _24673_ (.Y(_11061_),
    .A(_01525_),
    .B(net6349));
 sg13g2_o21ai_1 _24674_ (.B1(_11061_),
    .Y(_11062_),
    .A1(net6027),
    .A2(net6349));
 sg13g2_nand2_1 _24675_ (.Y(_11063_),
    .A(_01524_),
    .B(net6353));
 sg13g2_nand3_1 _24676_ (.B(_10189_),
    .C(_11060_),
    .A(_09150_),
    .Y(_11064_));
 sg13g2_o21ai_1 _24677_ (.B1(_11063_),
    .Y(_11065_),
    .A1(_09601_),
    .A2(net6353));
 sg13g2_nand2_1 _24678_ (.Y(_11066_),
    .A(_01523_),
    .B(net6354));
 sg13g2_o21ai_1 _24679_ (.B1(_11066_),
    .Y(_11067_),
    .A1(net6020),
    .A2(net6354));
 sg13g2_nand2_1 _24680_ (.Y(_11068_),
    .A(_01522_),
    .B(net6361));
 sg13g2_o21ai_1 _24681_ (.B1(_11068_),
    .Y(_11069_),
    .A1(net5847),
    .A2(net6361));
 sg13g2_nand2_1 _24682_ (.Y(_11070_),
    .A(_01521_),
    .B(net6354));
 sg13g2_o21ai_1 _24683_ (.B1(_11070_),
    .Y(_11071_),
    .A1(net6106),
    .A2(net6354));
 sg13g2_nand2_1 _24684_ (.Y(_11072_),
    .A(_01520_),
    .B(net6352));
 sg13g2_o21ai_1 _24685_ (.B1(_11072_),
    .Y(_11073_),
    .A1(net5867),
    .A2(net6101));
 sg13g2_or4_1 _24686_ (.A(net7670),
    .B(net6467),
    .C(_09680_),
    .D(_10092_),
    .X(_11074_));
 sg13g2_nor3_1 _24687_ (.A(net7671),
    .B(_09603_),
    .C(_10092_),
    .Y(_11075_));
 sg13g2_nand2_1 _24688_ (.Y(_11076_),
    .A(net7474),
    .B(net6335));
 sg13g2_nand2_1 _24689_ (.Y(_11077_),
    .A(_01519_),
    .B(net6342));
 sg13g2_o21ai_1 _24690_ (.B1(_11077_),
    .Y(_11078_),
    .A1(net5863),
    .A2(net6342));
 sg13g2_nand2_1 _24691_ (.Y(_11079_),
    .A(_01518_),
    .B(net6342));
 sg13g2_nand2b_1 _24692_ (.Y(_11080_),
    .B(net6381),
    .A_N(net6345));
 sg13g2_o21ai_1 _24693_ (.B1(_11079_),
    .Y(_11081_),
    .A1(net5855),
    .A2(_11080_));
 sg13g2_nand2_1 _24694_ (.Y(_11082_),
    .A(_01517_),
    .B(net6337));
 sg13g2_o21ai_1 _24695_ (.B1(_11082_),
    .Y(_11083_),
    .A1(net5808),
    .A2(net6100));
 sg13g2_nand2_1 _24696_ (.Y(_11084_),
    .A(_01516_),
    .B(net6345));
 sg13g2_mux2_1 _24697_ (.A0(_00995_),
    .A1(_01030_),
    .S(net7866),
    .X(_11085_));
 sg13g2_o21ai_1 _24698_ (.B1(_11084_),
    .Y(_11086_),
    .A1(net5850),
    .A2(net6345));
 sg13g2_nand2_1 _24699_ (.Y(_11087_),
    .A(_01515_),
    .B(net6343));
 sg13g2_o21ai_1 _24700_ (.B1(_11087_),
    .Y(_11088_),
    .A1(net5802),
    .A2(net6343));
 sg13g2_nand3_1 _24701_ (.B(net7526),
    .C(_11085_),
    .A(net7546),
    .Y(_11089_));
 sg13g2_nand2_1 _24702_ (.Y(_11090_),
    .A(_01514_),
    .B(net6340));
 sg13g2_o21ai_1 _24703_ (.B1(_11090_),
    .Y(_11091_),
    .A1(net5795),
    .A2(_11076_));
 sg13g2_nand2_1 _24704_ (.Y(_11092_),
    .A(_01513_),
    .B(net6341));
 sg13g2_nand2b_1 _24705_ (.Y(_11093_),
    .B(net6379),
    .A_N(net6341));
 sg13g2_o21ai_1 _24706_ (.B1(_11092_),
    .Y(_11094_),
    .A1(net5917),
    .A2(_11093_));
 sg13g2_nand2_1 _24707_ (.Y(_11095_),
    .A(_01512_),
    .B(net6337));
 sg13g2_o21ai_1 _24708_ (.B1(_11095_),
    .Y(_11096_),
    .A1(net5789),
    .A2(net6100));
 sg13g2_nand2_1 _24709_ (.Y(_11097_),
    .A(_01511_),
    .B(net6358));
 sg13g2_o21ai_1 _24710_ (.B1(_11097_),
    .Y(_11098_),
    .A1(net5803),
    .A2(net6358));
 sg13g2_nand2_1 _24711_ (.Y(_11099_),
    .A(_01510_),
    .B(_11074_));
 sg13g2_nand2b_1 _24712_ (.Y(_11100_),
    .B(net6374),
    .A_N(_11074_));
 sg13g2_o21ai_1 _24713_ (.B1(_11099_),
    .Y(_11101_),
    .A1(net5912),
    .A2(_11100_));
 sg13g2_nand2_1 _24714_ (.Y(_11102_),
    .A(_01509_),
    .B(net6340));
 sg13g2_mux2_1 _24715_ (.A0(_00924_),
    .A1(_00959_),
    .S(net7866),
    .X(_11103_));
 sg13g2_o21ai_1 _24716_ (.B1(_11102_),
    .Y(_11104_),
    .A1(net5778),
    .A2(net6100));
 sg13g2_nand2_1 _24717_ (.Y(_11105_),
    .A(_01508_),
    .B(net6341));
 sg13g2_nand2b_1 _24718_ (.Y(_11106_),
    .B(net6366),
    .A_N(net6341));
 sg13g2_o21ai_1 _24719_ (.B1(_11105_),
    .Y(_11107_),
    .A1(net5910),
    .A2(_11106_));
 sg13g2_nand3_1 _24720_ (.B(net7515),
    .C(_11103_),
    .A(net7546),
    .Y(_11108_));
 sg13g2_mux2_1 _24721_ (.A0(net5840),
    .A1(_01507_),
    .S(_11076_),
    .X(_11109_));
 sg13g2_nand2_1 _24722_ (.Y(_11110_),
    .A(_01506_),
    .B(net6340));
 sg13g2_o21ai_1 _24723_ (.B1(_11110_),
    .Y(_11111_),
    .A1(net5834),
    .A2(_11076_));
 sg13g2_nand2_1 _24724_ (.Y(_11112_),
    .A(_01505_),
    .B(net6337));
 sg13g2_o21ai_1 _24725_ (.B1(_11112_),
    .Y(_11113_),
    .A1(net5900),
    .A2(net6100));
 sg13g2_nand2_1 _24726_ (.Y(_11114_),
    .A(_01504_),
    .B(net6337));
 sg13g2_o21ai_1 _24727_ (.B1(_11114_),
    .Y(_11115_),
    .A1(net5895),
    .A2(net6100));
 sg13g2_nand2_1 _24728_ (.Y(_11116_),
    .A(_01503_),
    .B(net6338));
 sg13g2_o21ai_1 _24729_ (.B1(_11116_),
    .Y(_11117_),
    .A1(net5891),
    .A2(net6338));
 sg13g2_mux2_1 _24730_ (.A0(net5775),
    .A1(_01502_),
    .S(_11074_),
    .X(_11118_));
 sg13g2_nand2_1 _24731_ (.Y(_11119_),
    .A(_01501_),
    .B(net6340));
 sg13g2_o21ai_1 _24732_ (.B1(_11119_),
    .Y(_11120_),
    .A1(net5886),
    .A2(net6338));
 sg13g2_nand2_1 _24733_ (.Y(_11121_),
    .A(_01500_),
    .B(net6357));
 sg13g2_o21ai_1 _24734_ (.B1(_11121_),
    .Y(_11122_),
    .A1(net5792),
    .A2(_10986_));
 sg13g2_nand2_1 _24735_ (.Y(_11123_),
    .A(_01499_),
    .B(net6345));
 sg13g2_o21ai_1 _24736_ (.B1(_11123_),
    .Y(_11124_),
    .A1(net5927),
    .A2(net6345));
 sg13g2_nand2_1 _24737_ (.Y(_11125_),
    .A(_01498_),
    .B(net6343));
 sg13g2_nand4_1 _24738_ (.B(_11002_),
    .C(_11022_),
    .A(_10957_),
    .Y(_11126_),
    .D(_11089_));
 sg13g2_o21ai_1 _24739_ (.B1(_11125_),
    .Y(_11127_),
    .A1(net5966),
    .A2(net6343));
 sg13g2_nand2_1 _24740_ (.Y(_11128_),
    .A(_01497_),
    .B(net6339));
 sg13g2_o21ai_1 _24741_ (.B1(_11128_),
    .Y(_11129_),
    .A1(net6012),
    .A2(net6339));
 sg13g2_nand2_1 _24742_ (.Y(_11130_),
    .A(_01496_),
    .B(net6340));
 sg13g2_o21ai_1 _24743_ (.B1(_11130_),
    .Y(_11131_),
    .A1(net5958),
    .A2(net6100));
 sg13g2_nand2_1 _24744_ (.Y(_11132_),
    .A(_01495_),
    .B(net6343));
 sg13g2_o21ai_1 _24745_ (.B1(_11132_),
    .Y(_11133_),
    .A1(net6009),
    .A2(net6343));
 sg13g2_nand2_1 _24746_ (.Y(_11134_),
    .A(_01494_),
    .B(net6339));
 sg13g2_o21ai_1 _24747_ (.B1(_11134_),
    .Y(_11135_),
    .A1(net6003),
    .A2(net6339));
 sg13g2_nand2_1 _24748_ (.Y(_11136_),
    .A(_01493_),
    .B(net6344));
 sg13g2_nand4_1 _24749_ (.B(_11045_),
    .C(_11064_),
    .A(_10974_),
    .Y(_11137_),
    .D(_11108_));
 sg13g2_o21ai_1 _24750_ (.B1(_11136_),
    .Y(_11138_),
    .A1(net6118),
    .A2(net6344));
 sg13g2_nand2_1 _24751_ (.Y(_11139_),
    .A(_01492_),
    .B(net6343));
 sg13g2_o21ai_1 _24752_ (.B1(_11139_),
    .Y(_11140_),
    .A1(net6031),
    .A2(net6343));
 sg13g2_nand2_1 _24753_ (.Y(_11141_),
    .A(_01491_),
    .B(net6344));
 sg13g2_o21ai_1 _24754_ (.B1(_11141_),
    .Y(_11142_),
    .A1(net6113),
    .A2(net6344));
 sg13g2_nand2_1 _24755_ (.Y(_11143_),
    .A(_01490_),
    .B(net6344));
 sg13g2_o21ai_1 _24756_ (.B1(_11143_),
    .Y(_11144_),
    .A1(net6027),
    .A2(net6344));
 sg13g2_nand2_1 _24757_ (.Y(_11145_),
    .A(_01489_),
    .B(net6362));
 sg13g2_nand2b_1 _24758_ (.Y(_11146_),
    .B(net6378),
    .A_N(net6362));
 sg13g2_nor4_1 _24759_ (.A(_10858_),
    .B(_10945_),
    .C(_11126_),
    .D(_11137_),
    .Y(_11147_));
 sg13g2_o21ai_1 _24760_ (.B1(_11145_),
    .Y(_11148_),
    .A1(net5921),
    .A2(_11146_));
 sg13g2_nand2_1 _24761_ (.Y(_11149_),
    .A(_01488_),
    .B(net6338));
 sg13g2_or4_1 _24762_ (.A(_10858_),
    .B(_10945_),
    .C(_11126_),
    .D(_11137_),
    .X(_11150_));
 sg13g2_o21ai_1 _24763_ (.B1(_11149_),
    .Y(_11151_),
    .A1(_09601_),
    .A2(net6338));
 sg13g2_nand2_1 _24764_ (.Y(_11152_),
    .A(_01487_),
    .B(net6339));
 sg13g2_o21ai_1 _24765_ (.B1(_11152_),
    .Y(_11153_),
    .A1(net6020),
    .A2(net6339));
 sg13g2_nand2_1 _24766_ (.Y(_11154_),
    .A(_01486_),
    .B(net6339));
 sg13g2_o21ai_1 _24767_ (.B1(_11154_),
    .Y(_11155_),
    .A1(net6106),
    .A2(net6339));
 sg13g2_nand2_1 _24768_ (.Y(_11156_),
    .A(_01485_),
    .B(net6337));
 sg13g2_o21ai_1 _24769_ (.B1(_11156_),
    .Y(_11157_),
    .A1(net5867),
    .A2(net6100));
 sg13g2_nor2b_1 _24770_ (.A(_01917_),
    .B_N(_01887_),
    .Y(_11158_));
 sg13g2_nand2b_1 _24771_ (.Y(_11159_),
    .B(net7932),
    .A_N(net7666));
 sg13g2_nand4_1 _24772_ (.B(net6466),
    .C(_09681_),
    .A(net7669),
    .Y(_11160_),
    .D(_11158_));
 sg13g2_nand2_1 _24773_ (.Y(_11161_),
    .A(_09683_),
    .B(net7447));
 sg13g2_nand2_1 _24774_ (.Y(_11162_),
    .A(_01484_),
    .B(net6327));
 sg13g2_o21ai_1 _24775_ (.B1(_11162_),
    .Y(_11163_),
    .A1(net5862),
    .A2(net6327));
 sg13g2_nand2b_1 _24776_ (.Y(_11164_),
    .B(net8000),
    .A_N(_01634_));
 sg13g2_nand2_1 _24777_ (.Y(_11165_),
    .A(_01483_),
    .B(net6330));
 sg13g2_nand2b_1 _24778_ (.Y(_11166_),
    .B(net6383),
    .A_N(net6330));
 sg13g2_o21ai_1 _24779_ (.B1(_11165_),
    .Y(_11167_),
    .A1(net5857),
    .A2(_11166_));
 sg13g2_nand2_1 _24780_ (.Y(_11168_),
    .A(_01482_),
    .B(net6331));
 sg13g2_o21ai_1 _24781_ (.B1(_11164_),
    .Y(_11169_),
    .A1(_01629_),
    .A2(net7479));
 sg13g2_o21ai_1 _24782_ (.B1(_11168_),
    .Y(_11170_),
    .A1(net5808),
    .A2(_11161_));
 sg13g2_nand2_1 _24783_ (.Y(_11171_),
    .A(_01481_),
    .B(net6329));
 sg13g2_a21oi_1 _24784_ (.A1(net8006),
    .A2(net7283),
    .Y(_11172_),
    .B1(_11169_));
 sg13g2_o21ai_1 _24785_ (.B1(_11171_),
    .Y(_11173_),
    .A1(net5850),
    .A2(net6329));
 sg13g2_nand2_1 _24786_ (.Y(_11174_),
    .A(_01480_),
    .B(net6328));
 sg13g2_o21ai_1 _24787_ (.B1(_11174_),
    .Y(_11175_),
    .A1(net5800),
    .A2(net6328));
 sg13g2_nand2_1 _24788_ (.Y(_11176_),
    .A(_01479_),
    .B(net6331));
 sg13g2_o21ai_1 _24789_ (.B1(_11176_),
    .Y(_11177_),
    .A1(net5795),
    .A2(net5999));
 sg13g2_nand2_1 _24790_ (.Y(_11178_),
    .A(_01478_),
    .B(net6356));
 sg13g2_o21ai_1 _24791_ (.B1(_11178_),
    .Y(_11179_),
    .A1(net5786),
    .A2(_10986_));
 sg13g2_o21ai_1 _24792_ (.B1(_11172_),
    .Y(_11180_),
    .A1(_09277_),
    .A2(_10750_));
 sg13g2_nand2_1 _24793_ (.Y(_11181_),
    .A(_01477_),
    .B(net6330));
 sg13g2_nand2b_1 _24794_ (.Y(_11182_),
    .B(net6379),
    .A_N(net6330));
 sg13g2_o21ai_1 _24795_ (.B1(_11181_),
    .Y(_11183_),
    .A1(net5918),
    .A2(_11182_));
 sg13g2_nand2_1 _24796_ (.Y(_11184_),
    .A(_01476_),
    .B(net6331));
 sg13g2_o21ai_1 _24797_ (.B1(_11184_),
    .Y(_11185_),
    .A1(net5789),
    .A2(net5999));
 sg13g2_nand2_1 _24798_ (.Y(_11186_),
    .A(_01475_),
    .B(net6327));
 sg13g2_nand2b_1 _24799_ (.Y(_11187_),
    .B(net6374),
    .A_N(net6327));
 sg13g2_o21ai_1 _24800_ (.B1(_11186_),
    .Y(_11188_),
    .A1(net5912),
    .A2(_11187_));
 sg13g2_nand2_1 _24801_ (.Y(_11189_),
    .A(_01474_),
    .B(net6331));
 sg13g2_o21ai_1 _24802_ (.B1(_11189_),
    .Y(_11190_),
    .A1(net5778),
    .A2(_11161_));
 sg13g2_nand2_1 _24803_ (.Y(_11191_),
    .A(_01473_),
    .B(net6327));
 sg13g2_nand2b_1 _24804_ (.Y(_11192_),
    .B(net6366),
    .A_N(net6327));
 sg13g2_o21ai_1 _24805_ (.B1(_11191_),
    .Y(_11193_),
    .A1(net5910),
    .A2(_11192_));
 sg13g2_a22oi_1 _24806_ (.Y(_11194_),
    .B1(_11180_),
    .B2(net7377),
    .A2(_10788_),
    .A1(net6917));
 sg13g2_mux2_1 _24807_ (.A0(net5840),
    .A1(_01472_),
    .S(_11161_),
    .X(_11195_));
 sg13g2_nand2_1 _24808_ (.Y(_11196_),
    .A(_01471_),
    .B(net6334));
 sg13g2_o21ai_1 _24809_ (.B1(_11196_),
    .Y(_11197_),
    .A1(net5833),
    .A2(net5999));
 sg13g2_nand2_1 _24810_ (.Y(_11198_),
    .A(_01470_),
    .B(net6331));
 sg13g2_o21ai_1 _24811_ (.B1(_11198_),
    .Y(_11199_),
    .A1(net5900),
    .A2(net5999));
 sg13g2_nand2_1 _24812_ (.Y(_11200_),
    .A(_01469_),
    .B(net6331));
 sg13g2_o21ai_1 _24813_ (.B1(_11200_),
    .Y(_11201_),
    .A1(net5899),
    .A2(_11161_));
 sg13g2_nand2_1 _24814_ (.Y(_11202_),
    .A(_01468_),
    .B(net6334));
 sg13g2_o21ai_1 _24815_ (.B1(_11202_),
    .Y(_11203_),
    .A1(net5892),
    .A2(net6332));
 sg13g2_nand2_1 _24816_ (.Y(_11204_),
    .A(_01467_),
    .B(net6357));
 sg13g2_o21ai_1 _24817_ (.B1(_11194_),
    .Y(_11205_),
    .A1(net6981),
    .A2(_10788_));
 sg13g2_nand2b_1 _24818_ (.Y(_11206_),
    .B(net6369),
    .A_N(net6357));
 sg13g2_o21ai_1 _24819_ (.B1(_11204_),
    .Y(_11207_),
    .A1(net5915),
    .A2(_11206_));
 sg13g2_mux2_1 _24820_ (.A0(net5775),
    .A1(_01466_),
    .S(net6327),
    .X(_11208_));
 sg13g2_nand2_1 _24821_ (.Y(_11209_),
    .A(_01465_),
    .B(net6332));
 sg13g2_o21ai_1 _24822_ (.B1(_11209_),
    .Y(_11210_),
    .A1(net5882),
    .A2(net6332));
 sg13g2_nand2_1 _24823_ (.Y(_11211_),
    .A(_01464_),
    .B(net6328));
 sg13g2_o21ai_1 _24824_ (.B1(_11211_),
    .Y(_11212_),
    .A1(net5928),
    .A2(net6328));
 sg13g2_nand2_1 _24825_ (.Y(_11213_),
    .A(_01463_),
    .B(net6328));
 sg13g2_o21ai_1 _24826_ (.B1(_11213_),
    .Y(_11214_),
    .A1(net5966),
    .A2(net6328));
 sg13g2_nand2_1 _24827_ (.Y(_11215_),
    .A(_01462_),
    .B(net6333));
 sg13g2_o21ai_1 _24828_ (.B1(_11215_),
    .Y(_11216_),
    .A1(_10857_),
    .A2(net6333));
 sg13g2_nand2_1 _24829_ (.Y(_11217_),
    .A(_01461_),
    .B(net6331));
 sg13g2_o21ai_1 _24830_ (.B1(_11217_),
    .Y(_11218_),
    .A1(net5958),
    .A2(_11161_));
 sg13g2_nand2_1 _24831_ (.Y(_11219_),
    .A(_01460_),
    .B(net6333));
 sg13g2_o21ai_1 _24832_ (.B1(_11219_),
    .Y(_11220_),
    .A1(net6009),
    .A2(net6333));
 sg13g2_nand2_1 _24833_ (.Y(_11221_),
    .A(_01459_),
    .B(net6332));
 sg13g2_o21ai_1 _24834_ (.B1(_11221_),
    .Y(_11222_),
    .A1(net6003),
    .A2(net6334));
 sg13g2_a22oi_1 _24835_ (.Y(_11223_),
    .B1(_09397_),
    .B2(_01887_),
    .A2(_08800_),
    .A1(net7692));
 sg13g2_nand2_1 _24836_ (.Y(_11224_),
    .A(_01458_),
    .B(net6329));
 sg13g2_o21ai_1 _24837_ (.B1(_11224_),
    .Y(_11225_),
    .A1(net6119),
    .A2(net6329));
 sg13g2_nand2_1 _24838_ (.Y(_11226_),
    .A(_01457_),
    .B(net6333));
 sg13g2_o21ai_1 _24839_ (.B1(_11226_),
    .Y(_11227_),
    .A1(net6030),
    .A2(net6333));
 sg13g2_nand2_1 _24840_ (.Y(_11228_),
    .A(_01456_),
    .B(net6363));
 sg13g2_o21ai_1 _24841_ (.B1(_11228_),
    .Y(_11229_),
    .A1(net5783),
    .A2(net6000));
 sg13g2_nand2_1 _24842_ (.Y(_11230_),
    .A(_01455_),
    .B(net6329));
 sg13g2_o21ai_1 _24843_ (.B1(_11230_),
    .Y(_11231_),
    .A1(net6113),
    .A2(net6329));
 sg13g2_nand2_1 _24844_ (.Y(_11232_),
    .A(_01454_),
    .B(net6329));
 sg13g2_o21ai_1 _24845_ (.B1(_11232_),
    .Y(_11233_),
    .A1(net6024),
    .A2(net6329));
 sg13g2_nand2_1 _24846_ (.Y(_11234_),
    .A(_01453_),
    .B(net6332));
 sg13g2_o21ai_1 _24847_ (.B1(_11234_),
    .Y(_11235_),
    .A1(net6053),
    .A2(net6332));
 sg13g2_nand2_1 _24848_ (.Y(_11236_),
    .A(_01452_),
    .B(net6332));
 sg13g2_o21ai_1 _24849_ (.B1(_11236_),
    .Y(_11237_),
    .A1(net6020),
    .A2(net6332));
 sg13g2_nand2_1 _24850_ (.Y(_11238_),
    .A(_01451_),
    .B(net6333));
 sg13g2_o21ai_1 _24851_ (.B1(_11238_),
    .Y(_11239_),
    .A1(net6104),
    .A2(net6333));
 sg13g2_nand2_1 _24852_ (.Y(_11240_),
    .A(_01450_),
    .B(net6331));
 sg13g2_o21ai_1 _24853_ (.B1(_11240_),
    .Y(_11241_),
    .A1(net5867),
    .A2(_11161_));
 sg13g2_nand4_1 _24854_ (.B(net6466),
    .C(_10091_),
    .A(net7669),
    .Y(_11242_),
    .D(_11158_));
 sg13g2_nand2_1 _24855_ (.Y(_11243_),
    .A(_10094_),
    .B(net7447));
 sg13g2_nand2_1 _24856_ (.Y(_11244_),
    .A(_01449_),
    .B(net6322));
 sg13g2_o21ai_1 _24857_ (.B1(_11244_),
    .Y(_11245_),
    .A1(net5862),
    .A2(net6322));
 sg13g2_nand2_1 _24858_ (.Y(_11246_),
    .A(_01448_),
    .B(net6321));
 sg13g2_nand2b_1 _24859_ (.Y(_11247_),
    .B(net6383),
    .A_N(net6321));
 sg13g2_o21ai_1 _24860_ (.B1(_11246_),
    .Y(_11248_),
    .A1(net5857),
    .A2(_11247_));
 sg13g2_nand2_1 _24861_ (.Y(_11249_),
    .A(_01447_),
    .B(net6323));
 sg13g2_o21ai_1 _24862_ (.B1(_11249_),
    .Y(_11250_),
    .A1(net5808),
    .A2(_11243_));
 sg13g2_nand2_1 _24863_ (.Y(_11251_),
    .A(_01446_),
    .B(net6320));
 sg13g2_o21ai_1 _24864_ (.B1(_11251_),
    .Y(_11252_),
    .A1(net5850),
    .A2(net6320));
 sg13g2_nand2b_1 _24865_ (.Y(_11253_),
    .B(net6364),
    .A_N(net6357));
 sg13g2_nand2_1 _24866_ (.Y(_11254_),
    .A(_01445_),
    .B(net6357));
 sg13g2_o21ai_1 _24867_ (.B1(_11254_),
    .Y(_11255_),
    .A1(net5907),
    .A2(_11253_));
 sg13g2_nand2_1 _24868_ (.Y(_11256_),
    .A(_01444_),
    .B(net6319));
 sg13g2_o21ai_1 _24869_ (.B1(_11256_),
    .Y(_11257_),
    .A1(net5802),
    .A2(net6319));
 sg13g2_nand2_1 _24870_ (.Y(_11258_),
    .A(_01443_),
    .B(net6323));
 sg13g2_o21ai_1 _24871_ (.B1(_11258_),
    .Y(_11259_),
    .A1(net5795),
    .A2(net5998));
 sg13g2_nand2_1 _24872_ (.Y(_11260_),
    .A(_01442_),
    .B(net6321));
 sg13g2_nand2b_1 _24873_ (.Y(_11261_),
    .B(net6379),
    .A_N(net6321));
 sg13g2_o21ai_1 _24874_ (.B1(_11260_),
    .Y(_11262_),
    .A1(net5918),
    .A2(_11261_));
 sg13g2_nand2_1 _24875_ (.Y(_11263_),
    .A(_01441_),
    .B(net6323));
 sg13g2_o21ai_1 _24876_ (.B1(_11263_),
    .Y(_11264_),
    .A1(net5789),
    .A2(net5998));
 sg13g2_nand2_1 _24877_ (.Y(_11265_),
    .A(_01440_),
    .B(net6322));
 sg13g2_nand2b_1 _24878_ (.Y(_11266_),
    .B(net6374),
    .A_N(net6322));
 sg13g2_o21ai_1 _24879_ (.B1(_11265_),
    .Y(_11267_),
    .A1(net5912),
    .A2(_11266_));
 sg13g2_nand2_1 _24880_ (.Y(_11268_),
    .A(_01439_),
    .B(net6323));
 sg13g2_o21ai_1 _24881_ (.B1(_11268_),
    .Y(_11269_),
    .A1(net5778),
    .A2(_11243_));
 sg13g2_nand2_1 _24882_ (.Y(_11270_),
    .A(_01438_),
    .B(_11242_));
 sg13g2_nand2b_1 _24883_ (.Y(_11271_),
    .B(net6366),
    .A_N(net6321));
 sg13g2_mux4_1 _24884_ (.S0(net7765),
    .A0(_00791_),
    .A1(_00823_),
    .A2(_00855_),
    .A3(_00890_),
    .S1(net7725),
    .X(_11272_));
 sg13g2_o21ai_1 _24885_ (.B1(_11270_),
    .Y(_11273_),
    .A1(net5910),
    .A2(_11271_));
 sg13g2_nand2_1 _24886_ (.Y(_11274_),
    .A(net7605),
    .B(_11272_));
 sg13g2_mux2_1 _24887_ (.A0(net5840),
    .A1(_01437_),
    .S(_11243_),
    .X(_11275_));
 sg13g2_nand2_1 _24888_ (.Y(_11276_),
    .A(_01436_),
    .B(net6326));
 sg13g2_o21ai_1 _24889_ (.B1(_11276_),
    .Y(_11277_),
    .A1(net5833),
    .A2(net5998));
 sg13g2_nand2_1 _24890_ (.Y(_11278_),
    .A(_01435_),
    .B(net6323));
 sg13g2_o21ai_1 _24891_ (.B1(_11278_),
    .Y(_11279_),
    .A1(net5900),
    .A2(net5998));
 sg13g2_mux2_1 _24892_ (.A0(net5838),
    .A1(_01434_),
    .S(net6000),
    .X(_11280_));
 sg13g2_nand2_1 _24893_ (.Y(_11281_),
    .A(_01433_),
    .B(net6323));
 sg13g2_a21oi_1 _24894_ (.A1(_00895_),
    .A2(net7423),
    .Y(_11282_),
    .B1(net7687));
 sg13g2_o21ai_1 _24895_ (.B1(_11281_),
    .Y(_11283_),
    .A1(net5895),
    .A2(_11243_));
 sg13g2_nand2_1 _24896_ (.Y(_11284_),
    .A(_01432_),
    .B(net6326));
 sg13g2_o21ai_1 _24897_ (.B1(_11284_),
    .Y(_11285_),
    .A1(net5892),
    .A2(net6326));
 sg13g2_mux2_1 _24898_ (.A0(net5775),
    .A1(_01431_),
    .S(net6322),
    .X(_11286_));
 sg13g2_nand2_1 _24899_ (.Y(_11287_),
    .A(_01430_),
    .B(net6324));
 sg13g2_o21ai_1 _24900_ (.B1(_11287_),
    .Y(_11288_),
    .A1(net5882),
    .A2(net6324));
 sg13g2_nand2_1 _24901_ (.Y(_11289_),
    .A(_01429_),
    .B(net6319));
 sg13g2_o21ai_1 _24902_ (.B1(_11289_),
    .Y(_11290_),
    .A1(net5929),
    .A2(net6319));
 sg13g2_nand2_1 _24903_ (.Y(_11291_),
    .A(_01428_),
    .B(net6319));
 sg13g2_o21ai_1 _24904_ (.B1(_11291_),
    .Y(_11292_),
    .A1(net5966),
    .A2(net6319));
 sg13g2_mux2_1 _24905_ (.A0(_01599_),
    .A1(_00759_),
    .S(net7703),
    .X(_11293_));
 sg13g2_nand2_1 _24906_ (.Y(_11294_),
    .A(_01427_),
    .B(net6325));
 sg13g2_o21ai_1 _24907_ (.B1(_11294_),
    .Y(_11295_),
    .A1(net6013),
    .A2(net6325));
 sg13g2_nand2_1 _24908_ (.Y(_11296_),
    .A(_01426_),
    .B(net6323));
 sg13g2_o21ai_1 _24909_ (.B1(_11296_),
    .Y(_11297_),
    .A1(net5958),
    .A2(_11243_));
 sg13g2_nand2_1 _24910_ (.Y(_11298_),
    .A(_01425_),
    .B(net6325));
 sg13g2_o21ai_1 _24911_ (.B1(_11298_),
    .Y(_11299_),
    .A1(net6009),
    .A2(net6325));
 sg13g2_nand2_1 _24912_ (.Y(_11300_),
    .A(_01424_),
    .B(net6324));
 sg13g2_o21ai_1 _24913_ (.B1(_11300_),
    .Y(_11301_),
    .A1(net6007),
    .A2(net6324));
 sg13g2_nand2_1 _24914_ (.Y(_11302_),
    .A(_01423_),
    .B(net6356));
 sg13g2_o21ai_1 _24915_ (.B1(_11302_),
    .Y(_11303_),
    .A1(net5836),
    .A2(_10986_));
 sg13g2_nand2_1 _24916_ (.Y(_11304_),
    .A(_01422_),
    .B(net6320));
 sg13g2_a22oi_1 _24917_ (.Y(_11305_),
    .B1(_11293_),
    .B2(net7435),
    .A2(net7424),
    .A1(_01247_));
 sg13g2_o21ai_1 _24918_ (.B1(_11304_),
    .Y(_11306_),
    .A1(net6119),
    .A2(net6320));
 sg13g2_nand2_1 _24919_ (.Y(_11307_),
    .A(_01421_),
    .B(net6325));
 sg13g2_o21ai_1 _24920_ (.B1(_11307_),
    .Y(_11308_),
    .A1(net6030),
    .A2(net6325));
 sg13g2_nand2_1 _24921_ (.Y(_11309_),
    .A(_01420_),
    .B(net6320));
 sg13g2_o21ai_1 _24922_ (.B1(_11309_),
    .Y(_11310_),
    .A1(net6113),
    .A2(net6320));
 sg13g2_nand2_1 _24923_ (.Y(_11311_),
    .A(_01419_),
    .B(net6320));
 sg13g2_o21ai_1 _24924_ (.B1(_11311_),
    .Y(_11312_),
    .A1(net6024),
    .A2(net6320));
 sg13g2_nand2_1 _24925_ (.Y(_11313_),
    .A(_01418_),
    .B(net6326));
 sg13g2_o21ai_1 _24926_ (.B1(_11313_),
    .Y(_11314_),
    .A1(net6053),
    .A2(net6326));
 sg13g2_nand2_1 _24927_ (.Y(_11315_),
    .A(_01417_),
    .B(net6325));
 sg13g2_o21ai_1 _24928_ (.B1(_11315_),
    .Y(_11316_),
    .A1(net6021),
    .A2(net6325));
 sg13g2_nand2_1 _24929_ (.Y(_11317_),
    .A(_01416_),
    .B(net6324));
 sg13g2_o21ai_1 _24930_ (.B1(_11317_),
    .Y(_11318_),
    .A1(net6104),
    .A2(net6324));
 sg13g2_nand2_1 _24931_ (.Y(_11319_),
    .A(_01415_),
    .B(net6323));
 sg13g2_o21ai_1 _24932_ (.B1(_11319_),
    .Y(_11320_),
    .A1(net5867),
    .A2(_11243_));
 sg13g2_or4_1 _24933_ (.A(net7671),
    .B(net6467),
    .C(_09682_),
    .D(_11159_),
    .X(_11321_));
 sg13g2_nand2_1 _24934_ (.Y(_11322_),
    .A(net6346),
    .B(net7447));
 sg13g2_nand2_1 _24935_ (.Y(_11323_),
    .A(_01414_),
    .B(net6316));
 sg13g2_o21ai_1 _24936_ (.B1(_11323_),
    .Y(_11324_),
    .A1(net8286),
    .A2(net6316));
 sg13g2_nand2_1 _24937_ (.Y(_11325_),
    .A(_01413_),
    .B(net6318));
 sg13g2_nand2b_1 _24938_ (.Y(_11326_),
    .B(net6383),
    .A_N(_11321_));
 sg13g2_o21ai_1 _24939_ (.B1(_11325_),
    .Y(_11327_),
    .A1(net5857),
    .A2(_11326_));
 sg13g2_nand2_1 _24940_ (.Y(_11328_),
    .A(_01412_),
    .B(net6363));
 sg13g2_o21ai_1 _24941_ (.B1(_11328_),
    .Y(_11329_),
    .A1(net5902),
    .A2(net6000));
 sg13g2_nand2_1 _24942_ (.Y(_11330_),
    .A(_01411_),
    .B(net6314));
 sg13g2_o21ai_1 _24943_ (.B1(_11330_),
    .Y(_11331_),
    .A1(net5808),
    .A2(net6099));
 sg13g2_nand2_1 _24944_ (.Y(_11332_),
    .A(_01410_),
    .B(net6317));
 sg13g2_o21ai_1 _24945_ (.B1(_11332_),
    .Y(_11333_),
    .A1(net5849),
    .A2(net6317));
 sg13g2_nand2_1 _24946_ (.Y(_11334_),
    .A(_01409_),
    .B(net6318));
 sg13g2_o21ai_1 _24947_ (.B1(_11334_),
    .Y(_11335_),
    .A1(net5802),
    .A2(net6318));
 sg13g2_nand2_1 _24948_ (.Y(_11336_),
    .A(_01408_),
    .B(net6314));
 sg13g2_o21ai_1 _24949_ (.B1(_11336_),
    .Y(_11337_),
    .A1(net5795),
    .A2(net6099));
 sg13g2_nand2_1 _24950_ (.Y(_11338_),
    .A(_01407_),
    .B(_11321_));
 sg13g2_nand2b_1 _24951_ (.Y(_11339_),
    .B(net6379),
    .A_N(_11321_));
 sg13g2_o21ai_1 _24952_ (.B1(_11338_),
    .Y(_11340_),
    .A1(net5917),
    .A2(_11339_));
 sg13g2_nand2_1 _24953_ (.Y(_11341_),
    .A(_01406_),
    .B(net6314));
 sg13g2_o21ai_1 _24954_ (.B1(_11341_),
    .Y(_11342_),
    .A1(net5789),
    .A2(net6099));
 sg13g2_nand2_1 _24955_ (.Y(_11343_),
    .A(_01405_),
    .B(net6316));
 sg13g2_nand2b_1 _24956_ (.Y(_11344_),
    .B(net6374),
    .A_N(net6316));
 sg13g2_o21ai_1 _24957_ (.B1(_11343_),
    .Y(_11345_),
    .A1(net5912),
    .A2(_11344_));
 sg13g2_nand2_1 _24958_ (.Y(_11346_),
    .A(_01404_),
    .B(net6314));
 sg13g2_o21ai_1 _24959_ (.B1(_11346_),
    .Y(_11347_),
    .A1(net5778),
    .A2(net6099));
 sg13g2_nand2_1 _24960_ (.Y(_11348_),
    .A(_01403_),
    .B(net6316));
 sg13g2_nand2b_1 _24961_ (.Y(_11349_),
    .B(net6366),
    .A_N(net6316));
 sg13g2_o21ai_1 _24962_ (.B1(_11348_),
    .Y(_11350_),
    .A1(net5910),
    .A2(_11349_));
 sg13g2_mux2_1 _24963_ (.A0(net5840),
    .A1(_01402_),
    .S(_11322_),
    .X(_11351_));
 sg13g2_nand2_1 _24964_ (.Y(_11352_),
    .A(_01401_),
    .B(net6363));
 sg13g2_mux4_1 _24965_ (.S0(net7770),
    .A0(_00925_),
    .A1(_00960_),
    .A2(_00996_),
    .A3(_01031_),
    .S1(net7723),
    .X(_11353_));
 sg13g2_o21ai_1 _24966_ (.B1(_11352_),
    .Y(_11354_),
    .A1(net5897),
    .A2(_10986_));
 sg13g2_nand2_1 _24967_ (.Y(_11355_),
    .A(_01400_),
    .B(net6311));
 sg13g2_o21ai_1 _24968_ (.B1(_11355_),
    .Y(_11356_),
    .A1(net5833),
    .A2(net6099));
 sg13g2_nand2_1 _24969_ (.Y(_11357_),
    .A(_01399_),
    .B(net6314));
 sg13g2_o21ai_1 _24970_ (.B1(_11357_),
    .Y(_11358_),
    .A1(net5900),
    .A2(net6099));
 sg13g2_nand2_1 _24971_ (.Y(_11359_),
    .A(_01398_),
    .B(net6314));
 sg13g2_o21ai_1 _24972_ (.B1(_11359_),
    .Y(_11360_),
    .A1(net5895),
    .A2(net6099));
 sg13g2_nand2_1 _24973_ (.Y(_11361_),
    .A(_01397_),
    .B(net6311));
 sg13g2_o21ai_1 _24974_ (.B1(_11361_),
    .Y(_11362_),
    .A1(net5891),
    .A2(net6311));
 sg13g2_mux2_1 _24975_ (.A0(net5775),
    .A1(_01396_),
    .S(net6316),
    .X(_11363_));
 sg13g2_nand2_1 _24976_ (.Y(_11364_),
    .A(_01395_),
    .B(net6312));
 sg13g2_o21ai_1 _24977_ (.B1(_11364_),
    .Y(_11365_),
    .A1(net5882),
    .A2(net6312));
 sg13g2_nand2_1 _24978_ (.Y(_11366_),
    .A(_01394_),
    .B(net6318));
 sg13g2_mux2_1 _24979_ (.A0(_00663_),
    .A1(_00695_),
    .S(net7779),
    .X(_11367_));
 sg13g2_o21ai_1 _24980_ (.B1(_11366_),
    .Y(_11368_),
    .A1(net5928),
    .A2(net6318));
 sg13g2_nand2_1 _24981_ (.Y(_11369_),
    .A(_01393_),
    .B(net6318));
 sg13g2_o21ai_1 _24982_ (.B1(_11369_),
    .Y(_11370_),
    .A1(net5966),
    .A2(net6318));
 sg13g2_nand2_1 _24983_ (.Y(_11371_),
    .A(_01392_),
    .B(net6313));
 sg13g2_o21ai_1 _24984_ (.B1(_11371_),
    .Y(_11372_),
    .A1(net6013),
    .A2(net6313));
 sg13g2_nand2_1 _24985_ (.Y(_11373_),
    .A(_01391_),
    .B(net6314));
 sg13g2_o21ai_1 _24986_ (.B1(_11373_),
    .Y(_11374_),
    .A1(net5958),
    .A2(_11322_));
 sg13g2_nand2_1 _24987_ (.Y(_11375_),
    .A(_01390_),
    .B(net6356));
 sg13g2_o21ai_1 _24988_ (.B1(_11375_),
    .Y(_11376_),
    .A1(net5888),
    .A2(net6356));
 sg13g2_nand2_1 _24989_ (.Y(_11377_),
    .A(_01389_),
    .B(net6313));
 sg13g2_o21ai_1 _24990_ (.B1(_11377_),
    .Y(_11378_),
    .A1(net6009),
    .A2(net6313));
 sg13g2_nand2_1 _24991_ (.Y(_11379_),
    .A(_01388_),
    .B(net6312));
 sg13g2_o21ai_1 _24992_ (.B1(_11379_),
    .Y(_11380_),
    .A1(net6004),
    .A2(net6315));
 sg13g2_nand2_1 _24993_ (.Y(_11381_),
    .A(_01387_),
    .B(net6317));
 sg13g2_o21ai_1 _24994_ (.B1(_11381_),
    .Y(_11382_),
    .A1(_09678_),
    .A2(net6317));
 sg13g2_nand2_1 _24995_ (.Y(_11383_),
    .A(_01386_),
    .B(net6313));
 sg13g2_o21ai_1 _24996_ (.B1(_11383_),
    .Y(_11384_),
    .A1(net6030),
    .A2(net6313));
 sg13g2_nand2_1 _24997_ (.Y(_11385_),
    .A(_01385_),
    .B(net6317));
 sg13g2_o21ai_1 _24998_ (.B1(_11385_),
    .Y(_11386_),
    .A1(net6113),
    .A2(net6317));
 sg13g2_nand2_1 _24999_ (.Y(_11387_),
    .A(_01384_),
    .B(net6317));
 sg13g2_o21ai_1 _25000_ (.B1(_11387_),
    .Y(_11388_),
    .A1(net6028),
    .A2(net6317));
 sg13g2_nand2_1 _25001_ (.Y(_11389_),
    .A(_01383_),
    .B(net6311));
 sg13g2_o21ai_1 _25002_ (.B1(_11389_),
    .Y(_11390_),
    .A1(net6053),
    .A2(net6311));
 sg13g2_nand2_1 _25003_ (.Y(_11391_),
    .A(_01382_),
    .B(net6312));
 sg13g2_o21ai_1 _25004_ (.B1(_11391_),
    .Y(_11392_),
    .A1(net6020),
    .A2(net6312));
 sg13g2_nand2_1 _25005_ (.Y(_11393_),
    .A(_01381_),
    .B(net6313));
 sg13g2_o21ai_1 _25006_ (.B1(_11393_),
    .Y(_11394_),
    .A1(net6104),
    .A2(net6313));
 sg13g2_nand2_1 _25007_ (.Y(_11395_),
    .A(_01380_),
    .B(net6314));
 sg13g2_o21ai_1 _25008_ (.B1(_11395_),
    .Y(_11396_),
    .A1(net5867),
    .A2(net6099));
 sg13g2_mux2_1 _25009_ (.A0(net5773),
    .A1(_01379_),
    .S(net6357),
    .X(_11397_));
 sg13g2_or4_1 _25010_ (.A(net7671),
    .B(net6467),
    .C(_10092_),
    .D(_11159_),
    .X(_11398_));
 sg13g2_nand2_1 _25011_ (.Y(_11399_),
    .A(net6335),
    .B(net7447));
 sg13g2_nand2_1 _25012_ (.Y(_11400_),
    .A(_01378_),
    .B(net6308));
 sg13g2_a22oi_1 _25013_ (.Y(_11401_),
    .B1(_11367_),
    .B2(net7519),
    .A2(net7594),
    .A1(_00727_));
 sg13g2_o21ai_1 _25014_ (.B1(_11400_),
    .Y(_11402_),
    .A1(net8286),
    .A2(net6308));
 sg13g2_nand2_1 _25015_ (.Y(_11403_),
    .A(_01377_),
    .B(_11398_));
 sg13g2_nand2b_1 _25016_ (.Y(_11404_),
    .B(net6383),
    .A_N(_11398_));
 sg13g2_o21ai_1 _25017_ (.B1(_11403_),
    .Y(_11405_),
    .A1(net5857),
    .A2(_11404_));
 sg13g2_nand2_1 _25018_ (.Y(_11406_),
    .A(_01376_),
    .B(net6304));
 sg13g2_o21ai_1 _25019_ (.B1(_11406_),
    .Y(_11407_),
    .A1(net5808),
    .A2(net6098));
 sg13g2_nand2_1 _25020_ (.Y(_11408_),
    .A(_01375_),
    .B(net6309));
 sg13g2_o21ai_1 _25021_ (.B1(_11408_),
    .Y(_11409_),
    .A1(net5851),
    .A2(net6309));
 sg13g2_nand2_1 _25022_ (.Y(_11410_),
    .A(_01374_),
    .B(net6310));
 sg13g2_o21ai_1 _25023_ (.B1(_11410_),
    .Y(_11411_),
    .A1(net5802),
    .A2(net6310));
 sg13g2_nand2_1 _25024_ (.Y(_11412_),
    .A(_01373_),
    .B(net6304));
 sg13g2_o21ai_1 _25025_ (.B1(_11412_),
    .Y(_11413_),
    .A1(net5795),
    .A2(_11399_));
 sg13g2_nand2b_1 _25026_ (.Y(_11414_),
    .B(net6379),
    .A_N(_11398_));
 sg13g2_nand2_1 _25027_ (.Y(_11415_),
    .A(_01372_),
    .B(_11398_));
 sg13g2_o21ai_1 _25028_ (.B1(net7703),
    .Y(_11416_),
    .A1(net7532),
    .A2(_11353_));
 sg13g2_o21ai_1 _25029_ (.B1(_11415_),
    .Y(_11417_),
    .A1(net5918),
    .A2(_11414_));
 sg13g2_nand2_1 _25030_ (.Y(_11418_),
    .A(_01371_),
    .B(net6304));
 sg13g2_o21ai_1 _25031_ (.B1(_11418_),
    .Y(_11419_),
    .A1(net5789),
    .A2(_11399_));
 sg13g2_nand2b_1 _25032_ (.Y(_11420_),
    .B(net6374),
    .A_N(net6308));
 sg13g2_nand2_1 _25033_ (.Y(_11421_),
    .A(_01370_),
    .B(net6308));
 sg13g2_o21ai_1 _25034_ (.B1(_11421_),
    .Y(_11422_),
    .A1(net5912),
    .A2(_11420_));
 sg13g2_nand2_1 _25035_ (.Y(_11423_),
    .A(_01369_),
    .B(net6304));
 sg13g2_o21ai_1 _25036_ (.B1(_11423_),
    .Y(_11424_),
    .A1(net5778),
    .A2(net6098));
 sg13g2_nand2_1 _25037_ (.Y(_11425_),
    .A(_01368_),
    .B(net6356));
 sg13g2_o21ai_1 _25038_ (.B1(_11425_),
    .Y(_11426_),
    .A1(net5885),
    .A2(net6356));
 sg13g2_nand2b_1 _25039_ (.Y(_11427_),
    .B(net6366),
    .A_N(net6308));
 sg13g2_nand2_1 _25040_ (.Y(_11428_),
    .A(_01367_),
    .B(net6308));
 sg13g2_a21o_1 _25041_ (.A2(_11401_),
    .A1(net7532),
    .B1(_11416_),
    .X(_11429_));
 sg13g2_o21ai_1 _25042_ (.B1(_11428_),
    .Y(_11430_),
    .A1(net5910),
    .A2(_11427_));
 sg13g2_mux2_1 _25043_ (.A0(net5840),
    .A1(_01366_),
    .S(_11399_),
    .X(_11431_));
 sg13g2_nand4_1 _25044_ (.B(_11282_),
    .C(_11305_),
    .A(_11274_),
    .Y(_11432_),
    .D(_11429_));
 sg13g2_nand2_1 _25045_ (.Y(_11433_),
    .A(_01365_),
    .B(net6307));
 sg13g2_o21ai_1 _25046_ (.B1(_11433_),
    .Y(_11434_),
    .A1(net5833),
    .A2(_11399_));
 sg13g2_nand2_1 _25047_ (.Y(_11435_),
    .A(_01364_),
    .B(net6304));
 sg13g2_o21ai_1 _25048_ (.B1(_11435_),
    .Y(_11436_),
    .A1(net5904),
    .A2(net6098));
 sg13g2_nand2_1 _25049_ (.Y(_11437_),
    .A(_01363_),
    .B(net6304));
 sg13g2_o21ai_1 _25050_ (.B1(_11437_),
    .Y(_11438_),
    .A1(net5895),
    .A2(net6098));
 sg13g2_nand2_1 _25051_ (.Y(_11439_),
    .A(_01362_),
    .B(net6307));
 sg13g2_o21ai_1 _25052_ (.B1(_11439_),
    .Y(_11440_),
    .A1(net5891),
    .A2(net6307));
 sg13g2_mux2_1 _25053_ (.A0(net5775),
    .A1(_01361_),
    .S(net6308),
    .X(_11441_));
 sg13g2_nand2_1 _25054_ (.Y(_11442_),
    .A(_01360_),
    .B(net6305));
 sg13g2_o21ai_1 _25055_ (.B1(_11442_),
    .Y(_11443_),
    .A1(net5882),
    .A2(net6305));
 sg13g2_nand2_1 _25056_ (.Y(_11444_),
    .A(_01359_),
    .B(net6310));
 sg13g2_o21ai_1 _25057_ (.B1(_11444_),
    .Y(_11445_),
    .A1(net5928),
    .A2(net6310));
 sg13g2_nand2_1 _25058_ (.Y(_11446_),
    .A(_01358_),
    .B(net6310));
 sg13g2_o21ai_1 _25059_ (.B1(_11446_),
    .Y(_11447_),
    .A1(net5966),
    .A2(net6310));
 sg13g2_nand2_1 _25060_ (.Y(_11448_),
    .A(_01357_),
    .B(net6358));
 sg13g2_o21ai_1 _25061_ (.B1(_11448_),
    .Y(_11449_),
    .A1(net5925),
    .A2(net6358));
 sg13g2_nand2_1 _25062_ (.Y(_11450_),
    .A(_01356_),
    .B(net6306));
 sg13g2_o21ai_1 _25063_ (.B1(_11450_),
    .Y(_11451_),
    .A1(net6013),
    .A2(net6306));
 sg13g2_nand2_1 _25064_ (.Y(_11452_),
    .A(_01355_),
    .B(net6304));
 sg13g2_o21ai_1 _25065_ (.B1(_11452_),
    .Y(_11453_),
    .A1(net5958),
    .A2(_11399_));
 sg13g2_nand2_1 _25066_ (.Y(_11454_),
    .A(_01354_),
    .B(net6306));
 sg13g2_o21ai_1 _25067_ (.B1(_11454_),
    .Y(_11455_),
    .A1(net6009),
    .A2(net6306));
 sg13g2_nand2_1 _25068_ (.Y(_11456_),
    .A(_01353_),
    .B(net6305));
 sg13g2_o21ai_1 _25069_ (.B1(_11456_),
    .Y(_11457_),
    .A1(net6003),
    .A2(net6305));
 sg13g2_nand2_1 _25070_ (.Y(_11458_),
    .A(_01352_),
    .B(net6309));
 sg13g2_o21ai_1 _25071_ (.B1(_11458_),
    .Y(_11459_),
    .A1(net6119),
    .A2(net6309));
 sg13g2_nand2_1 _25072_ (.Y(_11460_),
    .A(_01351_),
    .B(net6306));
 sg13g2_o21ai_1 _25073_ (.B1(_11460_),
    .Y(_11461_),
    .A1(net6030),
    .A2(net6306));
 sg13g2_nand2_1 _25074_ (.Y(_11462_),
    .A(_01350_),
    .B(net6309));
 sg13g2_o21ai_1 _25075_ (.B1(_11462_),
    .Y(_11463_),
    .A1(net6113),
    .A2(net6309));
 sg13g2_nand2_1 _25076_ (.Y(_11464_),
    .A(_01349_),
    .B(net6309));
 sg13g2_o21ai_1 _25077_ (.B1(_11464_),
    .Y(_11465_),
    .A1(net6025),
    .A2(net6309));
 sg13g2_nand2_1 _25078_ (.Y(_11466_),
    .A(_01348_),
    .B(net6305));
 sg13g2_o21ai_1 _25079_ (.B1(_11466_),
    .Y(_11467_),
    .A1(net6053),
    .A2(net6305));
 sg13g2_nand2_1 _25080_ (.Y(_11468_),
    .A(_01347_),
    .B(net6306));
 sg13g2_o21ai_1 _25081_ (.B1(_11468_),
    .Y(_11469_),
    .A1(net6020),
    .A2(net6306));
 sg13g2_nand2_1 _25082_ (.Y(_11470_),
    .A(_01346_),
    .B(net6360));
 sg13g2_o21ai_1 _25083_ (.B1(_11470_),
    .Y(_11471_),
    .A1(net5962),
    .A2(net6360));
 sg13g2_nand2_1 _25084_ (.Y(_11472_),
    .A(_01345_),
    .B(net6307));
 sg13g2_o21ai_1 _25085_ (.B1(_11472_),
    .Y(_11473_),
    .A1(net6104),
    .A2(net6305));
 sg13g2_mux4_1 _25086_ (.S0(net7766),
    .A0(_01066_),
    .A1(_01101_),
    .A2(_01136_),
    .A3(_01172_),
    .S1(net7723),
    .X(_11474_));
 sg13g2_nand2_1 _25087_ (.Y(_11475_),
    .A(_01344_),
    .B(net6304));
 sg13g2_o21ai_1 _25088_ (.B1(_11475_),
    .Y(_11476_),
    .A1(net5867),
    .A2(net6098));
 sg13g2_nor2b_1 _25089_ (.A(_01887_),
    .B_N(_01917_),
    .Y(_11477_));
 sg13g2_nand2b_1 _25090_ (.Y(_11478_),
    .B(net7666),
    .A_N(net7932));
 sg13g2_nand4_1 _25091_ (.B(net6466),
    .C(_09681_),
    .A(net7669),
    .Y(_11479_),
    .D(_11477_));
 sg13g2_nor2_1 _25092_ (.A(_08389_),
    .B(_11474_),
    .Y(_11480_));
 sg13g2_nand2_1 _25093_ (.Y(_11481_),
    .A(_09683_),
    .B(net7446));
 sg13g2_nand2_1 _25094_ (.Y(_11482_),
    .A(_01343_),
    .B(net6303));
 sg13g2_o21ai_1 _25095_ (.B1(_11482_),
    .Y(_11483_),
    .A1(net8286),
    .A2(net6303));
 sg13g2_nand2_1 _25096_ (.Y(_11484_),
    .A(_01342_),
    .B(net6302));
 sg13g2_nand2b_1 _25097_ (.Y(_11485_),
    .B(net6383),
    .A_N(net6302));
 sg13g2_o21ai_1 _25098_ (.B1(_11484_),
    .Y(_11486_),
    .A1(net5857),
    .A2(_11485_));
 sg13g2_nand2_1 _25099_ (.Y(_11487_),
    .A(_01341_),
    .B(net6296));
 sg13g2_o21ai_1 _25100_ (.B1(_11487_),
    .Y(_11488_),
    .A1(net5807),
    .A2(net5997));
 sg13g2_nand2_1 _25101_ (.Y(_11489_),
    .A(_01340_),
    .B(net6301));
 sg13g2_o21ai_1 _25102_ (.B1(_11489_),
    .Y(_11490_),
    .A1(net5850),
    .A2(net6301));
 sg13g2_nand2_1 _25103_ (.Y(_11491_),
    .A(_01339_),
    .B(net6300));
 sg13g2_o21ai_1 _25104_ (.B1(_11491_),
    .Y(_11492_),
    .A1(net5801),
    .A2(net6300));
 sg13g2_nand2_1 _25105_ (.Y(_11493_),
    .A(_01338_),
    .B(net6296));
 sg13g2_o21ai_1 _25106_ (.B1(_11493_),
    .Y(_11494_),
    .A1(net5796),
    .A2(_11481_));
 sg13g2_nand2_1 _25107_ (.Y(_11495_),
    .A(_01337_),
    .B(_11479_));
 sg13g2_nand2b_1 _25108_ (.Y(_11496_),
    .B(net6380),
    .A_N(_11479_));
 sg13g2_o21ai_1 _25109_ (.B1(_11495_),
    .Y(_11497_),
    .A1(net5919),
    .A2(_11496_));
 sg13g2_nand2_1 _25110_ (.Y(_11498_),
    .A(_01336_),
    .B(net6295));
 sg13g2_o21ai_1 _25111_ (.B1(_11498_),
    .Y(_11499_),
    .A1(net5790),
    .A2(_11481_));
 sg13g2_nand2_1 _25112_ (.Y(_11500_),
    .A(_01335_),
    .B(net6359));
 sg13g2_o21ai_1 _25113_ (.B1(_11500_),
    .Y(_11501_),
    .A1(net6014),
    .A2(net6359));
 sg13g2_nand2_1 _25114_ (.Y(_11502_),
    .A(_01334_),
    .B(net6303));
 sg13g2_nand2b_1 _25115_ (.Y(_11503_),
    .B(net6371),
    .A_N(net6303));
 sg13g2_o21ai_1 _25116_ (.B1(_11502_),
    .Y(_11504_),
    .A1(net5913),
    .A2(_11503_));
 sg13g2_nand2_1 _25117_ (.Y(_11505_),
    .A(_01333_),
    .B(net6296));
 sg13g2_o21ai_1 _25118_ (.B1(_11505_),
    .Y(_11506_),
    .A1(net5781),
    .A2(net5997));
 sg13g2_nand2_1 _25119_ (.Y(_11507_),
    .A(_01332_),
    .B(net6303));
 sg13g2_nand2b_1 _25120_ (.Y(_11508_),
    .B(_10493_),
    .A_N(net6303));
 sg13g2_o21ai_1 _25121_ (.B1(_11507_),
    .Y(_11509_),
    .A1(net5908),
    .A2(_11508_));
 sg13g2_mux2_1 _25122_ (.A0(net5842),
    .A1(_01331_),
    .S(_11481_),
    .X(_11510_));
 sg13g2_nand2_1 _25123_ (.Y(_11511_),
    .A(_01330_),
    .B(net6295));
 sg13g2_o21ai_1 _25124_ (.B1(_11511_),
    .Y(_11512_),
    .A1(net5835),
    .A2(_11481_));
 sg13g2_nand2_1 _25125_ (.Y(_11513_),
    .A(_01329_),
    .B(net6295));
 sg13g2_o21ai_1 _25126_ (.B1(_11513_),
    .Y(_11514_),
    .A1(net5901),
    .A2(_11481_));
 sg13g2_nand2_1 _25127_ (.Y(_11515_),
    .A(_01328_),
    .B(net6296));
 sg13g2_o21ai_1 _25128_ (.B1(_11515_),
    .Y(_11516_),
    .A1(net5896),
    .A2(net5997));
 sg13g2_nand2_1 _25129_ (.Y(_11517_),
    .A(_01327_),
    .B(net6295));
 sg13g2_o21ai_1 _25130_ (.B1(_11517_),
    .Y(_11518_),
    .A1(net5893),
    .A2(net6295));
 sg13g2_mux2_1 _25131_ (.A0(net5776),
    .A1(_01326_),
    .S(net6303),
    .X(_11519_));
 sg13g2_mux4_1 _25132_ (.S0(net7766),
    .A0(_01207_),
    .A1(_01242_),
    .A2(_01277_),
    .A3(_01312_),
    .S1(net7723),
    .X(_11520_));
 sg13g2_nand2_1 _25133_ (.Y(_11521_),
    .A(_01325_),
    .B(net6297));
 sg13g2_o21ai_1 _25134_ (.B1(_11521_),
    .Y(_11522_),
    .A1(net5883),
    .A2(net6297));
 sg13g2_nand2_1 _25135_ (.Y(_11523_),
    .A(_01324_),
    .B(net6363));
 sg13g2_nor2_1 _25136_ (.A(net7587),
    .B(_11520_),
    .Y(_11524_));
 sg13g2_o21ai_1 _25137_ (.B1(_11523_),
    .Y(_11525_),
    .A1(net5957),
    .A2(net6000));
 sg13g2_nand2_1 _25138_ (.Y(_11526_),
    .A(_01323_),
    .B(net6301));
 sg13g2_o21ai_1 _25139_ (.B1(_11526_),
    .Y(_11527_),
    .A1(net5927),
    .A2(net6301));
 sg13g2_nand2_1 _25140_ (.Y(_11528_),
    .A(_01322_),
    .B(net6300));
 sg13g2_o21ai_1 _25141_ (.B1(_11528_),
    .Y(_11529_),
    .A1(net5965),
    .A2(net6300));
 sg13g2_nand2_1 _25142_ (.Y(_11530_),
    .A(_01321_),
    .B(net6298));
 sg13g2_o21ai_1 _25143_ (.B1(_11530_),
    .Y(_11531_),
    .A1(net6013),
    .A2(net6298));
 sg13g2_nand2_1 _25144_ (.Y(_11532_),
    .A(_01320_),
    .B(net6296));
 sg13g2_o21ai_1 _25145_ (.B1(_11532_),
    .Y(_11533_),
    .A1(net5960),
    .A2(_11481_));
 sg13g2_nand2_1 _25146_ (.Y(_11534_),
    .A(_01319_),
    .B(net6298));
 sg13g2_o21ai_1 _25147_ (.B1(_11534_),
    .Y(_11535_),
    .A1(net6008),
    .A2(net6298));
 sg13g2_nand2_1 _25148_ (.Y(_11536_),
    .A(_01318_),
    .B(net6299));
 sg13g2_o21ai_1 _25149_ (.B1(_11536_),
    .Y(_11537_),
    .A1(net6003),
    .A2(net6297));
 sg13g2_nand2_1 _25150_ (.Y(_11538_),
    .A(_01317_),
    .B(net6301));
 sg13g2_o21ai_1 _25151_ (.B1(_11538_),
    .Y(_11539_),
    .A1(net6120),
    .A2(net6301));
 sg13g2_nand2_1 _25152_ (.Y(_11540_),
    .A(_01316_),
    .B(net6298));
 sg13g2_o21ai_1 _25153_ (.B1(_11540_),
    .Y(_11541_),
    .A1(net6029),
    .A2(net6298));
 sg13g2_nand2_1 _25154_ (.Y(_11542_),
    .A(_01315_),
    .B(net6302));
 sg13g2_o21ai_1 _25155_ (.B1(_11542_),
    .Y(_11543_),
    .A1(net6111),
    .A2(net6300));
 sg13g2_nand2_1 _25156_ (.Y(_11544_),
    .A(_01314_),
    .B(net6301));
 sg13g2_mux2_1 _25157_ (.A0(_01348_),
    .A1(_01383_),
    .S(net7766),
    .X(_11545_));
 sg13g2_o21ai_1 _25158_ (.B1(_11544_),
    .Y(_11546_),
    .A1(net6025),
    .A2(net6301));
 sg13g2_nand2_1 _25159_ (.Y(_11547_),
    .A(_01313_),
    .B(net6359));
 sg13g2_o21ai_1 _25160_ (.B1(_11547_),
    .Y(_11548_),
    .A1(net6010),
    .A2(net6359));
 sg13g2_nor3_1 _25161_ (.A(net7579),
    .B(net7559),
    .C(_11545_),
    .Y(_11549_));
 sg13g2_nand2_1 _25162_ (.Y(_11550_),
    .A(_01312_),
    .B(net6297));
 sg13g2_o21ai_1 _25163_ (.B1(_11550_),
    .Y(_11551_),
    .A1(net6052),
    .A2(net6297));
 sg13g2_nand2_1 _25164_ (.Y(_11552_),
    .A(_01311_),
    .B(net6299));
 sg13g2_o21ai_1 _25165_ (.B1(_11552_),
    .Y(_11553_),
    .A1(net6019),
    .A2(net6299));
 sg13g2_nand2_1 _25166_ (.Y(_11554_),
    .A(_01310_),
    .B(net6298));
 sg13g2_o21ai_1 _25167_ (.B1(_11554_),
    .Y(_11555_),
    .A1(net6104),
    .A2(net6298));
 sg13g2_nand2_1 _25168_ (.Y(_11556_),
    .A(_01309_),
    .B(net6296));
 sg13g2_o21ai_1 _25169_ (.B1(_11556_),
    .Y(_11557_),
    .A1(net5866),
    .A2(net5997));
 sg13g2_nand4_1 _25170_ (.B(_09604_),
    .C(_10091_),
    .A(net7670),
    .Y(_11558_),
    .D(_11477_));
 sg13g2_nand2_1 _25171_ (.Y(_11559_),
    .A(_10094_),
    .B(net7446));
 sg13g2_nand2_1 _25172_ (.Y(_11560_),
    .A(_01308_),
    .B(net6294));
 sg13g2_o21ai_1 _25173_ (.B1(_11560_),
    .Y(_11561_),
    .A1(net8287),
    .A2(net6294));
 sg13g2_nand2_1 _25174_ (.Y(_11562_),
    .A(_01307_),
    .B(net6293));
 sg13g2_nand2b_1 _25175_ (.Y(_11563_),
    .B(net6383),
    .A_N(net6293));
 sg13g2_o21ai_1 _25176_ (.B1(_11562_),
    .Y(_11564_),
    .A1(net5857),
    .A2(_11563_));
 sg13g2_nand2_1 _25177_ (.Y(_11565_),
    .A(_01306_),
    .B(net6287));
 sg13g2_o21ai_1 _25178_ (.B1(_11565_),
    .Y(_11566_),
    .A1(net5807),
    .A2(_11559_));
 sg13g2_nand2_1 _25179_ (.Y(_11567_),
    .A(_01305_),
    .B(net6291));
 sg13g2_o21ai_1 _25180_ (.B1(_11567_),
    .Y(_11568_),
    .A1(net5850),
    .A2(net6291));
 sg13g2_nand2_1 _25181_ (.Y(_11569_),
    .A(_01304_),
    .B(net6292));
 sg13g2_o21ai_1 _25182_ (.B1(_11569_),
    .Y(_11570_),
    .A1(net5801),
    .A2(net6292));
 sg13g2_mux2_1 _25183_ (.A0(_01559_),
    .A1(_01594_),
    .S(net7766),
    .X(_11571_));
 sg13g2_nand2_1 _25184_ (.Y(_11572_),
    .A(_01303_),
    .B(net6286));
 sg13g2_o21ai_1 _25185_ (.B1(_11572_),
    .Y(_11573_),
    .A1(net5796),
    .A2(net5996));
 sg13g2_nand2_1 _25186_ (.Y(_11574_),
    .A(_01302_),
    .B(net6359));
 sg13g2_nor2_1 _25187_ (.A(net7551),
    .B(_11571_),
    .Y(_11575_));
 sg13g2_o21ai_1 _25188_ (.B1(_11574_),
    .Y(_11576_),
    .A1(net6006),
    .A2(net6359));
 sg13g2_nand2_1 _25189_ (.Y(_11577_),
    .A(_01301_),
    .B(net6293));
 sg13g2_nand2b_1 _25190_ (.Y(_11578_),
    .B(net6380),
    .A_N(net6290));
 sg13g2_o21ai_1 _25191_ (.B1(_11577_),
    .Y(_11579_),
    .A1(net5919),
    .A2(_11578_));
 sg13g2_nand2_1 _25192_ (.Y(_11580_),
    .A(_01300_),
    .B(net6286));
 sg13g2_o21ai_1 _25193_ (.B1(_11580_),
    .Y(_11581_),
    .A1(net5790),
    .A2(net5996));
 sg13g2_nand2_1 _25194_ (.Y(_11582_),
    .A(_01299_),
    .B(net6294));
 sg13g2_nand2b_1 _25195_ (.Y(_11583_),
    .B(net6371),
    .A_N(net6294));
 sg13g2_o21ai_1 _25196_ (.B1(_11582_),
    .Y(_11584_),
    .A1(net5913),
    .A2(_11583_));
 sg13g2_nand2_1 _25197_ (.Y(_11585_),
    .A(_01298_),
    .B(net6287));
 sg13g2_o21ai_1 _25198_ (.B1(_11585_),
    .Y(_11586_),
    .A1(net5781),
    .A2(_11559_));
 sg13g2_nand2_1 _25199_ (.Y(_11587_),
    .A(_01297_),
    .B(net6294));
 sg13g2_nand2b_1 _25200_ (.Y(_11588_),
    .B(_10493_),
    .A_N(net6294));
 sg13g2_o21ai_1 _25201_ (.B1(_11587_),
    .Y(_11589_),
    .A1(net5908),
    .A2(_11588_));
 sg13g2_mux2_1 _25202_ (.A0(net5842),
    .A1(_01296_),
    .S(_11559_),
    .X(_11590_));
 sg13g2_nand2_1 _25203_ (.Y(_11591_),
    .A(_01295_),
    .B(net6286));
 sg13g2_o21ai_1 _25204_ (.B1(_11591_),
    .Y(_11592_),
    .A1(net5835),
    .A2(net5996));
 sg13g2_nand2_1 _25205_ (.Y(_11593_),
    .A(_01294_),
    .B(net6286));
 sg13g2_o21ai_1 _25206_ (.B1(_11593_),
    .Y(_11594_),
    .A1(net5901),
    .A2(net5996));
 sg13g2_nand2_1 _25207_ (.Y(_11595_),
    .A(_01293_),
    .B(net6287));
 sg13g2_o21ai_1 _25208_ (.B1(_11595_),
    .Y(_11596_),
    .A1(net5896),
    .A2(_11559_));
 sg13g2_nand2_1 _25209_ (.Y(_11597_),
    .A(_01292_),
    .B(net6286));
 sg13g2_mux2_1 _25210_ (.A0(_01418_),
    .A1(_01453_),
    .S(net7766),
    .X(_11598_));
 sg13g2_o21ai_1 _25211_ (.B1(_11597_),
    .Y(_11599_),
    .A1(net5893),
    .A2(net6286));
 sg13g2_nand2_1 _25212_ (.Y(_11600_),
    .A(_01291_),
    .B(net6361));
 sg13g2_o21ai_1 _25213_ (.B1(_11600_),
    .Y(_11601_),
    .A1(_09678_),
    .A2(net6361));
 sg13g2_nor3_1 _25214_ (.A(net7579),
    .B(net7567),
    .C(_11598_),
    .Y(_11602_));
 sg13g2_mux2_1 _25215_ (.A0(net5776),
    .A1(_01290_),
    .S(net6294),
    .X(_11603_));
 sg13g2_nand2_1 _25216_ (.Y(_11604_),
    .A(_01289_),
    .B(net6288));
 sg13g2_o21ai_1 _25217_ (.B1(_11604_),
    .Y(_11605_),
    .A1(net5883),
    .A2(net6288));
 sg13g2_nand2_1 _25218_ (.Y(_11606_),
    .A(_01288_),
    .B(net6291));
 sg13g2_o21ai_1 _25219_ (.B1(_11606_),
    .Y(_11607_),
    .A1(net5927),
    .A2(net6291));
 sg13g2_nand2_1 _25220_ (.Y(_11608_),
    .A(_01287_),
    .B(net6292));
 sg13g2_o21ai_1 _25221_ (.B1(_11608_),
    .Y(_11609_),
    .A1(net5965),
    .A2(net6292));
 sg13g2_nand2_1 _25222_ (.Y(_11610_),
    .A(_01286_),
    .B(net6289));
 sg13g2_o21ai_1 _25223_ (.B1(_11610_),
    .Y(_11611_),
    .A1(net6013),
    .A2(net6289));
 sg13g2_nand2_1 _25224_ (.Y(_11612_),
    .A(_01285_),
    .B(net6287));
 sg13g2_o21ai_1 _25225_ (.B1(_11612_),
    .Y(_11613_),
    .A1(net5960),
    .A2(_11559_));
 sg13g2_nand2_1 _25226_ (.Y(_11614_),
    .A(_01284_),
    .B(net6289));
 sg13g2_o21ai_1 _25227_ (.B1(_11614_),
    .Y(_11615_),
    .A1(net6008),
    .A2(net6289));
 sg13g2_nand2_1 _25228_ (.Y(_11616_),
    .A(_01283_),
    .B(net6289));
 sg13g2_o21ai_1 _25229_ (.B1(_11616_),
    .Y(_11617_),
    .A1(net6003),
    .A2(net6288));
 sg13g2_nand2_1 _25230_ (.Y(_11618_),
    .A(_01282_),
    .B(net6291));
 sg13g2_o21ai_1 _25231_ (.B1(_11618_),
    .Y(_11619_),
    .A1(net6120),
    .A2(net6291));
 sg13g2_nand2_1 _25232_ (.Y(_11620_),
    .A(_01281_),
    .B(net6289));
 sg13g2_o21ai_1 _25233_ (.B1(_11620_),
    .Y(_11621_),
    .A1(net6029),
    .A2(net6289));
 sg13g2_nand2_1 _25234_ (.Y(_11622_),
    .A(_01280_),
    .B(net6360));
 sg13g2_mux2_1 _25235_ (.A0(_01488_),
    .A1(_01524_),
    .S(net7766),
    .X(_11623_));
 sg13g2_o21ai_1 _25236_ (.B1(_11622_),
    .Y(_11624_),
    .A1(net6033),
    .A2(net6360));
 sg13g2_nand2_1 _25237_ (.Y(_11625_),
    .A(_01279_),
    .B(net6293));
 sg13g2_o21ai_1 _25238_ (.B1(_11625_),
    .Y(_11626_),
    .A1(net6111),
    .A2(net6293));
 sg13g2_nor3_1 _25239_ (.A(net7579),
    .B(net7563),
    .C(_11623_),
    .Y(_11627_));
 sg13g2_nand2_1 _25240_ (.Y(_11628_),
    .A(_01278_),
    .B(net6291));
 sg13g2_o21ai_1 _25241_ (.B1(_11628_),
    .Y(_11629_),
    .A1(net6025),
    .A2(net6291));
 sg13g2_nand2_1 _25242_ (.Y(_11630_),
    .A(_01277_),
    .B(net6288));
 sg13g2_o21ai_1 _25243_ (.B1(_11630_),
    .Y(_11631_),
    .A1(net6052),
    .A2(net6288));
 sg13g2_nand2_1 _25244_ (.Y(_11632_),
    .A(_01276_),
    .B(net6290));
 sg13g2_o21ai_1 _25245_ (.B1(_11632_),
    .Y(_11633_),
    .A1(net6019),
    .A2(net6290));
 sg13g2_nand2_1 _25246_ (.Y(_11634_),
    .A(_01275_),
    .B(net6288));
 sg13g2_o21ai_1 _25247_ (.B1(_11634_),
    .Y(_11635_),
    .A1(net6105),
    .A2(net6288));
 sg13g2_nand2_1 _25248_ (.Y(_11636_),
    .A(_01274_),
    .B(net6287));
 sg13g2_o21ai_1 _25249_ (.B1(_11636_),
    .Y(_11637_),
    .A1(net5866),
    .A2(_11559_));
 sg13g2_or4_1 _25250_ (.A(net7667),
    .B(net6468),
    .C(_09682_),
    .D(_11478_),
    .X(_11638_));
 sg13g2_nand2_1 _25251_ (.Y(_11639_),
    .A(net6346),
    .B(net7446));
 sg13g2_nand2_1 _25252_ (.Y(_11640_),
    .A(_01273_),
    .B(net6278));
 sg13g2_o21ai_1 _25253_ (.B1(_11640_),
    .Y(_11641_),
    .A1(net8287),
    .A2(net6278));
 sg13g2_nand2_1 _25254_ (.Y(_11642_),
    .A(_01272_),
    .B(net6284));
 sg13g2_nand2b_1 _25255_ (.Y(_11643_),
    .B(net6383),
    .A_N(net6284));
 sg13g2_o21ai_1 _25256_ (.B1(_11642_),
    .Y(_11644_),
    .A1(net5857),
    .A2(_11643_));
 sg13g2_nand2_1 _25257_ (.Y(_11645_),
    .A(_01271_),
    .B(net6277));
 sg13g2_o21ai_1 _25258_ (.B1(_11645_),
    .Y(_11646_),
    .A1(net5807),
    .A2(net6097));
 sg13g2_nand2_1 _25259_ (.Y(_11647_),
    .A(_01270_),
    .B(net6283));
 sg13g2_or4_1 _25260_ (.A(_11549_),
    .B(_11575_),
    .C(_11602_),
    .D(_11627_),
    .X(_11648_));
 sg13g2_o21ai_1 _25261_ (.B1(_11647_),
    .Y(_11649_),
    .A1(net5850),
    .A2(net6283));
 sg13g2_nand2_1 _25262_ (.Y(_11650_),
    .A(_01269_),
    .B(net6358));
 sg13g2_o21ai_1 _25263_ (.B1(_11650_),
    .Y(_11651_),
    .A1(net6110),
    .A2(net6358));
 sg13g2_nand2_1 _25264_ (.Y(_11652_),
    .A(_01268_),
    .B(net6282));
 sg13g2_o21ai_1 _25265_ (.B1(_11652_),
    .Y(_11653_),
    .A1(net5801),
    .A2(net6282));
 sg13g2_nand2_1 _25266_ (.Y(_11654_),
    .A(_01267_),
    .B(_11638_));
 sg13g2_o21ai_1 _25267_ (.B1(_11654_),
    .Y(_11655_),
    .A1(net5796),
    .A2(net6097));
 sg13g2_nand2_1 _25268_ (.Y(_11656_),
    .A(_01266_),
    .B(net6285));
 sg13g2_nand2b_1 _25269_ (.Y(_11657_),
    .B(net6380),
    .A_N(net6285));
 sg13g2_o21ai_1 _25270_ (.B1(_11656_),
    .Y(_11658_),
    .A1(net5919),
    .A2(_11657_));
 sg13g2_nand2_1 _25271_ (.Y(_11659_),
    .A(_01265_),
    .B(net6277));
 sg13g2_nor3_1 _25272_ (.A(_11480_),
    .B(_11524_),
    .C(_11648_),
    .Y(_11660_));
 sg13g2_o21ai_1 _25273_ (.B1(_11659_),
    .Y(_11661_),
    .A1(net5790),
    .A2(net6097));
 sg13g2_nand2_1 _25274_ (.Y(_11662_),
    .A(_01264_),
    .B(net6278));
 sg13g2_nand2b_1 _25275_ (.Y(_11663_),
    .B(net6371),
    .A_N(net6278));
 sg13g2_o21ai_1 _25276_ (.B1(_11662_),
    .Y(_11664_),
    .A1(net5916),
    .A2(_11663_));
 sg13g2_and2_1 _25277_ (.A(_11432_),
    .B(_11660_),
    .X(_11665_));
 sg13g2_nand2_1 _25278_ (.Y(_11666_),
    .A(_01263_),
    .B(net6277));
 sg13g2_o21ai_1 _25279_ (.B1(_11666_),
    .Y(_11667_),
    .A1(net5781),
    .A2(net6097));
 sg13g2_nand2_1 _25280_ (.Y(_11668_),
    .A(_01262_),
    .B(net6278));
 sg13g2_nand2b_1 _25281_ (.Y(_11669_),
    .B(_10493_),
    .A_N(net6278));
 sg13g2_o21ai_1 _25282_ (.B1(_11668_),
    .Y(_11670_),
    .A1(net5908),
    .A2(_11669_));
 sg13g2_mux2_1 _25283_ (.A0(net5842),
    .A1(_01261_),
    .S(_11639_),
    .X(_11671_));
 sg13g2_nand2_1 _25284_ (.Y(_11672_),
    .A(_01260_),
    .B(_11638_));
 sg13g2_o21ai_1 _25285_ (.B1(_11672_),
    .Y(_11673_),
    .A1(net5835),
    .A2(net6097));
 sg13g2_nand2_1 _25286_ (.Y(_11674_),
    .A(_01259_),
    .B(net6277));
 sg13g2_o21ai_1 _25287_ (.B1(_11674_),
    .Y(_11675_),
    .A1(net5901),
    .A2(net6097));
 sg13g2_nand2_1 _25288_ (.Y(_11676_),
    .A(_01258_),
    .B(net6361));
 sg13g2_o21ai_1 _25289_ (.B1(_11676_),
    .Y(_11677_),
    .A1(_09902_),
    .A2(net6361));
 sg13g2_nand2_1 _25290_ (.Y(_11678_),
    .A(_01257_),
    .B(net6277));
 sg13g2_o21ai_1 _25291_ (.B1(_08634_),
    .Y(_11679_),
    .A1(_08616_),
    .A2(_11665_));
 sg13g2_o21ai_1 _25292_ (.B1(_11678_),
    .Y(_11680_),
    .A1(net5896),
    .A2(net6097));
 sg13g2_nand2_1 _25293_ (.Y(_11681_),
    .A(_01256_),
    .B(_11638_));
 sg13g2_a21oi_1 _25294_ (.A1(_08616_),
    .A2(_11223_),
    .Y(_11682_),
    .B1(_11679_));
 sg13g2_o21ai_1 _25295_ (.B1(_11681_),
    .Y(_11683_),
    .A1(net5893),
    .A2(_11638_));
 sg13g2_inv_1 _25296_ (.Y(_11684_),
    .A(net6953));
 sg13g2_mux2_1 _25297_ (.A0(net5774),
    .A1(_01255_),
    .S(net6278),
    .X(_11685_));
 sg13g2_nand2_1 _25298_ (.Y(_11686_),
    .A(_01254_),
    .B(net6280));
 sg13g2_o21ai_1 _25299_ (.B1(_11686_),
    .Y(_11687_),
    .A1(net5883),
    .A2(net6280));
 sg13g2_nand2_1 _25300_ (.Y(_11688_),
    .A(_01253_),
    .B(net6283));
 sg13g2_o21ai_1 _25301_ (.B1(_11688_),
    .Y(_11689_),
    .A1(net5927),
    .A2(net6283));
 sg13g2_nand2_1 _25302_ (.Y(_11690_),
    .A(_01252_),
    .B(net6282));
 sg13g2_o21ai_1 _25303_ (.B1(_11690_),
    .Y(_11691_),
    .A1(net5964),
    .A2(net6282));
 sg13g2_nand2_1 _25304_ (.Y(_11692_),
    .A(_01251_),
    .B(net6282));
 sg13g2_o21ai_1 _25305_ (.B1(_11692_),
    .Y(_11693_),
    .A1(net6013),
    .A2(net6282));
 sg13g2_nand2_1 _25306_ (.Y(_11694_),
    .A(_01250_),
    .B(_11638_));
 sg13g2_o21ai_1 _25307_ (.B1(_11694_),
    .Y(_11695_),
    .A1(net5960),
    .A2(net6097));
 sg13g2_nand2_1 _25308_ (.Y(_11696_),
    .A(_01249_),
    .B(net6281));
 sg13g2_o21ai_1 _25309_ (.B1(_11696_),
    .Y(_11697_),
    .A1(net6008),
    .A2(net6279));
 sg13g2_nand2_1 _25310_ (.Y(_11698_),
    .A(_01248_),
    .B(net6280));
 sg13g2_o21ai_1 _25311_ (.B1(_11698_),
    .Y(_11699_),
    .A1(net6003),
    .A2(net6280));
 sg13g2_nand2_1 _25312_ (.Y(_11700_),
    .A(_01247_),
    .B(net6356));
 sg13g2_o21ai_1 _25313_ (.B1(_11700_),
    .Y(_11701_),
    .A1(net6055),
    .A2(net6356));
 sg13g2_nand2_1 _25314_ (.Y(_11702_),
    .A(_01246_),
    .B(net6283));
 sg13g2_o21ai_1 _25315_ (.B1(_11702_),
    .Y(_11703_),
    .A1(net6120),
    .A2(net6283));
 sg13g2_nand2_1 _25316_ (.Y(_11704_),
    .A(_01245_),
    .B(net6282));
 sg13g2_o21ai_1 _25317_ (.B1(_11704_),
    .Y(_11705_),
    .A1(_09774_),
    .A2(net6281));
 sg13g2_nand2_1 _25318_ (.Y(_11706_),
    .A(_01244_),
    .B(net6284));
 sg13g2_o21ai_1 _25319_ (.B1(_11706_),
    .Y(_11707_),
    .A1(net6111),
    .A2(net6284));
 sg13g2_nand2_1 _25320_ (.Y(_11708_),
    .A(_01243_),
    .B(net6283));
 sg13g2_o21ai_1 _25321_ (.B1(_11708_),
    .Y(_11709_),
    .A1(net6025),
    .A2(net6283));
 sg13g2_nand2_1 _25322_ (.Y(_11710_),
    .A(_01242_),
    .B(net6280));
 sg13g2_o21ai_1 _25323_ (.B1(_11710_),
    .Y(_11711_),
    .A1(net6052),
    .A2(net6280));
 sg13g2_nand2_1 _25324_ (.Y(_11712_),
    .A(_01241_),
    .B(net6279));
 sg13g2_o21ai_1 _25325_ (.B1(_11712_),
    .Y(_11713_),
    .A1(net6019),
    .A2(net6279));
 sg13g2_nand2_1 _25326_ (.Y(_11714_),
    .A(_01240_),
    .B(net6280));
 sg13g2_o21ai_1 _25327_ (.B1(_11714_),
    .Y(_11715_),
    .A1(net6105),
    .A2(net6280));
 sg13g2_nand2_1 _25328_ (.Y(_11716_),
    .A(_01239_),
    .B(_11638_));
 sg13g2_o21ai_1 _25329_ (.B1(_11716_),
    .Y(_11717_),
    .A1(net5866),
    .A2(_11639_));
 sg13g2_or4_1 _25330_ (.A(net7667),
    .B(net6467),
    .C(_10092_),
    .D(_11478_),
    .X(_11718_));
 sg13g2_nand2_1 _25331_ (.Y(_11719_),
    .A(net6335),
    .B(net7446));
 sg13g2_nand2_1 _25332_ (.Y(_11720_),
    .A(_01238_),
    .B(net6268));
 sg13g2_o21ai_1 _25333_ (.B1(_11720_),
    .Y(_11721_),
    .A1(net8287),
    .A2(net6268));
 sg13g2_nand2_1 _25334_ (.Y(_11722_),
    .A(_01237_),
    .B(net6272));
 sg13g2_nand2b_1 _25335_ (.Y(_11723_),
    .B(net6383),
    .A_N(net6274));
 sg13g2_o21ai_1 _25336_ (.B1(_11722_),
    .Y(_11724_),
    .A1(net5857),
    .A2(_11723_));
 sg13g2_mux2_1 _25337_ (.A0(_01559_),
    .A1(_01594_),
    .S(net7915),
    .X(_11725_));
 sg13g2_nand2_1 _25338_ (.Y(_11726_),
    .A(_01236_),
    .B(net6360));
 sg13g2_o21ai_1 _25339_ (.B1(_11726_),
    .Y(_11727_),
    .A1(net6022),
    .A2(net6360));
 sg13g2_nor2_1 _25340_ (.A(net7449),
    .B(_11725_),
    .Y(_11728_));
 sg13g2_nand2_1 _25341_ (.Y(_11729_),
    .A(_01235_),
    .B(net6276));
 sg13g2_o21ai_1 _25342_ (.B1(_11729_),
    .Y(_11730_),
    .A1(net5807),
    .A2(net6096));
 sg13g2_nand2_1 _25343_ (.Y(_11731_),
    .A(_01234_),
    .B(net6271));
 sg13g2_o21ai_1 _25344_ (.B1(_11731_),
    .Y(_11732_),
    .A1(net5850),
    .A2(net6271));
 sg13g2_nand2_1 _25345_ (.Y(_11733_),
    .A(_01233_),
    .B(net6273));
 sg13g2_o21ai_1 _25346_ (.B1(_11733_),
    .Y(_11734_),
    .A1(net5801),
    .A2(net6273));
 sg13g2_nand2_1 _25347_ (.Y(_11735_),
    .A(_01232_),
    .B(net6275));
 sg13g2_o21ai_1 _25348_ (.B1(_11735_),
    .Y(_11736_),
    .A1(net5796),
    .A2(net6096));
 sg13g2_nand2b_1 _25349_ (.Y(_11737_),
    .B(net6380),
    .A_N(net6270));
 sg13g2_nand2_1 _25350_ (.Y(_11738_),
    .A(_01231_),
    .B(net6270));
 sg13g2_o21ai_1 _25351_ (.B1(_11738_),
    .Y(_11739_),
    .A1(net5919),
    .A2(_11737_));
 sg13g2_nand2_1 _25352_ (.Y(_11740_),
    .A(_01230_),
    .B(net6275));
 sg13g2_o21ai_1 _25353_ (.B1(_11740_),
    .Y(_11741_),
    .A1(net5790),
    .A2(net6096));
 sg13g2_nand2b_1 _25354_ (.Y(_11742_),
    .B(net6371),
    .A_N(net6268));
 sg13g2_nand2_1 _25355_ (.Y(_11743_),
    .A(_01229_),
    .B(net6268));
 sg13g2_o21ai_1 _25356_ (.B1(_11743_),
    .Y(_11744_),
    .A1(net5916),
    .A2(_11742_));
 sg13g2_nand2_1 _25357_ (.Y(_11745_),
    .A(_01228_),
    .B(net6276));
 sg13g2_o21ai_1 _25358_ (.B1(_11745_),
    .Y(_11746_),
    .A1(net5781),
    .A2(net6096));
 sg13g2_nand2b_1 _25359_ (.Y(_11747_),
    .B(_10493_),
    .A_N(_11718_));
 sg13g2_nand2_1 _25360_ (.Y(_11748_),
    .A(_01227_),
    .B(net6268));
 sg13g2_o21ai_1 _25361_ (.B1(_11748_),
    .Y(_11749_),
    .A1(net5908),
    .A2(_11747_));
 sg13g2_mux2_1 _25362_ (.A0(net5842),
    .A1(_01226_),
    .S(_11719_),
    .X(_11750_));
 sg13g2_nand2_1 _25363_ (.Y(_11751_),
    .A(_01225_),
    .B(net6362));
 sg13g2_mux2_1 _25364_ (.A0(_01488_),
    .A1(_01524_),
    .S(net7915),
    .X(_11752_));
 sg13g2_o21ai_1 _25365_ (.B1(_11751_),
    .Y(_11753_),
    .A1(net6108),
    .A2(net6362));
 sg13g2_nand2_1 _25366_ (.Y(_11754_),
    .A(_01224_),
    .B(net6275));
 sg13g2_o21ai_1 _25367_ (.B1(_11754_),
    .Y(_11755_),
    .A1(net5835),
    .A2(net6096));
 sg13g2_nor3_1 _25368_ (.A(_09028_),
    .B(net7487),
    .C(_11752_),
    .Y(_11756_));
 sg13g2_nand2_1 _25369_ (.Y(_11757_),
    .A(_01223_),
    .B(net6275));
 sg13g2_o21ai_1 _25370_ (.B1(_11757_),
    .Y(_11758_),
    .A1(net5901),
    .A2(net6096));
 sg13g2_nand2_1 _25371_ (.Y(_11759_),
    .A(_01222_),
    .B(net6276));
 sg13g2_o21ai_1 _25372_ (.B1(_11759_),
    .Y(_11760_),
    .A1(net5896),
    .A2(net6096));
 sg13g2_nand2_1 _25373_ (.Y(_11761_),
    .A(_01221_),
    .B(net6275));
 sg13g2_o21ai_1 _25374_ (.B1(_11761_),
    .Y(_11762_),
    .A1(net5893),
    .A2(net6275));
 sg13g2_mux2_1 _25375_ (.A0(net5774),
    .A1(_01220_),
    .S(net6268),
    .X(_11763_));
 sg13g2_nand2_1 _25376_ (.Y(_11764_),
    .A(_01219_),
    .B(net6269));
 sg13g2_o21ai_1 _25377_ (.B1(_11764_),
    .Y(_11765_),
    .A1(net5883),
    .A2(net6269));
 sg13g2_nand2_1 _25378_ (.Y(_11766_),
    .A(_01218_),
    .B(net6271));
 sg13g2_o21ai_1 _25379_ (.B1(_11766_),
    .Y(_11767_),
    .A1(net5927),
    .A2(net6271));
 sg13g2_nand2_1 _25380_ (.Y(_11768_),
    .A(_01217_),
    .B(net6273));
 sg13g2_o21ai_1 _25381_ (.B1(_11768_),
    .Y(_11769_),
    .A1(net5964),
    .A2(net6273));
 sg13g2_nand2_1 _25382_ (.Y(_11770_),
    .A(_01216_),
    .B(net6273));
 sg13g2_o21ai_1 _25383_ (.B1(_11770_),
    .Y(_11771_),
    .A1(net6014),
    .A2(net6273));
 sg13g2_nand2_1 _25384_ (.Y(_11772_),
    .A(_01215_),
    .B(net6276));
 sg13g2_o21ai_1 _25385_ (.B1(_11772_),
    .Y(_11773_),
    .A1(net5960),
    .A2(_11719_));
 sg13g2_nand2_1 _25386_ (.Y(_11774_),
    .A(_01214_),
    .B(net6363));
 sg13g2_o21ai_1 _25387_ (.B1(_11774_),
    .Y(_11775_),
    .A1(net5864),
    .A2(net6000));
 sg13g2_nand2_1 _25388_ (.Y(_11776_),
    .A(_01213_),
    .B(net6274));
 sg13g2_o21ai_1 _25389_ (.B1(_11776_),
    .Y(_11777_),
    .A1(net6008),
    .A2(net6274));
 sg13g2_nand2_1 _25390_ (.Y(_11778_),
    .A(_01212_),
    .B(net6269));
 sg13g2_o21ai_1 _25391_ (.B1(_11778_),
    .Y(_11779_),
    .A1(net6003),
    .A2(net6269));
 sg13g2_nand2_1 _25392_ (.Y(_11780_),
    .A(_01211_),
    .B(net6271));
 sg13g2_mux2_1 _25393_ (.A0(_00791_),
    .A1(_00823_),
    .S(net7913),
    .X(_11781_));
 sg13g2_o21ai_1 _25394_ (.B1(_11780_),
    .Y(_11782_),
    .A1(net6120),
    .A2(net6271));
 sg13g2_nand2_1 _25395_ (.Y(_11783_),
    .A(_01210_),
    .B(net6274));
 sg13g2_o21ai_1 _25396_ (.B1(_11783_),
    .Y(_11784_),
    .A1(_09774_),
    .A2(net6274));
 sg13g2_nor3_1 _25397_ (.A(net7540),
    .B(net7467),
    .C(_11781_),
    .Y(_11785_));
 sg13g2_nand2_1 _25398_ (.Y(_11786_),
    .A(_01209_),
    .B(net6272));
 sg13g2_o21ai_1 _25399_ (.B1(_11786_),
    .Y(_11787_),
    .A1(net6111),
    .A2(net6272));
 sg13g2_nand2_1 _25400_ (.Y(_11788_),
    .A(_01208_),
    .B(net6271));
 sg13g2_o21ai_1 _25401_ (.B1(_11788_),
    .Y(_11789_),
    .A1(net6025),
    .A2(net6271));
 sg13g2_nand2_1 _25402_ (.Y(_11790_),
    .A(_01207_),
    .B(net6269));
 sg13g2_o21ai_1 _25403_ (.B1(_11790_),
    .Y(_11791_),
    .A1(net6052),
    .A2(net6269));
 sg13g2_nand2_1 _25404_ (.Y(_11792_),
    .A(_01206_),
    .B(net6270));
 sg13g2_o21ai_1 _25405_ (.B1(_11792_),
    .Y(_11793_),
    .A1(net6019),
    .A2(net6270));
 sg13g2_nand2_1 _25406_ (.Y(_11794_),
    .A(_01205_),
    .B(net6269));
 sg13g2_o21ai_1 _25407_ (.B1(_11794_),
    .Y(_11795_),
    .A1(net6105),
    .A2(net6269));
 sg13g2_nand2_1 _25408_ (.Y(_11796_),
    .A(_01204_),
    .B(net6276));
 sg13g2_o21ai_1 _25409_ (.B1(_11796_),
    .Y(_11797_),
    .A1(net5866),
    .A2(_11719_));
 sg13g2_or4_1 _25410_ (.A(net7667),
    .B(_06620_),
    .C(net6468),
    .D(_09606_),
    .X(_11798_));
 sg13g2_nor3_1 _25411_ (.A(net7671),
    .B(_09603_),
    .C(_09606_),
    .Y(_11799_));
 sg13g2_nand2_1 _25412_ (.Y(_11800_),
    .A(net7627),
    .B(net6259));
 sg13g2_nand2_1 _25413_ (.Y(_11801_),
    .A(_01203_),
    .B(net6261));
 sg13g2_o21ai_1 _25414_ (.B1(_11801_),
    .Y(_11802_),
    .A1(net8286),
    .A2(net6261));
 sg13g2_nand4_1 _25415_ (.B(net7627),
    .C(net6466),
    .A(net7669),
    .Y(_11803_),
    .D(_09681_));
 sg13g2_nand2_1 _25416_ (.Y(_11804_),
    .A(_06619_),
    .B(_09683_));
 sg13g2_nand2_1 _25417_ (.Y(_11805_),
    .A(_01202_),
    .B(net6257));
 sg13g2_o21ai_1 _25418_ (.B1(_11805_),
    .Y(_11806_),
    .A1(net8287),
    .A2(net6257));
 sg13g2_nand2_1 _25419_ (.Y(_11807_),
    .A(_01201_),
    .B(net6256));
 sg13g2_nand2b_1 _25420_ (.Y(_11808_),
    .B(net6384),
    .A_N(net6258));
 sg13g2_o21ai_1 _25421_ (.B1(_11807_),
    .Y(_11809_),
    .A1(net5856),
    .A2(_11808_));
 sg13g2_nand2_1 _25422_ (.Y(_11810_),
    .A(_01200_),
    .B(net6251));
 sg13g2_mux2_1 _25423_ (.A0(_00855_),
    .A1(_00890_),
    .S(net7913),
    .X(_11811_));
 sg13g2_o21ai_1 _25424_ (.B1(_11810_),
    .Y(_11812_),
    .A1(net5807),
    .A2(_11804_));
 sg13g2_nand2_1 _25425_ (.Y(_11813_),
    .A(_01199_),
    .B(net6255));
 sg13g2_nor3_1 _25426_ (.A(net7540),
    .B(net7457),
    .C(_11811_),
    .Y(_11814_));
 sg13g2_o21ai_1 _25427_ (.B1(_11813_),
    .Y(_11815_),
    .A1(net5849),
    .A2(net6255));
 sg13g2_nand2_1 _25428_ (.Y(_11816_),
    .A(_01198_),
    .B(net6256));
 sg13g2_o21ai_1 _25429_ (.B1(_11816_),
    .Y(_11817_),
    .A1(net5801),
    .A2(net6256));
 sg13g2_nand2_1 _25430_ (.Y(_11818_),
    .A(_01197_),
    .B(net6250));
 sg13g2_o21ai_1 _25431_ (.B1(_11818_),
    .Y(_11819_),
    .A1(net5796),
    .A2(net5995));
 sg13g2_nand2_1 _25432_ (.Y(_11820_),
    .A(_01196_),
    .B(net6254));
 sg13g2_nand2b_1 _25433_ (.Y(_11821_),
    .B(net6380),
    .A_N(net6258));
 sg13g2_nor4_1 _25434_ (.A(_11728_),
    .B(_11756_),
    .C(_11785_),
    .D(_11814_),
    .Y(_11822_));
 sg13g2_o21ai_1 _25435_ (.B1(_11820_),
    .Y(_11823_),
    .A1(net5919),
    .A2(_11821_));
 sg13g2_nand2_1 _25436_ (.Y(_11824_),
    .A(_01195_),
    .B(net6250));
 sg13g2_o21ai_1 _25437_ (.B1(_11824_),
    .Y(_11825_),
    .A1(net5790),
    .A2(net5995));
 sg13g2_nand2_1 _25438_ (.Y(_11826_),
    .A(_01194_),
    .B(net6257));
 sg13g2_nand2b_1 _25439_ (.Y(_11827_),
    .B(net6371),
    .A_N(net6257));
 sg13g2_o21ai_1 _25440_ (.B1(_11826_),
    .Y(_11828_),
    .A1(net5913),
    .A2(_11827_));
 sg13g2_nand2_1 _25441_ (.Y(_11829_),
    .A(_01193_),
    .B(net6250));
 sg13g2_o21ai_1 _25442_ (.B1(_11829_),
    .Y(_11830_),
    .A1(net5781),
    .A2(_11804_));
 sg13g2_nand2_1 _25443_ (.Y(_11831_),
    .A(_01192_),
    .B(net6261));
 sg13g2_nand2b_1 _25444_ (.Y(_11832_),
    .B(net6382),
    .A_N(net6262));
 sg13g2_o21ai_1 _25445_ (.B1(_11831_),
    .Y(_11833_),
    .A1(net5854),
    .A2(_11832_));
 sg13g2_nand2_1 _25446_ (.Y(_11834_),
    .A(_01191_),
    .B(net6257));
 sg13g2_nand2b_1 _25447_ (.Y(_11835_),
    .B(net6364),
    .A_N(net6257));
 sg13g2_o21ai_1 _25448_ (.B1(_11834_),
    .Y(_11836_),
    .A1(net5907),
    .A2(_11835_));
 sg13g2_mux2_1 _25449_ (.A0(net5842),
    .A1(_01190_),
    .S(_11804_),
    .X(_11837_));
 sg13g2_nand2_1 _25450_ (.Y(_11838_),
    .A(_01189_),
    .B(net6250));
 sg13g2_o21ai_1 _25451_ (.B1(_11838_),
    .Y(_11839_),
    .A1(net5835),
    .A2(net5995));
 sg13g2_nand2_1 _25452_ (.Y(_11840_),
    .A(_01188_),
    .B(net6250));
 sg13g2_o21ai_1 _25453_ (.B1(_11840_),
    .Y(_11841_),
    .A1(net5901),
    .A2(net5995));
 sg13g2_nand2_1 _25454_ (.Y(_11842_),
    .A(_01187_),
    .B(net6250));
 sg13g2_mux2_1 _25455_ (.A0(_00996_),
    .A1(_01031_),
    .S(net7916),
    .X(_11843_));
 sg13g2_o21ai_1 _25456_ (.B1(_11842_),
    .Y(_11844_),
    .A1(net5896),
    .A2(_11804_));
 sg13g2_nand2_1 _25457_ (.Y(_11845_),
    .A(_01186_),
    .B(net6250));
 sg13g2_o21ai_1 _25458_ (.B1(_11845_),
    .Y(_11846_),
    .A1(net5893),
    .A2(net6250));
 sg13g2_nor3_1 _25459_ (.A(net7540),
    .B(net7524),
    .C(_11843_),
    .Y(_11847_));
 sg13g2_mux2_1 _25460_ (.A0(net5774),
    .A1(_01185_),
    .S(net6257),
    .X(_11848_));
 sg13g2_nand2_1 _25461_ (.Y(_11849_),
    .A(_01184_),
    .B(net6253));
 sg13g2_o21ai_1 _25462_ (.B1(_11849_),
    .Y(_11850_),
    .A1(net5883),
    .A2(net6253));
 sg13g2_nand2_1 _25463_ (.Y(_11851_),
    .A(_01183_),
    .B(net6256));
 sg13g2_o21ai_1 _25464_ (.B1(_11851_),
    .Y(_11852_),
    .A1(net5928),
    .A2(net6256));
 sg13g2_nand2_1 _25465_ (.Y(_11853_),
    .A(_01182_),
    .B(net6256));
 sg13g2_o21ai_1 _25466_ (.B1(_11853_),
    .Y(_11854_),
    .A1(net5965),
    .A2(net6256));
 sg13g2_nand2_1 _25467_ (.Y(_11855_),
    .A(_01181_),
    .B(net6264));
 sg13g2_o21ai_1 _25468_ (.B1(_11855_),
    .Y(_11856_),
    .A1(net5804),
    .A2(net6095));
 sg13g2_nand2_1 _25469_ (.Y(_11857_),
    .A(_01180_),
    .B(net6252));
 sg13g2_o21ai_1 _25470_ (.B1(_11857_),
    .Y(_11858_),
    .A1(_10857_),
    .A2(net6252));
 sg13g2_nand2_1 _25471_ (.Y(_11859_),
    .A(_01179_),
    .B(net6251));
 sg13g2_o21ai_1 _25472_ (.B1(_11859_),
    .Y(_11860_),
    .A1(net5960),
    .A2(_11804_));
 sg13g2_nand2_1 _25473_ (.Y(_11861_),
    .A(_01178_),
    .B(net6252));
 sg13g2_o21ai_1 _25474_ (.B1(_11861_),
    .Y(_11862_),
    .A1(net6008),
    .A2(net6252));
 sg13g2_nand2_1 _25475_ (.Y(_11863_),
    .A(_01177_),
    .B(net6254));
 sg13g2_o21ai_1 _25476_ (.B1(_11863_),
    .Y(_11864_),
    .A1(net6004),
    .A2(net6254));
 sg13g2_nand2_1 _25477_ (.Y(_11865_),
    .A(_01176_),
    .B(net6255));
 sg13g2_mux2_1 _25478_ (.A0(_00925_),
    .A1(_00960_),
    .S(net7916),
    .X(_11866_));
 sg13g2_o21ai_1 _25479_ (.B1(_11865_),
    .Y(_11867_),
    .A1(net6120),
    .A2(net6255));
 sg13g2_nand2_1 _25480_ (.Y(_11868_),
    .A(_01175_),
    .B(net6252));
 sg13g2_o21ai_1 _25481_ (.B1(_11868_),
    .Y(_11869_),
    .A1(net6029),
    .A2(net6252));
 sg13g2_nand2_1 _25482_ (.Y(_11870_),
    .A(_01174_),
    .B(net6255));
 sg13g2_nor3_1 _25483_ (.A(net7540),
    .B(_09028_),
    .C(_11866_),
    .Y(_11871_));
 sg13g2_o21ai_1 _25484_ (.B1(_11870_),
    .Y(_11872_),
    .A1(net6111),
    .A2(net6255));
 sg13g2_nand2_1 _25485_ (.Y(_11873_),
    .A(_01173_),
    .B(net6255));
 sg13g2_o21ai_1 _25486_ (.B1(_11873_),
    .Y(_11874_),
    .A1(net6028),
    .A2(net6255));
 sg13g2_nand2_1 _25487_ (.Y(_11875_),
    .A(_01172_),
    .B(net6253));
 sg13g2_o21ai_1 _25488_ (.B1(_11875_),
    .Y(_11876_),
    .A1(net6052),
    .A2(net6253));
 sg13g2_nand2_1 _25489_ (.Y(_11877_),
    .A(_01171_),
    .B(net6254));
 sg13g2_o21ai_1 _25490_ (.B1(_11877_),
    .Y(_11878_),
    .A1(net6019),
    .A2(net6254));
 sg13g2_nand2_1 _25491_ (.Y(_11879_),
    .A(_01170_),
    .B(net6260));
 sg13g2_o21ai_1 _25492_ (.B1(_11879_),
    .Y(_11880_),
    .A1(net5847),
    .A2(net6260));
 sg13g2_nand2_1 _25493_ (.Y(_11881_),
    .A(_01169_),
    .B(net6252));
 sg13g2_o21ai_1 _25494_ (.B1(_11881_),
    .Y(_11882_),
    .A1(net6106),
    .A2(net6252));
 sg13g2_nand2_1 _25495_ (.Y(_11883_),
    .A(_01168_),
    .B(net6251));
 sg13g2_o21ai_1 _25496_ (.B1(_11883_),
    .Y(_11884_),
    .A1(net5866),
    .A2(_11804_));
 sg13g2_nand4_1 _25497_ (.B(net7627),
    .C(net6466),
    .A(net7669),
    .Y(_11885_),
    .D(_10091_));
 sg13g2_nand2_1 _25498_ (.Y(_11886_),
    .A(_06619_),
    .B(_10094_));
 sg13g2_nand2_1 _25499_ (.Y(_11887_),
    .A(_01167_),
    .B(net6241));
 sg13g2_o21ai_1 _25500_ (.B1(_11887_),
    .Y(_11888_),
    .A1(net8286),
    .A2(net6241));
 sg13g2_nand2_1 _25501_ (.Y(_11889_),
    .A(_01166_),
    .B(net6247));
 sg13g2_nand2b_1 _25502_ (.Y(_11890_),
    .B(net6384),
    .A_N(net6247));
 sg13g2_o21ai_1 _25503_ (.B1(_11889_),
    .Y(_11891_),
    .A1(net5856),
    .A2(_11890_));
 sg13g2_nand2_1 _25504_ (.Y(_11892_),
    .A(_01165_),
    .B(net6249));
 sg13g2_o21ai_1 _25505_ (.B1(_11892_),
    .Y(_11893_),
    .A1(net5807),
    .A2(_11886_));
 sg13g2_nand2_1 _25506_ (.Y(_11894_),
    .A(_01164_),
    .B(net6247));
 sg13g2_o21ai_1 _25507_ (.B1(_11894_),
    .Y(_11895_),
    .A1(net5851),
    .A2(net6247));
 sg13g2_mux2_1 _25508_ (.A0(_01348_),
    .A1(_01383_),
    .S(net7915),
    .X(_11896_));
 sg13g2_nand2_1 _25509_ (.Y(_11897_),
    .A(_01163_),
    .B(net6245));
 sg13g2_o21ai_1 _25510_ (.B1(_11897_),
    .Y(_11898_),
    .A1(net5801),
    .A2(net6245));
 sg13g2_nand2_1 _25511_ (.Y(_11899_),
    .A(_01162_),
    .B(net6248));
 sg13g2_nor3_1 _25512_ (.A(_09152_),
    .B(net7470),
    .C(_11896_),
    .Y(_11900_));
 sg13g2_o21ai_1 _25513_ (.B1(_11899_),
    .Y(_11901_),
    .A1(net5796),
    .A2(net5994));
 sg13g2_nand2_1 _25514_ (.Y(_11902_),
    .A(_01161_),
    .B(net6244));
 sg13g2_nand2b_1 _25515_ (.Y(_11903_),
    .B(net6380),
    .A_N(net6244));
 sg13g2_o21ai_1 _25516_ (.B1(_11902_),
    .Y(_11904_),
    .A1(net5919),
    .A2(_11903_));
 sg13g2_nand2_1 _25517_ (.Y(_11905_),
    .A(_01160_),
    .B(net6248));
 sg13g2_o21ai_1 _25518_ (.B1(_11905_),
    .Y(_11906_),
    .A1(net5790),
    .A2(net5994));
 sg13g2_nand2_1 _25519_ (.Y(_11907_),
    .A(_01159_),
    .B(net6266));
 sg13g2_o21ai_1 _25520_ (.B1(_11907_),
    .Y(_11908_),
    .A1(net5803),
    .A2(net6266));
 sg13g2_nand2_1 _25521_ (.Y(_11909_),
    .A(_01158_),
    .B(net6241));
 sg13g2_nand2b_1 _25522_ (.Y(_11910_),
    .B(net6371),
    .A_N(net6241));
 sg13g2_o21ai_1 _25523_ (.B1(_11909_),
    .Y(_11911_),
    .A1(net5913),
    .A2(_11910_));
 sg13g2_nand2_1 _25524_ (.Y(_11912_),
    .A(_01157_),
    .B(net6248));
 sg13g2_o21ai_1 _25525_ (.B1(_11912_),
    .Y(_11913_),
    .A1(net5781),
    .A2(_11886_));
 sg13g2_nand2_1 _25526_ (.Y(_11914_),
    .A(_01156_),
    .B(net6241));
 sg13g2_nand2b_1 _25527_ (.Y(_11915_),
    .B(net6364),
    .A_N(net6241));
 sg13g2_o21ai_1 _25528_ (.B1(_11914_),
    .Y(_11916_),
    .A1(net5907),
    .A2(_11915_));
 sg13g2_mux2_1 _25529_ (.A0(net5842),
    .A1(_01155_),
    .S(_11886_),
    .X(_11917_));
 sg13g2_nand2_1 _25530_ (.Y(_11918_),
    .A(_01154_),
    .B(net6248));
 sg13g2_o21ai_1 _25531_ (.B1(_11918_),
    .Y(_11919_),
    .A1(net5835),
    .A2(net5994));
 sg13g2_nand2_1 _25532_ (.Y(_11920_),
    .A(_01153_),
    .B(net6248));
 sg13g2_mux2_1 _25533_ (.A0(_01418_),
    .A1(_01453_),
    .S(net7915),
    .X(_11921_));
 sg13g2_o21ai_1 _25534_ (.B1(_11920_),
    .Y(_11922_),
    .A1(net5901),
    .A2(_11886_));
 sg13g2_nand2_1 _25535_ (.Y(_11923_),
    .A(_01152_),
    .B(net6248));
 sg13g2_nor3_1 _25536_ (.A(_09152_),
    .B(net7460),
    .C(_11921_),
    .Y(_11924_));
 sg13g2_o21ai_1 _25537_ (.B1(_11923_),
    .Y(_11925_),
    .A1(net5896),
    .A2(_11886_));
 sg13g2_nand2_1 _25538_ (.Y(_11926_),
    .A(_01151_),
    .B(net6248));
 sg13g2_o21ai_1 _25539_ (.B1(_11926_),
    .Y(_11927_),
    .A1(net5893),
    .A2(net6248));
 sg13g2_mux2_1 _25540_ (.A0(net5774),
    .A1(_01150_),
    .S(net6241),
    .X(_11928_));
 sg13g2_nand2_1 _25541_ (.Y(_11929_),
    .A(_01149_),
    .B(net6242));
 sg13g2_o21ai_1 _25542_ (.B1(_11929_),
    .Y(_11930_),
    .A1(net5883),
    .A2(net6242));
 sg13g2_nand2_1 _25543_ (.Y(_11931_),
    .A(_01148_),
    .B(net6264));
 sg13g2_nor4_1 _25544_ (.A(_11847_),
    .B(_11871_),
    .C(_11900_),
    .D(_11924_),
    .Y(_11932_));
 sg13g2_o21ai_1 _25545_ (.B1(_11931_),
    .Y(_11933_),
    .A1(net5792),
    .A2(_11800_));
 sg13g2_nand2_1 _25546_ (.Y(_11934_),
    .A(_01147_),
    .B(net6246));
 sg13g2_o21ai_1 _25547_ (.B1(_11934_),
    .Y(_11935_),
    .A1(net5927),
    .A2(net6246));
 sg13g2_nand2_1 _25548_ (.Y(_11936_),
    .A(_01146_),
    .B(net6245));
 sg13g2_o21ai_1 _25549_ (.B1(_11936_),
    .Y(_11937_),
    .A1(net5965),
    .A2(net6245));
 sg13g2_nand2_1 _25550_ (.Y(_11938_),
    .A(_01145_),
    .B(net6243));
 sg13g2_o21ai_1 _25551_ (.B1(_11938_),
    .Y(_11939_),
    .A1(net6012),
    .A2(net6243));
 sg13g2_nand2_1 _25552_ (.Y(_11940_),
    .A(_01144_),
    .B(net6249));
 sg13g2_o21ai_1 _25553_ (.B1(_11940_),
    .Y(_11941_),
    .A1(net5960),
    .A2(_11886_));
 sg13g2_nand2_1 _25554_ (.Y(_11942_),
    .A(_01143_),
    .B(net6243));
 sg13g2_o21ai_1 _25555_ (.B1(_11942_),
    .Y(_11943_),
    .A1(net6008),
    .A2(net6243));
 sg13g2_nand2_1 _25556_ (.Y(_11944_),
    .A(_01142_),
    .B(net6242));
 sg13g2_o21ai_1 _25557_ (.B1(_11944_),
    .Y(_11945_),
    .A1(net6003),
    .A2(net6242));
 sg13g2_nand2_1 _25558_ (.Y(_11946_),
    .A(_01141_),
    .B(net6246));
 sg13g2_o21ai_1 _25559_ (.B1(_11946_),
    .Y(_11947_),
    .A1(net6120),
    .A2(net6246));
 sg13g2_nand2_1 _25560_ (.Y(_11948_),
    .A(_01140_),
    .B(net6243));
 sg13g2_o21ai_1 _25561_ (.B1(_11948_),
    .Y(_11949_),
    .A1(net6029),
    .A2(net6243));
 sg13g2_nand2_1 _25562_ (.Y(_11950_),
    .A(_01139_),
    .B(net6247));
 sg13g2_o21ai_1 _25563_ (.B1(_11950_),
    .Y(_11951_),
    .A1(net6111),
    .A2(net6247));
 sg13g2_nand2_1 _25564_ (.Y(_11952_),
    .A(_01138_),
    .B(net6246));
 sg13g2_o21ai_1 _25565_ (.B1(_11952_),
    .Y(_11953_),
    .A1(net6028),
    .A2(net6246));
 sg13g2_nand2_1 _25566_ (.Y(_11954_),
    .A(_01137_),
    .B(net6267));
 sg13g2_nand2b_1 _25567_ (.Y(_11955_),
    .B(net6379),
    .A_N(net6267));
 sg13g2_o21ai_1 _25568_ (.B1(_11954_),
    .Y(_11956_),
    .A1(net5918),
    .A2(_11955_));
 sg13g2_nand2_1 _25569_ (.Y(_11957_),
    .A(_01136_),
    .B(net6242));
 sg13g2_o21ai_1 _25570_ (.B1(_11957_),
    .Y(_11958_),
    .A1(net6052),
    .A2(net6242));
 sg13g2_nand2_1 _25571_ (.Y(_11959_),
    .A(_01135_),
    .B(net6244));
 sg13g2_o21ai_1 _25572_ (.B1(_11959_),
    .Y(_11960_),
    .A1(net6019),
    .A2(net6244));
 sg13g2_nand2_1 _25573_ (.Y(_11961_),
    .A(_01134_),
    .B(net6243));
 sg13g2_o21ai_1 _25574_ (.B1(_11961_),
    .Y(_11962_),
    .A1(net6105),
    .A2(net6243));
 sg13g2_nand2_1 _25575_ (.Y(_11963_),
    .A(_01133_),
    .B(net6249));
 sg13g2_o21ai_1 _25576_ (.B1(_11963_),
    .Y(_11964_),
    .A1(net5866),
    .A2(_11886_));
 sg13g2_or4_1 _25577_ (.A(net7667),
    .B(_06620_),
    .C(net6468),
    .D(_09682_),
    .X(_11965_));
 sg13g2_nand2_1 _25578_ (.Y(_11966_),
    .A(_06619_),
    .B(net6346));
 sg13g2_nand2_1 _25579_ (.Y(_11967_),
    .A(_01132_),
    .B(net6235));
 sg13g2_o21ai_1 _25580_ (.B1(_11967_),
    .Y(_11968_),
    .A1(net5860),
    .A2(net6235));
 sg13g2_nand2_1 _25581_ (.Y(_11969_),
    .A(_01131_),
    .B(net6240));
 sg13g2_nand2b_1 _25582_ (.Y(_11970_),
    .B(net6384),
    .A_N(_11965_));
 sg13g2_o21ai_1 _25583_ (.B1(_11969_),
    .Y(_11971_),
    .A1(net5856),
    .A2(_11970_));
 sg13g2_nand2_1 _25584_ (.Y(_11972_),
    .A(_01130_),
    .B(net6234));
 sg13g2_o21ai_1 _25585_ (.B1(_11972_),
    .Y(_11973_),
    .A1(net5807),
    .A2(net6093));
 sg13g2_nand2_1 _25586_ (.Y(_11974_),
    .A(_01129_),
    .B(net6239));
 sg13g2_mux2_1 _25587_ (.A0(_01247_),
    .A1(_01599_),
    .S(net7858),
    .X(_11975_));
 sg13g2_o21ai_1 _25588_ (.B1(_11974_),
    .Y(_11976_),
    .A1(net5851),
    .A2(net6239));
 sg13g2_nand2_1 _25589_ (.Y(_11977_),
    .A(_01128_),
    .B(net6240));
 sg13g2_o21ai_1 _25590_ (.B1(_11977_),
    .Y(_11978_),
    .A1(net5801),
    .A2(net6240));
 sg13g2_nand2_1 _25591_ (.Y(_11979_),
    .A(_01127_),
    .B(net6233));
 sg13g2_o21ai_1 _25592_ (.B1(_11979_),
    .Y(_11980_),
    .A1(net5796),
    .A2(net6094));
 sg13g2_nand2_1 _25593_ (.Y(_11981_),
    .A(_01126_),
    .B(net6263));
 sg13g2_o21ai_1 _25594_ (.B1(_11981_),
    .Y(_11982_),
    .A1(net5786),
    .A2(net6095));
 sg13g2_nand2_1 _25595_ (.Y(_11983_),
    .A(_01125_),
    .B(net6238));
 sg13g2_nand2b_1 _25596_ (.Y(_11984_),
    .B(net6380),
    .A_N(net6238));
 sg13g2_o21ai_1 _25597_ (.B1(_11983_),
    .Y(_11985_),
    .A1(net5919),
    .A2(_11984_));
 sg13g2_nand2_1 _25598_ (.Y(_11986_),
    .A(_01124_),
    .B(net6233));
 sg13g2_o21ai_1 _25599_ (.B1(_11986_),
    .Y(_11987_),
    .A1(net5790),
    .A2(net6094));
 sg13g2_nand2_1 _25600_ (.Y(_11988_),
    .A(_01123_),
    .B(net6235));
 sg13g2_nand2b_1 _25601_ (.Y(_11989_),
    .B(net6371),
    .A_N(net6235));
 sg13g2_o21ai_1 _25602_ (.B1(_11988_),
    .Y(_11990_),
    .A1(net5913),
    .A2(_11989_));
 sg13g2_nand2_1 _25603_ (.Y(_11991_),
    .A(_01122_),
    .B(net6234));
 sg13g2_o21ai_1 _25604_ (.B1(_11991_),
    .Y(_11992_),
    .A1(net5781),
    .A2(net6093));
 sg13g2_nand2_1 _25605_ (.Y(_11993_),
    .A(_01121_),
    .B(net6235));
 sg13g2_nand2b_1 _25606_ (.Y(_11994_),
    .B(net6364),
    .A_N(net6235));
 sg13g2_o21ai_1 _25607_ (.B1(_11993_),
    .Y(_11995_),
    .A1(net5907),
    .A2(_11994_));
 sg13g2_mux2_1 _25608_ (.A0(net5842),
    .A1(_01120_),
    .S(net6093),
    .X(_11996_));
 sg13g2_nand2_1 _25609_ (.Y(_11997_),
    .A(_01119_),
    .B(net6233));
 sg13g2_o21ai_1 _25610_ (.B1(_11997_),
    .Y(_11998_),
    .A1(net5835),
    .A2(net6094));
 sg13g2_nand2_1 _25611_ (.Y(_11999_),
    .A(_01118_),
    .B(net6233));
 sg13g2_o21ai_1 _25612_ (.B1(_11999_),
    .Y(_12000_),
    .A1(net5901),
    .A2(net6094));
 sg13g2_nand2_1 _25613_ (.Y(_12001_),
    .A(_01117_),
    .B(net6234));
 sg13g2_o21ai_1 _25614_ (.B1(_12001_),
    .Y(_12002_),
    .A1(net5896),
    .A2(net6093));
 sg13g2_nand2_1 _25615_ (.Y(_12003_),
    .A(_01116_),
    .B(net6233));
 sg13g2_o21ai_1 _25616_ (.B1(_12003_),
    .Y(_12004_),
    .A1(net5893),
    .A2(net6233));
 sg13g2_nand2b_1 _25617_ (.Y(_12005_),
    .B(net6370),
    .A_N(_11798_));
 sg13g2_nand2_1 _25618_ (.Y(_12006_),
    .A(_01115_),
    .B(_11798_));
 sg13g2_o21ai_1 _25619_ (.B1(_12006_),
    .Y(_12007_),
    .A1(net5915),
    .A2(_12005_));
 sg13g2_mux2_1 _25620_ (.A0(net5774),
    .A1(_01114_),
    .S(net6235),
    .X(_12008_));
 sg13g2_nand2_1 _25621_ (.Y(_12009_),
    .A(_01113_),
    .B(net6237));
 sg13g2_o21ai_1 _25622_ (.B1(_12009_),
    .Y(_12010_),
    .A1(net5883),
    .A2(net6237));
 sg13g2_nand2_1 _25623_ (.Y(_12011_),
    .A(_01112_),
    .B(net6240));
 sg13g2_o21ai_1 _25624_ (.B1(_12011_),
    .Y(_12012_),
    .A1(net5928),
    .A2(net6240));
 sg13g2_nand2_1 _25625_ (.Y(_12013_),
    .A(_01111_),
    .B(net6240));
 sg13g2_o21ai_1 _25626_ (.B1(_12013_),
    .Y(_12014_),
    .A1(net5965),
    .A2(net6240));
 sg13g2_nand2_1 _25627_ (.Y(_12015_),
    .A(_01110_),
    .B(net6236));
 sg13g2_o21ai_1 _25628_ (.B1(_12015_),
    .Y(_12016_),
    .A1(net6012),
    .A2(net6236));
 sg13g2_nand2_1 _25629_ (.Y(_12017_),
    .A(_01109_),
    .B(net6234));
 sg13g2_o21ai_1 _25630_ (.B1(_12017_),
    .Y(_12018_),
    .A1(net5960),
    .A2(net6093));
 sg13g2_nand2_1 _25631_ (.Y(_12019_),
    .A(_01108_),
    .B(net6236));
 sg13g2_o21ai_1 _25632_ (.B1(_12019_),
    .Y(_12020_),
    .A1(net6008),
    .A2(net6236));
 sg13g2_nand2_1 _25633_ (.Y(_12021_),
    .A(_01107_),
    .B(net6238));
 sg13g2_o21ai_1 _25634_ (.B1(_12021_),
    .Y(_12022_),
    .A1(net6004),
    .A2(net6238));
 sg13g2_nand2_1 _25635_ (.Y(_12023_),
    .A(_01106_),
    .B(net6239));
 sg13g2_mux4_1 _25636_ (.S0(net7858),
    .A0(_00663_),
    .A1(_00695_),
    .A2(_00727_),
    .A3(_00759_),
    .S1(net7832),
    .X(_12024_));
 sg13g2_o21ai_1 _25637_ (.B1(_12023_),
    .Y(_12025_),
    .A1(net6120),
    .A2(net6239));
 sg13g2_nand2_1 _25638_ (.Y(_12026_),
    .A(_01105_),
    .B(net6236));
 sg13g2_o21ai_1 _25639_ (.B1(_12026_),
    .Y(_12027_),
    .A1(net6029),
    .A2(net6236));
 sg13g2_nand2_1 _25640_ (.Y(_12028_),
    .A(_01104_),
    .B(net6264));
 sg13g2_o21ai_1 _25641_ (.B1(_12028_),
    .Y(_12029_),
    .A1(net5783),
    .A2(net6095));
 sg13g2_nand2_1 _25642_ (.Y(_12030_),
    .A(_01103_),
    .B(net6239));
 sg13g2_o21ai_1 _25643_ (.B1(_12030_),
    .Y(_12031_),
    .A1(net6111),
    .A2(net6239));
 sg13g2_nand2_1 _25644_ (.Y(_12032_),
    .A(_01102_),
    .B(net6239));
 sg13g2_o21ai_1 _25645_ (.B1(_12032_),
    .Y(_12033_),
    .A1(net6025),
    .A2(net6239));
 sg13g2_nand2_1 _25646_ (.Y(_12034_),
    .A(_01101_),
    .B(net6237));
 sg13g2_o21ai_1 _25647_ (.B1(_12034_),
    .Y(_12035_),
    .A1(net6052),
    .A2(net6237));
 sg13g2_nand2_1 _25648_ (.Y(_12036_),
    .A(_01100_),
    .B(net6238));
 sg13g2_o21ai_1 _25649_ (.B1(_12036_),
    .Y(_12037_),
    .A1(net6019),
    .A2(net6238));
 sg13g2_nand2_1 _25650_ (.Y(_12038_),
    .A(_01099_),
    .B(net6236));
 sg13g2_o21ai_1 _25651_ (.B1(_12038_),
    .Y(_12039_),
    .A1(net6105),
    .A2(net6236));
 sg13g2_nand2_1 _25652_ (.Y(_12040_),
    .A(_01098_),
    .B(net6234));
 sg13g2_o21ai_1 _25653_ (.B1(_12040_),
    .Y(_12041_),
    .A1(net5866),
    .A2(net6093));
 sg13g2_nand2_2 _25654_ (.Y(_12042_),
    .A(net7627),
    .B(_11075_));
 sg13g2_nand2_1 _25655_ (.Y(_12043_),
    .A(_01097_),
    .B(net6086));
 sg13g2_nor2_1 _25656_ (.A(net7484),
    .B(_12024_),
    .Y(_12044_));
 sg13g2_o21ai_1 _25657_ (.B1(_12043_),
    .Y(_12045_),
    .A1(net5860),
    .A2(net6086));
 sg13g2_nand3_1 _25658_ (.B(_10162_),
    .C(net6336),
    .A(net7627),
    .Y(_12046_));
 sg13g2_nand2_1 _25659_ (.Y(_12047_),
    .A(_01096_),
    .B(net6092));
 sg13g2_o21ai_1 _25660_ (.B1(_12047_),
    .Y(_12048_),
    .A1(net5854),
    .A2(_12046_));
 sg13g2_nand2_1 _25661_ (.Y(_12049_),
    .A(_01095_),
    .B(net6083));
 sg13g2_o21ai_1 _25662_ (.B1(_12049_),
    .Y(_12050_),
    .A1(net5807),
    .A2(net6083));
 sg13g2_nand2_1 _25663_ (.Y(_12051_),
    .A(_01094_),
    .B(net6091));
 sg13g2_o21ai_1 _25664_ (.B1(_12051_),
    .Y(_12052_),
    .A1(net5849),
    .A2(net6091));
 sg13g2_nand2b_1 _25665_ (.Y(_12053_),
    .B(net6365),
    .A_N(_11798_));
 sg13g2_nand2_1 _25666_ (.Y(_12054_),
    .A(_01093_),
    .B(_11798_));
 sg13g2_o21ai_1 _25667_ (.B1(_12054_),
    .Y(_12055_),
    .A1(net5908),
    .A2(_12053_));
 sg13g2_nand2_1 _25668_ (.Y(_12056_),
    .A(_01092_),
    .B(net6090));
 sg13g2_o21ai_1 _25669_ (.B1(_12056_),
    .Y(_12057_),
    .A1(net5801),
    .A2(net6090));
 sg13g2_nand2_1 _25670_ (.Y(_12058_),
    .A(_01091_),
    .B(net6084));
 sg13g2_o21ai_1 _25671_ (.B1(_12058_),
    .Y(_12059_),
    .A1(net5796),
    .A2(net6084));
 sg13g2_nand3_1 _25672_ (.B(_10341_),
    .C(net6336),
    .A(net7627),
    .Y(_12060_));
 sg13g2_a221oi_1 _25673_ (.B2(net7835),
    .C1(_01894_),
    .B1(_11975_),
    .A1(_00895_),
    .Y(_12061_),
    .A2(_08988_));
 sg13g2_nand2_1 _25674_ (.Y(_12062_),
    .A(_01090_),
    .B(net6086));
 sg13g2_o21ai_1 _25675_ (.B1(_12062_),
    .Y(_12063_),
    .A1(net5920),
    .A2(_12060_));
 sg13g2_nand2_1 _25676_ (.Y(_12064_),
    .A(_01089_),
    .B(net6085));
 sg13g2_o21ai_1 _25677_ (.B1(_12064_),
    .Y(_12065_),
    .A1(net5790),
    .A2(net6085));
 sg13g2_nand3_1 _25678_ (.B(_10415_),
    .C(net6336),
    .A(net7627),
    .Y(_12066_));
 sg13g2_nand2_1 _25679_ (.Y(_12067_),
    .A(_01088_),
    .B(net6086));
 sg13g2_o21ai_1 _25680_ (.B1(_12067_),
    .Y(_12068_),
    .A1(net5916),
    .A2(_12066_));
 sg13g2_nand2_1 _25681_ (.Y(_12069_),
    .A(_01087_),
    .B(net6083));
 sg13g2_o21ai_1 _25682_ (.B1(_12069_),
    .Y(_12070_),
    .A1(net5781),
    .A2(net6083));
 sg13g2_nand3_1 _25683_ (.B(net6367),
    .C(net6336),
    .A(net7627),
    .Y(_12071_));
 sg13g2_nand2_1 _25684_ (.Y(_12072_),
    .A(_01086_),
    .B(net6086));
 sg13g2_o21ai_1 _25685_ (.B1(_12072_),
    .Y(_12073_),
    .A1(net5909),
    .A2(_12071_));
 sg13g2_o21ai_1 _25686_ (.B1(_08973_),
    .Y(_12074_),
    .A1(_12044_),
    .A2(_12061_));
 sg13g2_mux2_1 _25687_ (.A0(net5842),
    .A1(_01085_),
    .S(_12042_),
    .X(_12075_));
 sg13g2_nand2_1 _25688_ (.Y(_12076_),
    .A(_01084_),
    .B(net6084));
 sg13g2_o21ai_1 _25689_ (.B1(_12076_),
    .Y(_12077_),
    .A1(net5835),
    .A2(net6084));
 sg13g2_nand2_1 _25690_ (.Y(_12078_),
    .A(_01083_),
    .B(net6085));
 sg13g2_o21ai_1 _25691_ (.B1(_12078_),
    .Y(_12079_),
    .A1(net5901),
    .A2(net6085));
 sg13g2_mux2_1 _25692_ (.A0(net5838),
    .A1(_01082_),
    .S(net6095),
    .X(_12080_));
 sg13g2_nand2_1 _25693_ (.Y(_12081_),
    .A(_01081_),
    .B(net6085));
 sg13g2_o21ai_1 _25694_ (.B1(_12081_),
    .Y(_12082_),
    .A1(net5896),
    .A2(net6085));
 sg13g2_nand2_1 _25695_ (.Y(_12083_),
    .A(_01080_),
    .B(net6084));
 sg13g2_o21ai_1 _25696_ (.B1(_12083_),
    .Y(_12084_),
    .A1(net5893),
    .A2(net6084));
 sg13g2_mux2_1 _25697_ (.A0(net5774),
    .A1(_01079_),
    .S(net6086),
    .X(_12085_));
 sg13g2_nand2_1 _25698_ (.Y(_12086_),
    .A(_01078_),
    .B(net6088));
 sg13g2_o21ai_1 _25699_ (.B1(_12086_),
    .Y(_12087_),
    .A1(net5883),
    .A2(net6088));
 sg13g2_nand2_1 _25700_ (.Y(_12088_),
    .A(_01077_),
    .B(net6090));
 sg13g2_o21ai_1 _25701_ (.B1(_12088_),
    .Y(_12089_),
    .A1(net5928),
    .A2(net6090));
 sg13g2_nand2_1 _25702_ (.Y(_12090_),
    .A(_01076_),
    .B(net6090));
 sg13g2_o21ai_1 _25703_ (.B1(_12090_),
    .Y(_12091_),
    .A1(net5965),
    .A2(net6090));
 sg13g2_nand2_1 _25704_ (.Y(_12092_),
    .A(_01075_),
    .B(net6089));
 sg13g2_o21ai_1 _25705_ (.B1(_12092_),
    .Y(_12093_),
    .A1(net6012),
    .A2(net6089));
 sg13g2_nand2_1 _25706_ (.Y(_12094_),
    .A(_01074_),
    .B(net6083));
 sg13g2_o21ai_1 _25707_ (.B1(_12094_),
    .Y(_12095_),
    .A1(net5960),
    .A2(net6083));
 sg13g2_nand2_1 _25708_ (.Y(_12096_),
    .A(_01073_),
    .B(net6089));
 sg13g2_o21ai_1 _25709_ (.B1(_12096_),
    .Y(_12097_),
    .A1(net6008),
    .A2(net6089));
 sg13g2_nand2_1 _25710_ (.Y(_12098_),
    .A(_01072_),
    .B(net6087));
 sg13g2_o21ai_1 _25711_ (.B1(_12098_),
    .Y(_12099_),
    .A1(net6004),
    .A2(net6087));
 sg13g2_nand2_1 _25712_ (.Y(_12100_),
    .A(_01071_),
    .B(net6263));
 sg13g2_o21ai_1 _25713_ (.B1(_12100_),
    .Y(_12101_),
    .A1(net5836),
    .A2(_11800_));
 sg13g2_nand2_1 _25714_ (.Y(_12102_),
    .A(_01070_),
    .B(net6091));
 sg13g2_o21ai_1 _25715_ (.B1(_12102_),
    .Y(_12103_),
    .A1(net6120),
    .A2(net6091));
 sg13g2_nand2_1 _25716_ (.Y(_12104_),
    .A(_01069_),
    .B(net6089));
 sg13g2_o21ai_1 _25717_ (.B1(_12104_),
    .Y(_12105_),
    .A1(net6029),
    .A2(net6089));
 sg13g2_nand2_1 _25718_ (.Y(_12106_),
    .A(_01068_),
    .B(net6092));
 sg13g2_o21ai_1 _25719_ (.B1(_12106_),
    .Y(_12107_),
    .A1(net6111),
    .A2(net6092));
 sg13g2_nand2_1 _25720_ (.Y(_12108_),
    .A(_01067_),
    .B(net6091));
 sg13g2_o21ai_1 _25721_ (.B1(_12108_),
    .Y(_12109_),
    .A1(net6025),
    .A2(net6091));
 sg13g2_nand2_1 _25722_ (.Y(_12110_),
    .A(_01066_),
    .B(net6088));
 sg13g2_o21ai_1 _25723_ (.B1(_12110_),
    .Y(_12111_),
    .A1(net6052),
    .A2(net6088));
 sg13g2_nand2_1 _25724_ (.Y(_12112_),
    .A(_01065_),
    .B(net6087));
 sg13g2_o21ai_1 _25725_ (.B1(_12112_),
    .Y(_12113_),
    .A1(net6019),
    .A2(net6087));
 sg13g2_nand2_1 _25726_ (.Y(_12114_),
    .A(_01064_),
    .B(net6089));
 sg13g2_o21ai_1 _25727_ (.B1(_12114_),
    .Y(_12115_),
    .A1(net6105),
    .A2(net6089));
 sg13g2_nand2_1 _25728_ (.Y(_12116_),
    .A(_01063_),
    .B(net6083));
 sg13g2_o21ai_1 _25729_ (.B1(_12116_),
    .Y(_12117_),
    .A1(net5866),
    .A2(net6083));
 sg13g2_nand4_1 _25730_ (.B(_09604_),
    .C(_09605_),
    .A(net7668),
    .Y(_12118_),
    .D(net7474));
 sg13g2_nand2_1 _25731_ (.Y(_12119_),
    .A(_09608_),
    .B(net7474));
 sg13g2_nand2_1 _25732_ (.Y(_12120_),
    .A(_01062_),
    .B(net6231));
 sg13g2_o21ai_1 _25733_ (.B1(_12120_),
    .Y(_12121_),
    .A1(net5862),
    .A2(net6231));
 sg13g2_nand2_1 _25734_ (.Y(_12122_),
    .A(_01061_),
    .B(net6231));
 sg13g2_nand2b_1 _25735_ (.Y(_12123_),
    .B(net6381),
    .A_N(net6231));
 sg13g2_o21ai_1 _25736_ (.B1(_12122_),
    .Y(_12124_),
    .A1(net5855),
    .A2(_12123_));
 sg13g2_nand2_1 _25737_ (.Y(_12125_),
    .A(_01060_),
    .B(net6264));
 sg13g2_o21ai_1 _25738_ (.B1(_12125_),
    .Y(_12126_),
    .A1(net5902),
    .A2(net6095));
 sg13g2_nand2_1 _25739_ (.Y(_12127_),
    .A(_01059_),
    .B(net6225));
 sg13g2_o21ai_1 _25740_ (.B1(_12127_),
    .Y(_12128_),
    .A1(net5806),
    .A2(net5993));
 sg13g2_nand2_1 _25741_ (.Y(_12129_),
    .A(_01058_),
    .B(net6229));
 sg13g2_o21ai_1 _25742_ (.B1(_12129_),
    .Y(_12130_),
    .A1(net5847),
    .A2(net6229));
 sg13g2_nand2_1 _25743_ (.Y(_12131_),
    .A(_01057_),
    .B(net6230));
 sg13g2_mux4_1 _25744_ (.S0(net7915),
    .A0(_01066_),
    .A1(_01101_),
    .A2(_01136_),
    .A3(_01172_),
    .S1(net7828),
    .X(_12132_));
 sg13g2_o21ai_1 _25745_ (.B1(_12131_),
    .Y(_12133_),
    .A1(net5798),
    .A2(net6230));
 sg13g2_nand2_1 _25746_ (.Y(_12134_),
    .A(_01056_),
    .B(net6225));
 sg13g2_nor2_1 _25747_ (.A(net7814),
    .B(net7500),
    .Y(_12135_));
 sg13g2_o21ai_1 _25748_ (.B1(_12134_),
    .Y(_12136_),
    .A1(net5797),
    .A2(_12119_));
 sg13g2_nand2_1 _25749_ (.Y(_12137_),
    .A(_01055_),
    .B(net6231));
 sg13g2_nand2b_1 _25750_ (.Y(_12138_),
    .B(net6377),
    .A_N(net6231));
 sg13g2_nand2_1 _25751_ (.Y(_12139_),
    .A(net7485),
    .B(_09070_));
 sg13g2_o21ai_1 _25752_ (.B1(_12137_),
    .Y(_12140_),
    .A1(net5920),
    .A2(_12138_));
 sg13g2_nand2_1 _25753_ (.Y(_12141_),
    .A(_01054_),
    .B(net6225));
 sg13g2_nor3_1 _25754_ (.A(net7814),
    .B(net7500),
    .C(_12132_),
    .Y(_12142_));
 sg13g2_o21ai_1 _25755_ (.B1(_12141_),
    .Y(_12143_),
    .A1(net5788),
    .A2(_12119_));
 sg13g2_nand2_1 _25756_ (.Y(_12144_),
    .A(_01053_),
    .B(net6232));
 sg13g2_nand2b_1 _25757_ (.Y(_12145_),
    .B(net6376),
    .A_N(net6232));
 sg13g2_o21ai_1 _25758_ (.B1(_12144_),
    .Y(_12146_),
    .A1(net5916),
    .A2(_12145_));
 sg13g2_nand2_1 _25759_ (.Y(_12147_),
    .A(_01052_),
    .B(net6225));
 sg13g2_o21ai_1 _25760_ (.B1(_12147_),
    .Y(_12148_),
    .A1(net5780),
    .A2(net5993));
 sg13g2_nand2_1 _25761_ (.Y(_12149_),
    .A(_01051_),
    .B(net6232));
 sg13g2_nand2b_1 _25762_ (.Y(_12150_),
    .B(net6367),
    .A_N(net6232));
 sg13g2_o21ai_1 _25763_ (.B1(_12149_),
    .Y(_12151_),
    .A1(net5909),
    .A2(_12150_));
 sg13g2_mux2_1 _25764_ (.A0(net5841),
    .A1(_01050_),
    .S(net5993),
    .X(_12152_));
 sg13g2_nand2_1 _25765_ (.Y(_12153_),
    .A(_01049_),
    .B(net6264));
 sg13g2_o21ai_1 _25766_ (.B1(_12153_),
    .Y(_12154_),
    .A1(net5897),
    .A2(net6095));
 sg13g2_nand2_1 _25767_ (.Y(_12155_),
    .A(_01048_),
    .B(net6228));
 sg13g2_o21ai_1 _25768_ (.B1(_12155_),
    .Y(_12156_),
    .A1(net5834),
    .A2(_12119_));
 sg13g2_nand2_1 _25769_ (.Y(_12157_),
    .A(_01047_),
    .B(net6225));
 sg13g2_o21ai_1 _25770_ (.B1(_12157_),
    .Y(_12158_),
    .A1(net5904),
    .A2(_12119_));
 sg13g2_nand2_1 _25771_ (.Y(_12159_),
    .A(_01046_),
    .B(net6225));
 sg13g2_o21ai_1 _25772_ (.B1(_12159_),
    .Y(_12160_),
    .A1(net5898),
    .A2(net5993));
 sg13g2_nand2_1 _25773_ (.Y(_12161_),
    .A(_01045_),
    .B(net6228));
 sg13g2_o21ai_1 _25774_ (.B1(_12161_),
    .Y(_12162_),
    .A1(net5890),
    .A2(net6228));
 sg13g2_mux2_1 _25775_ (.A0(net5773),
    .A1(_01044_),
    .S(net6232),
    .X(_12163_));
 sg13g2_nand2_1 _25776_ (.Y(_12164_),
    .A(_01043_),
    .B(net6228));
 sg13g2_o21ai_1 _25777_ (.B1(_12164_),
    .Y(_12165_),
    .A1(net5882),
    .A2(net6228));
 sg13g2_nand2_1 _25778_ (.Y(_12166_),
    .A(_01042_),
    .B(net6230));
 sg13g2_o21ai_1 _25779_ (.B1(_12166_),
    .Y(_12167_),
    .A1(net5926),
    .A2(net6230));
 sg13g2_nand2_1 _25780_ (.Y(_12168_),
    .A(_01041_),
    .B(net6230));
 sg13g2_o21ai_1 _25781_ (.B1(_12168_),
    .Y(_12169_),
    .A1(net5963),
    .A2(net6230));
 sg13g2_nand2_1 _25782_ (.Y(_12170_),
    .A(_01040_),
    .B(net6226));
 sg13g2_o21ai_1 _25783_ (.B1(_12170_),
    .Y(_12171_),
    .A1(net6015),
    .A2(net6226));
 sg13g2_nand2_1 _25784_ (.Y(_12172_),
    .A(_01039_),
    .B(net6225));
 sg13g2_o21ai_1 _25785_ (.B1(_12172_),
    .Y(_12173_),
    .A1(net5961),
    .A2(net5993));
 sg13g2_nand2_1 _25786_ (.Y(_12174_),
    .A(_01038_),
    .B(net6263));
 sg13g2_o21ai_1 _25787_ (.B1(_12174_),
    .Y(_12175_),
    .A1(net5888),
    .A2(net6263));
 sg13g2_nand2_1 _25788_ (.Y(_12176_),
    .A(_01037_),
    .B(net6226));
 sg13g2_o21ai_1 _25789_ (.B1(_12176_),
    .Y(_12177_),
    .A1(net6011),
    .A2(net6226));
 sg13g2_nand2_1 _25790_ (.Y(_12178_),
    .A(_01036_),
    .B(net6226));
 sg13g2_o21ai_1 _25791_ (.B1(_12178_),
    .Y(_12179_),
    .A1(net6005),
    .A2(net6226));
 sg13g2_nand2_1 _25792_ (.Y(_12180_),
    .A(_01035_),
    .B(net6229));
 sg13g2_mux4_1 _25793_ (.S0(net7915),
    .A0(_01207_),
    .A1(_01242_),
    .A2(_01277_),
    .A3(_01312_),
    .S1(net7828),
    .X(_12181_));
 sg13g2_o21ai_1 _25794_ (.B1(_12180_),
    .Y(_12182_),
    .A1(net6117),
    .A2(net6229));
 sg13g2_nand2_1 _25795_ (.Y(_12183_),
    .A(_01034_),
    .B(net6230));
 sg13g2_o21ai_1 _25796_ (.B1(_12183_),
    .Y(_12184_),
    .A1(net6032),
    .A2(net6230));
 sg13g2_nand2_1 _25797_ (.Y(_12185_),
    .A(_01033_),
    .B(net6229));
 sg13g2_o21ai_1 _25798_ (.B1(_12185_),
    .Y(_12186_),
    .A1(net6112),
    .A2(net6229));
 sg13g2_nand3b_1 _25799_ (.B(net7813),
    .C(net7806),
    .Y(_12187_),
    .A_N(net7808));
 sg13g2_nand2_1 _25800_ (.Y(_12188_),
    .A(_01032_),
    .B(net6229));
 sg13g2_o21ai_1 _25801_ (.B1(_12188_),
    .Y(_12189_),
    .A1(net6023),
    .A2(net6229));
 sg13g2_nor2_1 _25802_ (.A(_12181_),
    .B(net7445),
    .Y(_12190_));
 sg13g2_nand2_1 _25803_ (.Y(_12191_),
    .A(_01031_),
    .B(net6227));
 sg13g2_o21ai_1 _25804_ (.B1(_12191_),
    .Y(_12192_),
    .A1(net6054),
    .A2(net6228));
 sg13g2_nand2_1 _25805_ (.Y(_12193_),
    .A(_01030_),
    .B(net6226));
 sg13g2_o21ai_1 _25806_ (.B1(_12193_),
    .Y(_12194_),
    .A1(net6021),
    .A2(net6226));
 sg13g2_nand2_1 _25807_ (.Y(_12195_),
    .A(_01029_),
    .B(net6227));
 sg13g2_o21ai_1 _25808_ (.B1(_12195_),
    .Y(_12196_),
    .A1(net6107),
    .A2(net6227));
 sg13g2_nand2_1 _25809_ (.Y(_12197_),
    .A(_01028_),
    .B(net6225));
 sg13g2_o21ai_1 _25810_ (.B1(_12197_),
    .Y(_12198_),
    .A1(net5865),
    .A2(net5993));
 sg13g2_mux2_1 _25811_ (.A0(net5773),
    .A1(_01027_),
    .S(_11798_),
    .X(_12199_));
 sg13g2_nand4_1 _25812_ (.B(_06621_),
    .C(net6466),
    .A(net7669),
    .Y(_12200_),
    .D(_09679_));
 sg13g2_nand2_1 _25813_ (.Y(_12201_),
    .A(net7474),
    .B(_10985_));
 sg13g2_nand2_1 _25814_ (.Y(_12202_),
    .A(_01026_),
    .B(net6221));
 sg13g2_o21ai_1 _25815_ (.B1(_12202_),
    .Y(_12203_),
    .A1(net5862),
    .A2(net6221));
 sg13g2_nand2b_1 _25816_ (.Y(_12204_),
    .B(net6384),
    .A_N(net6221));
 sg13g2_nand2_1 _25817_ (.Y(_12205_),
    .A(_01025_),
    .B(net6221));
 sg13g2_o21ai_1 _25818_ (.B1(_12205_),
    .Y(_12206_),
    .A1(net5856),
    .A2(_12204_));
 sg13g2_nand2_1 _25819_ (.Y(_12207_),
    .A(_01024_),
    .B(net6217));
 sg13g2_o21ai_1 _25820_ (.B1(_12207_),
    .Y(_12208_),
    .A1(net5809),
    .A2(net5992));
 sg13g2_nand2_1 _25821_ (.Y(_12209_),
    .A(_01023_),
    .B(net6219));
 sg13g2_o21ai_1 _25822_ (.B1(_12209_),
    .Y(_12210_),
    .A1(net5848),
    .A2(net6219));
 sg13g2_nand2_1 _25823_ (.Y(_12211_),
    .A(_01022_),
    .B(net6220));
 sg13g2_o21ai_1 _25824_ (.B1(_12211_),
    .Y(_12212_),
    .A1(net5798),
    .A2(net6220));
 sg13g2_nand2_1 _25825_ (.Y(_12213_),
    .A(_01021_),
    .B(net6218));
 sg13g2_o21ai_1 _25826_ (.B1(_12213_),
    .Y(_12214_),
    .A1(net5794),
    .A2(_12201_));
 sg13g2_nand2b_1 _25827_ (.Y(_12215_),
    .B(net6377),
    .A_N(net6224));
 sg13g2_nand2_1 _25828_ (.Y(_12216_),
    .A(_01020_),
    .B(_12200_));
 sg13g2_o21ai_1 _25829_ (.B1(_12216_),
    .Y(_12217_),
    .A1(net5920),
    .A2(_12215_));
 sg13g2_nand2_1 _25830_ (.Y(_12218_),
    .A(_01019_),
    .B(net6218));
 sg13g2_o21ai_1 _25831_ (.B1(_12218_),
    .Y(_12219_),
    .A1(net5788),
    .A2(_12201_));
 sg13g2_nand2b_1 _25832_ (.Y(_12220_),
    .B(net6372),
    .A_N(net6221));
 sg13g2_nand2_1 _25833_ (.Y(_12221_),
    .A(_01018_),
    .B(net6221));
 sg13g2_o21ai_1 _25834_ (.B1(_12221_),
    .Y(_12222_),
    .A1(net5914),
    .A2(_12220_));
 sg13g2_nor2_1 _25835_ (.A(_12142_),
    .B(_12190_),
    .Y(_12223_));
 sg13g2_nand2_1 _25836_ (.Y(_12224_),
    .A(_01017_),
    .B(net6217));
 sg13g2_and4_1 _25837_ (.A(_11822_),
    .B(_11932_),
    .C(_12074_),
    .D(_12223_),
    .X(_12225_));
 sg13g2_o21ai_1 _25838_ (.B1(_12224_),
    .Y(_12226_),
    .A1(net5780),
    .A2(net5992));
 sg13g2_nand2_1 _25839_ (.Y(_12227_),
    .A(_01016_),
    .B(net6263));
 sg13g2_nand4_1 _25840_ (.B(_11932_),
    .C(_12074_),
    .A(_11822_),
    .Y(_12228_),
    .D(_12223_));
 sg13g2_o21ai_1 _25841_ (.B1(_12227_),
    .Y(_12229_),
    .A1(net5885),
    .A2(net6263));
 sg13g2_nand2b_1 _25842_ (.Y(_12230_),
    .B(net6367),
    .A_N(net6224));
 sg13g2_nand2_1 _25843_ (.Y(_12231_),
    .A(_01015_),
    .B(_12200_));
 sg13g2_o21ai_1 _25844_ (.B1(_12231_),
    .Y(_12232_),
    .A1(net5909),
    .A2(_12230_));
 sg13g2_mux2_1 _25845_ (.A0(net5843),
    .A1(_01014_),
    .S(net5992),
    .X(_12233_));
 sg13g2_nand2_1 _25846_ (.Y(_12234_),
    .A(_01013_),
    .B(net6218));
 sg13g2_o21ai_1 _25847_ (.B1(_12234_),
    .Y(_12235_),
    .A1(net5834),
    .A2(_12201_));
 sg13g2_nand2_1 _25848_ (.Y(_12236_),
    .A(_01012_),
    .B(net6218));
 sg13g2_o21ai_1 _25849_ (.B1(_12236_),
    .Y(_12237_),
    .A1(net5903),
    .A2(_12201_));
 sg13g2_nand2b_1 _25850_ (.Y(_12238_),
    .B(net8000),
    .A_N(_01635_));
 sg13g2_nand2_1 _25851_ (.Y(_12239_),
    .A(_01011_),
    .B(net6217));
 sg13g2_o21ai_1 _25852_ (.B1(_12239_),
    .Y(_12240_),
    .A1(net5898),
    .A2(net5992));
 sg13g2_nand2_1 _25853_ (.Y(_12241_),
    .A(_01010_),
    .B(net6222));
 sg13g2_o21ai_1 _25854_ (.B1(_12241_),
    .Y(_12242_),
    .A1(net5890),
    .A2(net6222));
 sg13g2_o21ai_1 _25855_ (.B1(_12238_),
    .Y(_12243_),
    .A1(_01638_),
    .A2(net7479));
 sg13g2_mux2_1 _25856_ (.A0(net5774),
    .A1(_01009_),
    .S(_12200_),
    .X(_12244_));
 sg13g2_a21oi_1 _25857_ (.A1(net8006),
    .A2(net7282),
    .Y(_12245_),
    .B1(_12243_));
 sg13g2_nand2_1 _25858_ (.Y(_12246_),
    .A(_01008_),
    .B(net6222));
 sg13g2_o21ai_1 _25859_ (.B1(_12246_),
    .Y(_12247_),
    .A1(net5884),
    .A2(net6222));
 sg13g2_nand2_1 _25860_ (.Y(_12248_),
    .A(_01007_),
    .B(net6220));
 sg13g2_o21ai_1 _25861_ (.B1(_12248_),
    .Y(_12249_),
    .A1(net5926),
    .A2(net6220));
 sg13g2_nand2_1 _25862_ (.Y(_12250_),
    .A(_01006_),
    .B(net6220));
 sg13g2_o21ai_1 _25863_ (.B1(_12250_),
    .Y(_12251_),
    .A1(net5963),
    .A2(net6220));
 sg13g2_nand2_1 _25864_ (.Y(_12252_),
    .A(_01005_),
    .B(net6261));
 sg13g2_o21ai_1 _25865_ (.B1(_12252_),
    .Y(_12253_),
    .A1(net5925),
    .A2(net6261));
 sg13g2_nand2_1 _25866_ (.Y(_12254_),
    .A(_01004_),
    .B(net6223));
 sg13g2_o21ai_1 _25867_ (.B1(_12254_),
    .Y(_12255_),
    .A1(net6015),
    .A2(net6223));
 sg13g2_o21ai_1 _25868_ (.B1(_12245_),
    .Y(_12256_),
    .A1(_09277_),
    .A2(_11665_));
 sg13g2_nand2_1 _25869_ (.Y(_12257_),
    .A(_01003_),
    .B(net6217));
 sg13g2_o21ai_1 _25870_ (.B1(_12257_),
    .Y(_12258_),
    .A1(net5959),
    .A2(net5992));
 sg13g2_nand2_1 _25871_ (.Y(_12259_),
    .A(_01002_),
    .B(net6223));
 sg13g2_o21ai_1 _25872_ (.B1(_12259_),
    .Y(_12260_),
    .A1(net6011),
    .A2(net6223));
 sg13g2_nand2_1 _25873_ (.Y(_12261_),
    .A(_01001_),
    .B(net6223));
 sg13g2_o21ai_1 _25874_ (.B1(_12261_),
    .Y(_12262_),
    .A1(net6005),
    .A2(net6223));
 sg13g2_nand2_1 _25875_ (.Y(_12263_),
    .A(_01000_),
    .B(net6219));
 sg13g2_o21ai_1 _25876_ (.B1(_12263_),
    .Y(_12264_),
    .A1(net6117),
    .A2(net6219));
 sg13g2_nand2_1 _25877_ (.Y(_12265_),
    .A(_00999_),
    .B(net6220));
 sg13g2_o21ai_1 _25878_ (.B1(_12265_),
    .Y(_12266_),
    .A1(net6032),
    .A2(net6220));
 sg13g2_nand2_1 _25879_ (.Y(_12267_),
    .A(_00998_),
    .B(net6219));
 sg13g2_o21ai_1 _25880_ (.B1(_12267_),
    .Y(_12268_),
    .A1(net6112),
    .A2(net6219));
 sg13g2_nand2_1 _25881_ (.Y(_12269_),
    .A(_00997_),
    .B(net6219));
 sg13g2_o21ai_1 _25882_ (.B1(_12269_),
    .Y(_12270_),
    .A1(net6023),
    .A2(net6219));
 sg13g2_a22oi_1 _25883_ (.Y(_12271_),
    .B1(_12256_),
    .B2(net7377),
    .A2(_11682_),
    .A1(net6917));
 sg13g2_nand2_1 _25884_ (.Y(_12272_),
    .A(_00996_),
    .B(net6222));
 sg13g2_o21ai_1 _25885_ (.B1(_12272_),
    .Y(_12273_),
    .A1(net6054),
    .A2(net6222));
 sg13g2_nand2_1 _25886_ (.Y(_12274_),
    .A(_00995_),
    .B(net6223));
 sg13g2_o21ai_1 _25887_ (.B1(_12274_),
    .Y(_12275_),
    .A1(net6021),
    .A2(net6223));
 sg13g2_nand2_1 _25888_ (.Y(_12276_),
    .A(_00994_),
    .B(net6266));
 sg13g2_o21ai_1 _25889_ (.B1(_12276_),
    .Y(_12277_),
    .A1(net5962),
    .A2(net6266));
 sg13g2_nand2_1 _25890_ (.Y(_12278_),
    .A(_00993_),
    .B(net6224));
 sg13g2_o21ai_1 _25891_ (.B1(_12278_),
    .Y(_12279_),
    .A1(net6108),
    .A2(net6224));
 sg13g2_nand2_1 _25892_ (.Y(_12280_),
    .A(_00992_),
    .B(net6217));
 sg13g2_o21ai_1 _25893_ (.B1(_12280_),
    .Y(_12281_),
    .A1(_10088_),
    .A2(net5992));
 sg13g2_nand2_2 _25894_ (.Y(_12282_),
    .A(_09679_),
    .B(_11799_));
 sg13g2_nand2_1 _25895_ (.Y(_12283_),
    .A(_00991_),
    .B(net6074));
 sg13g2_o21ai_1 _25896_ (.B1(_12283_),
    .Y(_12284_),
    .A1(net5862),
    .A2(net6074));
 sg13g2_nand3_1 _25897_ (.B(_10162_),
    .C(net6259),
    .A(_09679_),
    .Y(_12285_));
 sg13g2_o21ai_1 _25898_ (.B1(_12271_),
    .Y(_12286_),
    .A1(net6981),
    .A2(_11682_));
 sg13g2_nand2_1 _25899_ (.Y(_12287_),
    .A(_00990_),
    .B(net6074));
 sg13g2_o21ai_1 _25900_ (.B1(_12287_),
    .Y(_12288_),
    .A1(net5854),
    .A2(_12285_));
 sg13g2_nand2_1 _25901_ (.Y(_12289_),
    .A(_00989_),
    .B(net6080));
 sg13g2_o21ai_1 _25902_ (.B1(_12289_),
    .Y(_12290_),
    .A1(net5806),
    .A2(net6080));
 sg13g2_nand2_1 _25903_ (.Y(_12291_),
    .A(_00988_),
    .B(net6073));
 sg13g2_o21ai_1 _25904_ (.B1(_12291_),
    .Y(_12292_),
    .A1(net5848),
    .A2(net6073));
 sg13g2_nand2_1 _25905_ (.Y(_12293_),
    .A(_00987_),
    .B(net6077));
 sg13g2_o21ai_1 _25906_ (.B1(_12293_),
    .Y(_12294_),
    .A1(net5798),
    .A2(net6077));
 sg13g2_nand2_1 _25907_ (.Y(_12295_),
    .A(_00986_),
    .B(net6079));
 sg13g2_o21ai_1 _25908_ (.B1(_12295_),
    .Y(_12296_),
    .A1(net5794),
    .A2(net6079));
 sg13g2_nand3_1 _25909_ (.B(_10341_),
    .C(net6259),
    .A(_09679_),
    .Y(_12297_));
 sg13g2_nand2_1 _25910_ (.Y(_12298_),
    .A(_00985_),
    .B(net6074));
 sg13g2_o21ai_1 _25911_ (.B1(_12298_),
    .Y(_12299_),
    .A1(net5920),
    .A2(_12297_));
 sg13g2_nand2_1 _25912_ (.Y(_12300_),
    .A(_00984_),
    .B(net6079));
 sg13g2_o21ai_1 _25913_ (.B1(_12300_),
    .Y(_12301_),
    .A1(net5788),
    .A2(net6079));
 sg13g2_nand2_1 _25914_ (.Y(_12302_),
    .A(_00983_),
    .B(net6265));
 sg13g2_o21ai_1 _25915_ (.B1(_12302_),
    .Y(_12303_),
    .A1(net6014),
    .A2(net6265));
 sg13g2_nand3_1 _25916_ (.B(_10415_),
    .C(net6259),
    .A(_09679_),
    .Y(_12304_));
 sg13g2_nand2_1 _25917_ (.Y(_12305_),
    .A(_00982_),
    .B(net6074));
 sg13g2_o21ai_1 _25918_ (.B1(_12305_),
    .Y(_12306_),
    .A1(net5914),
    .A2(_12304_));
 sg13g2_nand2_1 _25919_ (.Y(_12307_),
    .A(_00981_),
    .B(net6080));
 sg13g2_o21ai_1 _25920_ (.B1(_12307_),
    .Y(_12308_),
    .A1(net5779),
    .A2(net6080));
 sg13g2_nand3_1 _25921_ (.B(net6367),
    .C(net6259),
    .A(_09679_),
    .Y(_12309_));
 sg13g2_nand2_1 _25922_ (.Y(_12310_),
    .A(_00980_),
    .B(net6074));
 sg13g2_o21ai_1 _25923_ (.B1(_12310_),
    .Y(_12311_),
    .A1(net5909),
    .A2(_12309_));
 sg13g2_mux2_1 _25924_ (.A0(net5843),
    .A1(_00979_),
    .S(net6081),
    .X(_12312_));
 sg13g2_nand2_1 _25925_ (.Y(_12313_),
    .A(_00978_),
    .B(net6082));
 sg13g2_o21ai_1 _25926_ (.B1(_12313_),
    .Y(_12314_),
    .A1(net5833),
    .A2(net6082));
 sg13g2_nand2_1 _25927_ (.Y(_12315_),
    .A(_00977_),
    .B(net6079));
 sg13g2_o21ai_1 _25928_ (.B1(_12315_),
    .Y(_12316_),
    .A1(net5904),
    .A2(net6079));
 sg13g2_nand2_1 _25929_ (.Y(_12317_),
    .A(_00976_),
    .B(net6080));
 sg13g2_o21ai_1 _25930_ (.B1(_12317_),
    .Y(_12318_),
    .A1(net5898),
    .A2(net6080));
 sg13g2_nand2_1 _25931_ (.Y(_12319_),
    .A(_00975_),
    .B(net6082));
 sg13g2_o21ai_1 _25932_ (.B1(_12319_),
    .Y(_12320_),
    .A1(net5890),
    .A2(net6075));
 sg13g2_mux2_1 _25933_ (.A0(net5773),
    .A1(_00974_),
    .S(net6074),
    .X(_12321_));
 sg13g2_nand2_1 _25934_ (.Y(_12322_),
    .A(_00973_),
    .B(net6075));
 sg13g2_o21ai_1 _25935_ (.B1(_12322_),
    .Y(_12323_),
    .A1(net5886),
    .A2(net6075));
 sg13g2_nand2_1 _25936_ (.Y(_12324_),
    .A(_00972_),
    .B(net6264));
 sg13g2_o21ai_1 _25937_ (.B1(_12324_),
    .Y(_12325_),
    .A1(net5957),
    .A2(net6095));
 sg13g2_nand2_1 _25938_ (.Y(_12326_),
    .A(_00971_),
    .B(net6077));
 sg13g2_o21ai_1 _25939_ (.B1(_12326_),
    .Y(_12327_),
    .A1(net5926),
    .A2(net6077));
 sg13g2_nand2_1 _25940_ (.Y(_12328_),
    .A(_00970_),
    .B(net6077));
 sg13g2_o21ai_1 _25941_ (.B1(_12328_),
    .Y(_12329_),
    .A1(net5963),
    .A2(net6077));
 sg13g2_nand2_1 _25942_ (.Y(_12330_),
    .A(_00969_),
    .B(net6078));
 sg13g2_a221oi_1 _25943_ (.B2(_01888_),
    .C1(_08614_),
    .B1(_09397_),
    .A1(net7685),
    .Y(_12331_),
    .A2(_08800_));
 sg13g2_o21ai_1 _25944_ (.B1(_12330_),
    .Y(_12332_),
    .A1(net6015),
    .A2(net6078));
 sg13g2_nand2_1 _25945_ (.Y(_12333_),
    .A(_00968_),
    .B(net6081));
 sg13g2_o21ai_1 _25946_ (.B1(_12333_),
    .Y(_12334_),
    .A1(net5961),
    .A2(net6081));
 sg13g2_nand2_1 _25947_ (.Y(_12335_),
    .A(_00967_),
    .B(net6078));
 sg13g2_o21ai_1 _25948_ (.B1(_12335_),
    .Y(_12336_),
    .A1(net6011),
    .A2(net6078));
 sg13g2_nand2_1 _25949_ (.Y(_12337_),
    .A(_00966_),
    .B(net6076));
 sg13g2_o21ai_1 _25950_ (.B1(_12337_),
    .Y(_12338_),
    .A1(net6001),
    .A2(net6076));
 sg13g2_nand2_1 _25951_ (.Y(_12339_),
    .A(_00965_),
    .B(net6073));
 sg13g2_o21ai_1 _25952_ (.B1(_12339_),
    .Y(_12340_),
    .A1(net6117),
    .A2(net6073));
 sg13g2_nand2_1 _25953_ (.Y(_12341_),
    .A(_00964_),
    .B(net6077));
 sg13g2_o21ai_1 _25954_ (.B1(_12341_),
    .Y(_12342_),
    .A1(net6032),
    .A2(net6078));
 sg13g2_nand2_1 _25955_ (.Y(_12343_),
    .A(_00963_),
    .B(net6073));
 sg13g2_o21ai_1 _25956_ (.B1(_12343_),
    .Y(_12344_),
    .A1(net6112),
    .A2(net6073));
 sg13g2_nand2_1 _25957_ (.Y(_12345_),
    .A(_00962_),
    .B(net6073));
 sg13g2_o21ai_1 _25958_ (.B1(_12345_),
    .Y(_12346_),
    .A1(net6023),
    .A2(net6073));
 sg13g2_nand2_1 _25959_ (.Y(_12347_),
    .A(_00961_),
    .B(net6265));
 sg13g2_o21ai_1 _25960_ (.B1(_12347_),
    .Y(_12348_),
    .A1(net6010),
    .A2(net6265));
 sg13g2_nand2_1 _25961_ (.Y(_12349_),
    .A(_00960_),
    .B(net6075));
 sg13g2_o21ai_1 _25962_ (.B1(_12349_),
    .Y(_12350_),
    .A1(net6054),
    .A2(net6075));
 sg13g2_nand2_1 _25963_ (.Y(_12351_),
    .A(_00959_),
    .B(net6076));
 sg13g2_o21ai_1 _25964_ (.B1(_12351_),
    .Y(_12352_),
    .A1(net6021),
    .A2(net6076));
 sg13g2_nand2_1 _25965_ (.Y(_12353_),
    .A(_00958_),
    .B(net6075));
 sg13g2_o21ai_1 _25966_ (.B1(_12353_),
    .Y(_12354_),
    .A1(net6107),
    .A2(net6075));
 sg13g2_nand2_1 _25967_ (.Y(_12355_),
    .A(_00957_),
    .B(net6080));
 sg13g2_o21ai_1 _25968_ (.B1(_12355_),
    .Y(_12356_),
    .A1(net5865),
    .A2(net6080));
 sg13g2_or4_1 _25969_ (.A(net7670),
    .B(_06622_),
    .C(net6467),
    .D(_09680_),
    .X(_12357_));
 sg13g2_nand3_1 _25970_ (.B(net7474),
    .C(_10990_),
    .A(_06621_),
    .Y(_12358_));
 sg13g2_nand2_1 _25971_ (.Y(_12359_),
    .A(_00956_),
    .B(net6210));
 sg13g2_o21ai_1 _25972_ (.B1(_12359_),
    .Y(_12360_),
    .A1(net5862),
    .A2(net6210));
 sg13g2_nand2_1 _25973_ (.Y(_12361_),
    .A(_00955_),
    .B(net6210));
 sg13g2_nand2b_1 _25974_ (.Y(_12362_),
    .B(net6382),
    .A_N(net6210));
 sg13g2_o21ai_1 _25975_ (.B1(_12361_),
    .Y(_12363_),
    .A1(net5858),
    .A2(_12362_));
 sg13g2_nand2_1 _25976_ (.Y(_12364_),
    .A(_00954_),
    .B(net6216));
 sg13g2_o21ai_1 _25977_ (.B1(_12364_),
    .Y(_12365_),
    .A1(net5806),
    .A2(net6072));
 sg13g2_nand2_1 _25978_ (.Y(_12366_),
    .A(_00953_),
    .B(net6209));
 sg13g2_o21ai_1 _25979_ (.B1(_12366_),
    .Y(_12367_),
    .A1(net5848),
    .A2(net6209));
 sg13g2_nand2_1 _25980_ (.Y(_12368_),
    .A(_00952_),
    .B(net6214));
 sg13g2_o21ai_1 _25981_ (.B1(_12368_),
    .Y(_12369_),
    .A1(net5798),
    .A2(net6214));
 sg13g2_nand2_1 _25982_ (.Y(_12370_),
    .A(_00951_),
    .B(_12357_));
 sg13g2_o21ai_1 _25983_ (.B1(_12370_),
    .Y(_12371_),
    .A1(net5794),
    .A2(_12358_));
 sg13g2_nand2_1 _25984_ (.Y(_12372_),
    .A(_00950_),
    .B(net6265));
 sg13g2_o21ai_1 _25985_ (.B1(_12372_),
    .Y(_12373_),
    .A1(net6006),
    .A2(net6265));
 sg13g2_nand2_1 _25986_ (.Y(_12374_),
    .A(_00949_),
    .B(net6210));
 sg13g2_nand2b_1 _25987_ (.Y(_12375_),
    .B(net6378),
    .A_N(net6215));
 sg13g2_o21ai_1 _25988_ (.B1(_12374_),
    .Y(_12376_),
    .A1(net5920),
    .A2(_12375_));
 sg13g2_nand2_1 _25989_ (.Y(_12377_),
    .A(_00948_),
    .B(net6216));
 sg13g2_o21ai_1 _25990_ (.B1(_12377_),
    .Y(_12378_),
    .A1(net5788),
    .A2(_12358_));
 sg13g2_nand2b_1 _25991_ (.Y(_12379_),
    .B(net6372),
    .A_N(_12357_));
 sg13g2_nand2_1 _25992_ (.Y(_12380_),
    .A(_00947_),
    .B(_12357_));
 sg13g2_o21ai_1 _25993_ (.B1(_12380_),
    .Y(_12381_),
    .A1(net5914),
    .A2(_12379_));
 sg13g2_nand2_1 _25994_ (.Y(_12382_),
    .A(_00946_),
    .B(net6216));
 sg13g2_o21ai_1 _25995_ (.B1(_12382_),
    .Y(_12383_),
    .A1(net5779),
    .A2(net6072));
 sg13g2_nand2_1 _25996_ (.Y(_12384_),
    .A(_00945_),
    .B(_12357_));
 sg13g2_nand2b_1 _25997_ (.Y(_12385_),
    .B(net6367),
    .A_N(net6210));
 sg13g2_mux4_1 _25998_ (.S0(net7795),
    .A0(_00792_),
    .A1(_00824_),
    .A2(_00856_),
    .A3(_00891_),
    .S1(net7738),
    .X(_12386_));
 sg13g2_o21ai_1 _25999_ (.B1(_12384_),
    .Y(_12387_),
    .A1(net5909),
    .A2(_12385_));
 sg13g2_and2_1 _26000_ (.A(net7604),
    .B(_12386_),
    .X(_12388_));
 sg13g2_mux2_1 _26001_ (.A0(net5841),
    .A1(_00944_),
    .S(_12358_),
    .X(_12389_));
 sg13g2_nand2_1 _26002_ (.Y(_12390_),
    .A(_00943_),
    .B(net6216));
 sg13g2_o21ai_1 _26003_ (.B1(_12390_),
    .Y(_12391_),
    .A1(net5834),
    .A2(_12358_));
 sg13g2_nand2_1 _26004_ (.Y(_12392_),
    .A(_00942_),
    .B(net6216));
 sg13g2_nand2_1 _26005_ (.Y(_12393_),
    .A(net7708),
    .B(_00760_));
 sg13g2_o21ai_1 _26006_ (.B1(_12392_),
    .Y(_12394_),
    .A1(net5904),
    .A2(net6072));
 sg13g2_nand2_1 _26007_ (.Y(_12395_),
    .A(_00941_),
    .B(net6216));
 sg13g2_o21ai_1 _26008_ (.B1(_12395_),
    .Y(_12396_),
    .A1(net5898),
    .A2(_12358_));
 sg13g2_nand2b_1 _26009_ (.Y(_12397_),
    .B(_00618_),
    .A_N(net7708));
 sg13g2_nand2_1 _26010_ (.Y(_12398_),
    .A(_00940_),
    .B(net6211));
 sg13g2_o21ai_1 _26011_ (.B1(_12398_),
    .Y(_12399_),
    .A1(net5890),
    .A2(net6211));
 sg13g2_nand2_1 _26012_ (.Y(_12400_),
    .A(_00939_),
    .B(net6260));
 sg13g2_o21ai_1 _26013_ (.B1(_12400_),
    .Y(_12401_),
    .A1(net6117),
    .A2(net6260));
 sg13g2_a21oi_1 _26014_ (.A1(_12393_),
    .A2(_12397_),
    .Y(_12402_),
    .B1(net7600));
 sg13g2_mux2_1 _26015_ (.A0(net5773),
    .A1(_00938_),
    .S(_12357_),
    .X(_12403_));
 sg13g2_nand2_1 _26016_ (.Y(_12404_),
    .A(_00937_),
    .B(net6211));
 sg13g2_o21ai_1 _26017_ (.B1(_12404_),
    .Y(_12405_),
    .A1(net5886),
    .A2(net6211));
 sg13g2_nand2_1 _26018_ (.Y(_12406_),
    .A(_00936_),
    .B(net6214));
 sg13g2_o21ai_1 _26019_ (.B1(_12406_),
    .Y(_12407_),
    .A1(net5926),
    .A2(net6214));
 sg13g2_nand2_1 _26020_ (.Y(_12408_),
    .A(_00935_),
    .B(net6214));
 sg13g2_o21ai_1 _26021_ (.B1(_12408_),
    .Y(_12409_),
    .A1(net5963),
    .A2(net6214));
 sg13g2_nand2_1 _26022_ (.Y(_12410_),
    .A(_00934_),
    .B(net6213));
 sg13g2_nand3b_1 _26023_ (.B(net7796),
    .C(_00906_),
    .Y(_12411_),
    .A_N(net7738));
 sg13g2_o21ai_1 _26024_ (.B1(_12410_),
    .Y(_12412_),
    .A1(net6012),
    .A2(net6213));
 sg13g2_nand2_1 _26025_ (.Y(_12413_),
    .A(_00933_),
    .B(net6216));
 sg13g2_o21ai_1 _26026_ (.B1(_12413_),
    .Y(_12414_),
    .A1(net5959),
    .A2(_12358_));
 sg13g2_nand2_1 _26027_ (.Y(_12415_),
    .A(_00932_),
    .B(net6212));
 sg13g2_nand3b_1 _26028_ (.B(_01258_),
    .C(net7738),
    .Y(_12416_),
    .A_N(net7796));
 sg13g2_o21ai_1 _26029_ (.B1(_12415_),
    .Y(_12417_),
    .A1(net6011),
    .A2(net6213));
 sg13g2_nand2_1 _26030_ (.Y(_12418_),
    .A(_00931_),
    .B(net6211));
 sg13g2_o21ai_1 _26031_ (.B1(_12418_),
    .Y(_12419_),
    .A1(net6002),
    .A2(net6212));
 sg13g2_nand2_1 _26032_ (.Y(_12420_),
    .A(_00930_),
    .B(net6209));
 sg13g2_a21oi_1 _26033_ (.A1(_12411_),
    .A2(_12416_),
    .Y(_12421_),
    .B1(net7598));
 sg13g2_o21ai_1 _26034_ (.B1(_12420_),
    .Y(_12422_),
    .A1(net6117),
    .A2(net6209));
 sg13g2_nand2_1 _26035_ (.Y(_12423_),
    .A(_00929_),
    .B(net6214));
 sg13g2_o21ai_1 _26036_ (.B1(_12423_),
    .Y(_12424_),
    .A1(net6032),
    .A2(net6214));
 sg13g2_nand2_1 _26037_ (.Y(_12425_),
    .A(_00928_),
    .B(net6266));
 sg13g2_o21ai_1 _26038_ (.B1(_12425_),
    .Y(_12426_),
    .A1(net6033),
    .A2(net6266));
 sg13g2_nand2_1 _26039_ (.Y(_12427_),
    .A(_00927_),
    .B(net6209));
 sg13g2_o21ai_1 _26040_ (.B1(_12427_),
    .Y(_12428_),
    .A1(net6112),
    .A2(net6209));
 sg13g2_nor4_1 _26041_ (.A(net7690),
    .B(_12388_),
    .C(_12402_),
    .D(_12421_),
    .Y(_12429_));
 sg13g2_nand2_1 _26042_ (.Y(_12430_),
    .A(_00926_),
    .B(net6209));
 sg13g2_o21ai_1 _26043_ (.B1(_12430_),
    .Y(_12431_),
    .A1(net6023),
    .A2(net6209));
 sg13g2_nand2_1 _26044_ (.Y(_12432_),
    .A(_00925_),
    .B(net6211));
 sg13g2_o21ai_1 _26045_ (.B1(_12432_),
    .Y(_12433_),
    .A1(net6054),
    .A2(net6211));
 sg13g2_nand2_1 _26046_ (.Y(_12434_),
    .A(_00924_),
    .B(net6212));
 sg13g2_o21ai_1 _26047_ (.B1(_12434_),
    .Y(_12435_),
    .A1(net6021),
    .A2(net6212));
 sg13g2_nand2_1 _26048_ (.Y(_12436_),
    .A(_00923_),
    .B(net6215));
 sg13g2_o21ai_1 _26049_ (.B1(_12436_),
    .Y(_12437_),
    .A1(_10022_),
    .A2(net6215));
 sg13g2_nand2_1 _26050_ (.Y(_12438_),
    .A(_00922_),
    .B(net6216));
 sg13g2_o21ai_1 _26051_ (.B1(_12438_),
    .Y(_12439_),
    .A1(net5865),
    .A2(_12358_));
 sg13g2_nor2_1 _26052_ (.A(_09609_),
    .B(_11159_),
    .Y(_12440_));
 sg13g2_nand2_1 _26053_ (.Y(_12441_),
    .A(_09608_),
    .B(net7447));
 sg13g2_mux2_1 _26054_ (.A0(_00664_),
    .A1(_00696_),
    .S(net7796),
    .X(_12442_));
 sg13g2_nand2_1 _26055_ (.Y(_12443_),
    .A(_00921_),
    .B(net5982));
 sg13g2_o21ai_1 _26056_ (.B1(_12443_),
    .Y(_12444_),
    .A1(net5861),
    .A2(_12441_));
 sg13g2_nand2_1 _26057_ (.Y(_12445_),
    .A(net6382),
    .B(_12440_));
 sg13g2_nand2_1 _26058_ (.Y(_12446_),
    .A(_00920_),
    .B(net5982));
 sg13g2_o21ai_1 _26059_ (.B1(_12446_),
    .Y(_12447_),
    .A1(net5853),
    .A2(_12445_));
 sg13g2_nand2_1 _26060_ (.Y(_12448_),
    .A(_00919_),
    .B(net5984));
 sg13g2_o21ai_1 _26061_ (.B1(_12448_),
    .Y(_12449_),
    .A1(net5804),
    .A2(net5985));
 sg13g2_nand2_1 _26062_ (.Y(_12450_),
    .A(_00918_),
    .B(net5983));
 sg13g2_o21ai_1 _26063_ (.B1(_12450_),
    .Y(_12451_),
    .A1(net5851),
    .A2(net5983));
 sg13g2_nand2_1 _26064_ (.Y(_12452_),
    .A(_00917_),
    .B(net6261));
 sg13g2_o21ai_1 _26065_ (.B1(_12452_),
    .Y(_12453_),
    .A1(net6110),
    .A2(net6261));
 sg13g2_nand2_1 _26066_ (.Y(_12454_),
    .A(_00916_),
    .B(net5990));
 sg13g2_o21ai_1 _26067_ (.B1(_12454_),
    .Y(_12455_),
    .A1(net5799),
    .A2(net5990));
 sg13g2_nand2_1 _26068_ (.Y(_12456_),
    .A(_00915_),
    .B(net5986));
 sg13g2_o21ai_1 _26069_ (.B1(_12456_),
    .Y(_12457_),
    .A1(net5793),
    .A2(net5986));
 sg13g2_nand2_1 _26070_ (.Y(_12458_),
    .A(_00914_),
    .B(net5982));
 sg13g2_nand2_1 _26071_ (.Y(_12459_),
    .A(net6377),
    .B(_12440_));
 sg13g2_o21ai_1 _26072_ (.B1(_12458_),
    .Y(_12460_),
    .A1(net5921),
    .A2(_12459_));
 sg13g2_nand2_1 _26073_ (.Y(_12461_),
    .A(_00913_),
    .B(net5984));
 sg13g2_o21ai_1 _26074_ (.B1(_12461_),
    .Y(_12462_),
    .A1(net5787),
    .A2(net5984));
 sg13g2_nand2_1 _26075_ (.Y(_12463_),
    .A(net6374),
    .B(_12440_));
 sg13g2_a22oi_1 _26076_ (.Y(_12464_),
    .B1(_12442_),
    .B2(net7516),
    .A2(net7595),
    .A1(_00728_));
 sg13g2_nand2_1 _26077_ (.Y(_12465_),
    .A(_00912_),
    .B(net5982));
 sg13g2_o21ai_1 _26078_ (.B1(_12465_),
    .Y(_12466_),
    .A1(net5914),
    .A2(_12463_));
 sg13g2_nand2_1 _26079_ (.Y(_12467_),
    .A(_00911_),
    .B(net5985));
 sg13g2_o21ai_1 _26080_ (.B1(_12467_),
    .Y(_12468_),
    .A1(net5783),
    .A2(net5985));
 sg13g2_nand2_1 _26081_ (.Y(_12469_),
    .A(net6368),
    .B(_12440_));
 sg13g2_nand2_1 _26082_ (.Y(_12470_),
    .A(_00910_),
    .B(net5982));
 sg13g2_o21ai_1 _26083_ (.B1(_12470_),
    .Y(_12471_),
    .A1(net5911),
    .A2(_12469_));
 sg13g2_mux2_1 _26084_ (.A0(_00909_),
    .A1(net5838),
    .S(_12440_),
    .X(_12472_));
 sg13g2_nand2_1 _26085_ (.Y(_12473_),
    .A(_00908_),
    .B(net5986));
 sg13g2_o21ai_1 _26086_ (.B1(_12473_),
    .Y(_12474_),
    .A1(net5833),
    .A2(net5986));
 sg13g2_nand2_1 _26087_ (.Y(_12475_),
    .A(_00907_),
    .B(net5984));
 sg13g2_o21ai_1 _26088_ (.B1(_12475_),
    .Y(_12476_),
    .A1(net5902),
    .A2(net5984));
 sg13g2_nand2_1 _26089_ (.Y(_12477_),
    .A(_00906_),
    .B(net6260));
 sg13g2_o21ai_1 _26090_ (.B1(_12477_),
    .Y(_12478_),
    .A1(_09902_),
    .A2(net6260));
 sg13g2_nand2_1 _26091_ (.Y(_12479_),
    .A(_00905_),
    .B(net5985));
 sg13g2_o21ai_1 _26092_ (.B1(_12479_),
    .Y(_12480_),
    .A1(net5899),
    .A2(net5985));
 sg13g2_nand2_1 _26093_ (.Y(_12481_),
    .A(_00904_),
    .B(net5987));
 sg13g2_o21ai_1 _26094_ (.B1(_12481_),
    .Y(_12482_),
    .A1(net5889),
    .A2(net5987));
 sg13g2_mux2_1 _26095_ (.A0(_00903_),
    .A1(net5772),
    .S(_12440_),
    .X(_12483_));
 sg13g2_nand2_1 _26096_ (.Y(_12484_),
    .A(_00902_),
    .B(net5991));
 sg13g2_o21ai_1 _26097_ (.B1(_12484_),
    .Y(_12485_),
    .A1(net5884),
    .A2(net5987));
 sg13g2_nand2_1 _26098_ (.Y(_12486_),
    .A(_00901_),
    .B(net5990));
 sg13g2_o21ai_1 _26099_ (.B1(_12486_),
    .Y(_12487_),
    .A1(net5926),
    .A2(net5990));
 sg13g2_nand2_1 _26100_ (.Y(_12488_),
    .A(_00900_),
    .B(net5990));
 sg13g2_o21ai_1 _26101_ (.B1(_12488_),
    .Y(_12489_),
    .A1(net5963),
    .A2(net5990));
 sg13g2_nand2_1 _26102_ (.Y(_12490_),
    .A(_00899_),
    .B(net5989));
 sg13g2_o21ai_1 _26103_ (.B1(_12490_),
    .Y(_12491_),
    .A1(net6015),
    .A2(net5989));
 sg13g2_nand2_1 _26104_ (.Y(_12492_),
    .A(_00898_),
    .B(net5984));
 sg13g2_o21ai_1 _26105_ (.B1(_12492_),
    .Y(_12493_),
    .A1(net5959),
    .A2(net5984));
 sg13g2_nand2_1 _26106_ (.Y(_12494_),
    .A(_00897_),
    .B(net5988));
 sg13g2_o21ai_1 _26107_ (.B1(_12494_),
    .Y(_12495_),
    .A1(_10929_),
    .A2(net5988));
 sg13g2_nand2_1 _26108_ (.Y(_12496_),
    .A(_00896_),
    .B(net5988));
 sg13g2_o21ai_1 _26109_ (.B1(_12496_),
    .Y(_12497_),
    .A1(net6001),
    .A2(net5988));
 sg13g2_nand2_1 _26110_ (.Y(_12498_),
    .A(_00895_),
    .B(net6263));
 sg13g2_o21ai_1 _26111_ (.B1(_12498_),
    .Y(_12499_),
    .A1(net6055),
    .A2(net6263));
 sg13g2_nand2_1 _26112_ (.Y(_12500_),
    .A(_00894_),
    .B(net5983));
 sg13g2_o21ai_1 _26113_ (.B1(_12500_),
    .Y(_12501_),
    .A1(net6118),
    .A2(net5983));
 sg13g2_nand2_1 _26114_ (.Y(_12502_),
    .A(_00893_),
    .B(net5989));
 sg13g2_o21ai_1 _26115_ (.B1(_12502_),
    .Y(_12503_),
    .A1(net6031),
    .A2(net5989));
 sg13g2_nand2_1 _26116_ (.Y(_12504_),
    .A(_00892_),
    .B(net5983));
 sg13g2_o21ai_1 _26117_ (.B1(_12504_),
    .Y(_12505_),
    .A1(net6112),
    .A2(net5983));
 sg13g2_nand2_1 _26118_ (.Y(_12506_),
    .A(_00891_),
    .B(net5983));
 sg13g2_o21ai_1 _26119_ (.B1(_12506_),
    .Y(_12507_),
    .A1(net6023),
    .A2(net5983));
 sg13g2_nand2_1 _26120_ (.Y(_12508_),
    .A(_00890_),
    .B(net5987));
 sg13g2_o21ai_1 _26121_ (.B1(_12508_),
    .Y(_12509_),
    .A1(net6051),
    .A2(net5987));
 sg13g2_nand2_1 _26122_ (.Y(_12510_),
    .A(_00889_),
    .B(net5988));
 sg13g2_o21ai_1 _26123_ (.B1(_12510_),
    .Y(_12511_),
    .A1(net6021),
    .A2(net5988));
 sg13g2_nand2_1 _26124_ (.Y(_12512_),
    .A(_00888_),
    .B(net5988));
 sg13g2_o21ai_1 _26125_ (.B1(_12512_),
    .Y(_12513_),
    .A1(net6107),
    .A2(net5988));
 sg13g2_nand2_1 _26126_ (.Y(_12514_),
    .A(_00887_),
    .B(net5985));
 sg13g2_o21ai_1 _26127_ (.B1(_12514_),
    .Y(_12515_),
    .A1(net5864),
    .A2(net5985));
 sg13g2_nand4_1 _26128_ (.B(_06621_),
    .C(net6466),
    .A(net7670),
    .Y(_12516_),
    .D(_11158_));
 sg13g2_nand2_1 _26129_ (.Y(_12517_),
    .A(_10985_),
    .B(net7447));
 sg13g2_nand2_1 _26130_ (.Y(_12518_),
    .A(_00886_),
    .B(net6202));
 sg13g2_o21ai_1 _26131_ (.B1(_12518_),
    .Y(_12519_),
    .A1(net5861),
    .A2(net6202));
 sg13g2_nand2_1 _26132_ (.Y(_12520_),
    .A(_00885_),
    .B(net6202));
 sg13g2_nand2b_1 _26133_ (.Y(_12521_),
    .B(net6381),
    .A_N(net6202));
 sg13g2_o21ai_1 _26134_ (.B1(_12520_),
    .Y(_12522_),
    .A1(net5855),
    .A2(_12521_));
 sg13g2_nand2_1 _26135_ (.Y(_12523_),
    .A(_00884_),
    .B(net6267));
 sg13g2_o21ai_1 _26136_ (.B1(_12523_),
    .Y(_12524_),
    .A1(net6022),
    .A2(net6267));
 sg13g2_nand2_1 _26137_ (.Y(_12525_),
    .A(_00883_),
    .B(net6207));
 sg13g2_o21ai_1 _26138_ (.B1(_12525_),
    .Y(_12526_),
    .A1(net5805),
    .A2(net5981));
 sg13g2_nand2_1 _26139_ (.Y(_12527_),
    .A(_00882_),
    .B(net6201));
 sg13g2_o21ai_1 _26140_ (.B1(_12527_),
    .Y(_12528_),
    .A1(net5848),
    .A2(net6201));
 sg13g2_nand2_1 _26141_ (.Y(_12529_),
    .A(_00881_),
    .B(net6205));
 sg13g2_o21ai_1 _26142_ (.B1(_12529_),
    .Y(_12530_),
    .A1(net5798),
    .A2(net6205));
 sg13g2_nand2_1 _26143_ (.Y(_12531_),
    .A(_00880_),
    .B(net6208));
 sg13g2_o21ai_1 _26144_ (.B1(_12531_),
    .Y(_12532_),
    .A1(net5793),
    .A2(_12517_));
 sg13g2_nand2_1 _26145_ (.Y(_12533_),
    .A(_00879_),
    .B(net6203));
 sg13g2_mux4_1 _26146_ (.S0(net7794),
    .A0(_00926_),
    .A1(_00962_),
    .A2(_00997_),
    .A3(_01032_),
    .S1(net7738),
    .X(_12534_));
 sg13g2_nand2b_1 _26147_ (.Y(_12535_),
    .B(net6378),
    .A_N(net6203));
 sg13g2_o21ai_1 _26148_ (.B1(_12533_),
    .Y(_12536_),
    .A1(net5917),
    .A2(_12535_));
 sg13g2_nand2_1 _26149_ (.Y(_12537_),
    .A(_00878_),
    .B(net6207));
 sg13g2_o21ai_1 _26150_ (.B1(_12537_),
    .Y(_12538_),
    .A1(net5787),
    .A2(_12517_));
 sg13g2_nand2_1 _26151_ (.Y(_12539_),
    .A(_00877_),
    .B(net6202));
 sg13g2_nand2b_1 _26152_ (.Y(_12540_),
    .B(net6371),
    .A_N(net6202));
 sg13g2_o21ai_1 _26153_ (.B1(_12539_),
    .Y(_12541_),
    .A1(net5913),
    .A2(_12540_));
 sg13g2_nand2_1 _26154_ (.Y(_12542_),
    .A(_00876_),
    .B(net6207));
 sg13g2_o21ai_1 _26155_ (.B1(net7707),
    .Y(_12543_),
    .A1(net7531),
    .A2(_12534_));
 sg13g2_o21ai_1 _26156_ (.B1(_12542_),
    .Y(_12544_),
    .A1(net5782),
    .A2(net5981));
 sg13g2_nand2_1 _26157_ (.Y(_12545_),
    .A(_00875_),
    .B(net6203));
 sg13g2_nand2b_1 _26158_ (.Y(_12546_),
    .B(net6365),
    .A_N(net6203));
 sg13g2_o21ai_1 _26159_ (.B1(_12545_),
    .Y(_12547_),
    .A1(net5907),
    .A2(_12546_));
 sg13g2_mux2_1 _26160_ (.A0(net5839),
    .A1(_00874_),
    .S(net5981),
    .X(_12548_));
 sg13g2_nand2_1 _26161_ (.Y(_12549_),
    .A(_00873_),
    .B(net6267));
 sg13g2_o21ai_1 _26162_ (.B1(_12549_),
    .Y(_12550_),
    .A1(net6108),
    .A2(net6267));
 sg13g2_nand2_1 _26163_ (.Y(_12551_),
    .A(_00872_),
    .B(net6208));
 sg13g2_o21ai_1 _26164_ (.B1(_12551_),
    .Y(_12552_),
    .A1(net5837),
    .A2(_12517_));
 sg13g2_a21o_1 _26165_ (.A2(_12464_),
    .A1(net7531),
    .B1(_12543_),
    .X(_12553_));
 sg13g2_nand2_1 _26166_ (.Y(_12554_),
    .A(_00871_),
    .B(net6207));
 sg13g2_o21ai_1 _26167_ (.B1(_12554_),
    .Y(_12555_),
    .A1(net5903),
    .A2(_12517_));
 sg13g2_nand2_1 _26168_ (.Y(_12556_),
    .A(_00870_),
    .B(net6207));
 sg13g2_o21ai_1 _26169_ (.B1(_12556_),
    .Y(_12557_),
    .A1(net5897),
    .A2(net5981));
 sg13g2_nand2_1 _26170_ (.Y(_12558_),
    .A(_12429_),
    .B(_12553_));
 sg13g2_nand2_1 _26171_ (.Y(_12559_),
    .A(_00869_),
    .B(net6208));
 sg13g2_o21ai_1 _26172_ (.B1(_12559_),
    .Y(_12560_),
    .A1(net5889),
    .A2(net6208));
 sg13g2_mux2_1 _26173_ (.A0(net5773),
    .A1(_00868_),
    .S(net6203),
    .X(_12561_));
 sg13g2_nand2_1 _26174_ (.Y(_12562_),
    .A(_00867_),
    .B(net6204));
 sg13g2_o21ai_1 _26175_ (.B1(_12562_),
    .Y(_12563_),
    .A1(net5885),
    .A2(net6204));
 sg13g2_nand2_1 _26176_ (.Y(_12564_),
    .A(_00866_),
    .B(net6205));
 sg13g2_o21ai_1 _26177_ (.B1(_12564_),
    .Y(_12565_),
    .A1(net5926),
    .A2(net6205));
 sg13g2_nand2_1 _26178_ (.Y(_12566_),
    .A(_00865_),
    .B(net6205));
 sg13g2_o21ai_1 _26179_ (.B1(_12566_),
    .Y(_12567_),
    .A1(_10822_),
    .A2(net6205));
 sg13g2_nand2_1 _26180_ (.Y(_12568_),
    .A(_00864_),
    .B(net6206));
 sg13g2_o21ai_1 _26181_ (.B1(_12568_),
    .Y(_12569_),
    .A1(net6015),
    .A2(net6206));
 sg13g2_nand2_1 _26182_ (.Y(_12570_),
    .A(_00863_),
    .B(net6207));
 sg13g2_o21ai_1 _26183_ (.B1(_12570_),
    .Y(_12571_),
    .A1(net5961),
    .A2(net5981));
 sg13g2_nand2_1 _26184_ (.Y(_12572_),
    .A(_00862_),
    .B(net6264));
 sg13g2_o21ai_1 _26185_ (.B1(_12572_),
    .Y(_12573_),
    .A1(net5864),
    .A2(net6095));
 sg13g2_nand2_1 _26186_ (.Y(_12574_),
    .A(_00861_),
    .B(net6206));
 sg13g2_o21ai_1 _26187_ (.B1(_12574_),
    .Y(_12575_),
    .A1(net6011),
    .A2(net6206));
 sg13g2_mux2_1 _26188_ (.A0(_01349_),
    .A1(_01384_),
    .S(net7793),
    .X(_12576_));
 sg13g2_nand2_1 _26189_ (.Y(_12577_),
    .A(_00860_),
    .B(net6204));
 sg13g2_o21ai_1 _26190_ (.B1(_12577_),
    .Y(_12578_),
    .A1(net6001),
    .A2(net6204));
 sg13g2_nand2_1 _26191_ (.Y(_12579_),
    .A(_00859_),
    .B(net6201));
 sg13g2_nor3_1 _26192_ (.A(net7573),
    .B(net7558),
    .C(_12576_),
    .Y(_12580_));
 sg13g2_o21ai_1 _26193_ (.B1(_12579_),
    .Y(_12581_),
    .A1(net6118),
    .A2(net6201));
 sg13g2_nand2_1 _26194_ (.Y(_12582_),
    .A(_00858_),
    .B(net6205));
 sg13g2_o21ai_1 _26195_ (.B1(_12582_),
    .Y(_12583_),
    .A1(net6032),
    .A2(net6205));
 sg13g2_nand2_1 _26196_ (.Y(_12584_),
    .A(_00857_),
    .B(net6201));
 sg13g2_o21ai_1 _26197_ (.B1(_12584_),
    .Y(_12585_),
    .A1(net6112),
    .A2(net6201));
 sg13g2_nand2_1 _26198_ (.Y(_12586_),
    .A(_00856_),
    .B(net6201));
 sg13g2_o21ai_1 _26199_ (.B1(_12586_),
    .Y(_12587_),
    .A1(net6023),
    .A2(net6201));
 sg13g2_nand2_1 _26200_ (.Y(_12588_),
    .A(_00855_),
    .B(net6204));
 sg13g2_o21ai_1 _26201_ (.B1(_12588_),
    .Y(_12589_),
    .A1(net6051),
    .A2(net6208));
 sg13g2_nand2_1 _26202_ (.Y(_12590_),
    .A(_00854_),
    .B(net6206));
 sg13g2_o21ai_1 _26203_ (.B1(_12590_),
    .Y(_12591_),
    .A1(net6021),
    .A2(net6206));
 sg13g2_nand2_1 _26204_ (.Y(_12592_),
    .A(_00853_),
    .B(net6204));
 sg13g2_o21ai_1 _26205_ (.B1(_12592_),
    .Y(_12593_),
    .A1(net6107),
    .A2(net6204));
 sg13g2_nand2_1 _26206_ (.Y(_12594_),
    .A(_00852_),
    .B(net6207));
 sg13g2_o21ai_1 _26207_ (.B1(_12594_),
    .Y(_12595_),
    .A1(net5865),
    .A2(net5981));
 sg13g2_or4_1 _26208_ (.A(net7667),
    .B(net6468),
    .C(_09606_),
    .D(_11159_),
    .X(_12596_));
 sg13g2_nand2_1 _26209_ (.Y(_12597_),
    .A(net7447),
    .B(_11799_));
 sg13g2_nand2_1 _26210_ (.Y(_12598_),
    .A(_00851_),
    .B(net6200));
 sg13g2_o21ai_1 _26211_ (.B1(_12598_),
    .Y(_12599_),
    .A1(net5861),
    .A2(net6200));
 sg13g2_nand2_1 _26212_ (.Y(_12600_),
    .A(_00850_),
    .B(net6200));
 sg13g2_nand2b_1 _26213_ (.Y(_12601_),
    .B(net6381),
    .A_N(net6200));
 sg13g2_o21ai_1 _26214_ (.B1(_12600_),
    .Y(_12602_),
    .A1(net5855),
    .A2(_12601_));
 sg13g2_mux2_1 _26215_ (.A0(_01490_),
    .A1(_01525_),
    .S(net7793),
    .X(_12603_));
 sg13g2_nand2_1 _26216_ (.Y(_12604_),
    .A(_00849_),
    .B(net6194));
 sg13g2_o21ai_1 _26217_ (.B1(_12604_),
    .Y(_12605_),
    .A1(net5809),
    .A2(net6071));
 sg13g2_nand2_1 _26218_ (.Y(_12606_),
    .A(_00848_),
    .B(net6199));
 sg13g2_nor3_1 _26219_ (.A(net7573),
    .B(net7562),
    .C(_12603_),
    .Y(_12607_));
 sg13g2_o21ai_1 _26220_ (.B1(_12606_),
    .Y(_12608_),
    .A1(net5848),
    .A2(net6199));
 sg13g2_nand2_1 _26221_ (.Y(_12609_),
    .A(_00847_),
    .B(net6198));
 sg13g2_o21ai_1 _26222_ (.B1(_12609_),
    .Y(_12610_),
    .A1(net5799),
    .A2(net6198));
 sg13g2_nand2_1 _26223_ (.Y(_12611_),
    .A(_00846_),
    .B(net6197));
 sg13g2_o21ai_1 _26224_ (.B1(_12611_),
    .Y(_12612_),
    .A1(net5794),
    .A2(_12597_));
 sg13g2_nand2_1 _26225_ (.Y(_12613_),
    .A(_00845_),
    .B(_12596_));
 sg13g2_nand2b_1 _26226_ (.Y(_12614_),
    .B(net6378),
    .A_N(_12596_));
 sg13g2_o21ai_1 _26227_ (.B1(_12613_),
    .Y(_12615_),
    .A1(net5917),
    .A2(_12614_));
 sg13g2_nand2_1 _26228_ (.Y(_12616_),
    .A(_00844_),
    .B(net6194));
 sg13g2_o21ai_1 _26229_ (.B1(_12616_),
    .Y(_12617_),
    .A1(net5787),
    .A2(_12597_));
 sg13g2_nand2_1 _26230_ (.Y(_12618_),
    .A(_00843_),
    .B(net6200));
 sg13g2_nand2b_1 _26231_ (.Y(_12619_),
    .B(net6375),
    .A_N(_12596_));
 sg13g2_o21ai_1 _26232_ (.B1(_12618_),
    .Y(_12620_),
    .A1(net5912),
    .A2(_12619_));
 sg13g2_nand2_1 _26233_ (.Y(_12621_),
    .A(_00842_),
    .B(net6194));
 sg13g2_o21ai_1 _26234_ (.B1(_12621_),
    .Y(_12622_),
    .A1(net5782),
    .A2(net6071));
 sg13g2_nand2_1 _26235_ (.Y(_12623_),
    .A(_00841_),
    .B(_12596_));
 sg13g2_nand2b_1 _26236_ (.Y(_12624_),
    .B(net6368),
    .A_N(_12596_));
 sg13g2_o21ai_1 _26237_ (.B1(_12623_),
    .Y(_12625_),
    .A1(net5911),
    .A2(_12624_));
 sg13g2_mux2_1 _26238_ (.A0(net5840),
    .A1(_00840_),
    .S(_12597_),
    .X(_12626_));
 sg13g2_nand2_1 _26239_ (.Y(_12627_),
    .A(_00839_),
    .B(net6194));
 sg13g2_o21ai_1 _26240_ (.B1(_12627_),
    .Y(_12628_),
    .A1(net5837),
    .A2(_12597_));
 sg13g2_nand2_1 _26241_ (.Y(_12629_),
    .A(_00838_),
    .B(net6194));
 sg13g2_o21ai_1 _26242_ (.B1(_12629_),
    .Y(_12630_),
    .A1(net5903),
    .A2(_12597_));
 sg13g2_mux2_1 _26243_ (.A0(_01419_),
    .A1(_01454_),
    .S(net7793),
    .X(_12631_));
 sg13g2_nand2_1 _26244_ (.Y(_12632_),
    .A(_00837_),
    .B(net6194));
 sg13g2_o21ai_1 _26245_ (.B1(_12632_),
    .Y(_12633_),
    .A1(net5899),
    .A2(net6071));
 sg13g2_nand2_1 _26246_ (.Y(_12634_),
    .A(_00836_),
    .B(net6197));
 sg13g2_nor3_1 _26247_ (.A(net7573),
    .B(net7571),
    .C(_12631_),
    .Y(_12635_));
 sg13g2_o21ai_1 _26248_ (.B1(_12634_),
    .Y(_12636_),
    .A1(net5889),
    .A2(net6197));
 sg13g2_mux2_1 _26249_ (.A0(net5773),
    .A1(_00835_),
    .S(_12596_),
    .X(_12637_));
 sg13g2_nand2_1 _26250_ (.Y(_12638_),
    .A(_00834_),
    .B(net6197));
 sg13g2_o21ai_1 _26251_ (.B1(_12638_),
    .Y(_12639_),
    .A1(net5884),
    .A2(net6195));
 sg13g2_nand2_1 _26252_ (.Y(_12640_),
    .A(_00833_),
    .B(net6198));
 sg13g2_o21ai_1 _26253_ (.B1(_12640_),
    .Y(_12641_),
    .A1(net5926),
    .A2(net6198));
 sg13g2_nand2_1 _26254_ (.Y(_12642_),
    .A(_00832_),
    .B(net6196));
 sg13g2_o21ai_1 _26255_ (.B1(_12642_),
    .Y(_12643_),
    .A1(net5964),
    .A2(net6196));
 sg13g2_nand2_1 _26256_ (.Y(_12644_),
    .A(_00831_),
    .B(net6196));
 sg13g2_o21ai_1 _26257_ (.B1(_12644_),
    .Y(_12645_),
    .A1(net6015),
    .A2(net6196));
 sg13g2_nand2_1 _26258_ (.Y(_12646_),
    .A(_00830_),
    .B(net6194));
 sg13g2_o21ai_1 _26259_ (.B1(_12646_),
    .Y(_12647_),
    .A1(net5959),
    .A2(_12597_));
 sg13g2_nand2_1 _26260_ (.Y(_12648_),
    .A(_00829_),
    .B(net6196));
 sg13g2_o21ai_1 _26261_ (.B1(_12648_),
    .Y(_12649_),
    .A1(net6011),
    .A2(net6196));
 sg13g2_nand2_1 _26262_ (.Y(_12650_),
    .A(_00828_),
    .B(net6195));
 sg13g2_o21ai_1 _26263_ (.B1(_12650_),
    .Y(_12651_),
    .A1(net6001),
    .A2(net6195));
 sg13g2_nand2_1 _26264_ (.Y(_12652_),
    .A(_00827_),
    .B(net6199));
 sg13g2_o21ai_1 _26265_ (.B1(_12652_),
    .Y(_12653_),
    .A1(net6118),
    .A2(net6199));
 sg13g2_nand2_1 _26266_ (.Y(_12654_),
    .A(_00826_),
    .B(net6196));
 sg13g2_mux2_1 _26267_ (.A0(_01560_),
    .A1(_01595_),
    .S(net7793),
    .X(_12655_));
 sg13g2_o21ai_1 _26268_ (.B1(_12654_),
    .Y(_12656_),
    .A1(net6032),
    .A2(net6196));
 sg13g2_nand2_1 _26269_ (.Y(_12657_),
    .A(_00825_),
    .B(net6199));
 sg13g2_o21ai_1 _26270_ (.B1(_12657_),
    .Y(_12658_),
    .A1(net6114),
    .A2(net6199));
 sg13g2_nor2_1 _26271_ (.A(net7555),
    .B(_12655_),
    .Y(_12659_));
 sg13g2_nand2_1 _26272_ (.Y(_12660_),
    .A(_00824_),
    .B(net6199));
 sg13g2_o21ai_1 _26273_ (.B1(_12660_),
    .Y(_12661_),
    .A1(net6023),
    .A2(net6199));
 sg13g2_nand2_1 _26274_ (.Y(_12662_),
    .A(_00823_),
    .B(net6195));
 sg13g2_o21ai_1 _26275_ (.B1(_12662_),
    .Y(_12663_),
    .A1(net6055),
    .A2(net6195));
 sg13g2_nand2_1 _26276_ (.Y(_12664_),
    .A(_00822_),
    .B(net6195));
 sg13g2_o21ai_1 _26277_ (.B1(_12664_),
    .Y(_12665_),
    .A1(net6020),
    .A2(net6197));
 sg13g2_nand2_1 _26278_ (.Y(_12666_),
    .A(_00821_),
    .B(net6195));
 sg13g2_o21ai_1 _26279_ (.B1(_12666_),
    .Y(_12667_),
    .A1(net6107),
    .A2(net6195));
 sg13g2_nand2_1 _26280_ (.Y(_12668_),
    .A(_00820_),
    .B(net6194));
 sg13g2_or4_1 _26281_ (.A(_12580_),
    .B(_12607_),
    .C(_12635_),
    .D(_12659_),
    .X(_12669_));
 sg13g2_o21ai_1 _26282_ (.B1(_12668_),
    .Y(_12670_),
    .A1(net5865),
    .A2(net6071));
 sg13g2_or4_1 _26283_ (.A(net7667),
    .B(_06622_),
    .C(net6468),
    .D(_11159_),
    .X(_12671_));
 sg13g2_nand3_1 _26284_ (.B(_10990_),
    .C(net7447),
    .A(_06621_),
    .Y(_12672_));
 sg13g2_nand2_1 _26285_ (.Y(_12673_),
    .A(_00819_),
    .B(net6187));
 sg13g2_o21ai_1 _26286_ (.B1(_12673_),
    .Y(_12674_),
    .A1(net5861),
    .A2(net6187));
 sg13g2_nand2_1 _26287_ (.Y(_12675_),
    .A(_00818_),
    .B(net6187));
 sg13g2_nand2b_1 _26288_ (.Y(_12676_),
    .B(net6381),
    .A_N(net6189));
 sg13g2_o21ai_1 _26289_ (.B1(_12675_),
    .Y(_12677_),
    .A1(net5855),
    .A2(_12676_));
 sg13g2_nand2_1 _26290_ (.Y(_12678_),
    .A(_00817_),
    .B(net6190));
 sg13g2_o21ai_1 _26291_ (.B1(_12678_),
    .Y(_12679_),
    .A1(net5809),
    .A2(net6070));
 sg13g2_nand2_1 _26292_ (.Y(_12680_),
    .A(_00816_),
    .B(net6188));
 sg13g2_o21ai_1 _26293_ (.B1(_12680_),
    .Y(_12681_),
    .A1(net5848),
    .A2(net6188));
 sg13g2_nand2_1 _26294_ (.Y(_12682_),
    .A(_00815_),
    .B(net6188));
 sg13g2_o21ai_1 _26295_ (.B1(_12682_),
    .Y(_12683_),
    .A1(net5798),
    .A2(net6188));
 sg13g2_nand2_1 _26296_ (.Y(_12684_),
    .A(_00814_),
    .B(net6193));
 sg13g2_o21ai_1 _26297_ (.B1(_12684_),
    .Y(_12685_),
    .A1(net5794),
    .A2(net6070));
 sg13g2_nand2_1 _26298_ (.Y(_12686_),
    .A(_00813_),
    .B(net6186));
 sg13g2_nand2b_1 _26299_ (.Y(_12687_),
    .B(net6378),
    .A_N(net6186));
 sg13g2_o21ai_1 _26300_ (.B1(_12686_),
    .Y(_12688_),
    .A1(net5917),
    .A2(_12687_));
 sg13g2_nand2_1 _26301_ (.Y(_12689_),
    .A(_00812_),
    .B(net6190));
 sg13g2_o21ai_1 _26302_ (.B1(_12689_),
    .Y(_12690_),
    .A1(net5787),
    .A2(net6070));
 sg13g2_nand2_1 _26303_ (.Y(_12691_),
    .A(_00811_),
    .B(net6189));
 sg13g2_nand2b_1 _26304_ (.Y(_12692_),
    .B(net6374),
    .A_N(_12671_));
 sg13g2_o21ai_1 _26305_ (.B1(_12691_),
    .Y(_12693_),
    .A1(net5912),
    .A2(_12692_));
 sg13g2_nand2_1 _26306_ (.Y(_12694_),
    .A(_00810_),
    .B(net6190));
 sg13g2_o21ai_1 _26307_ (.B1(_12694_),
    .Y(_12695_),
    .A1(net5782),
    .A2(net6070));
 sg13g2_nand2_1 _26308_ (.Y(_12696_),
    .A(_00809_),
    .B(net6186));
 sg13g2_nand2b_1 _26309_ (.Y(_12697_),
    .B(net6368),
    .A_N(_12671_));
 sg13g2_o21ai_1 _26310_ (.B1(_12696_),
    .Y(_12698_),
    .A1(net5909),
    .A2(_12697_));
 sg13g2_mux4_1 _26311_ (.S0(net7791),
    .A0(_01208_),
    .A1(_01243_),
    .A2(_01278_),
    .A3(_01314_),
    .S1(net7741),
    .X(_12699_));
 sg13g2_mux2_1 _26312_ (.A0(net5839),
    .A1(_00808_),
    .S(_12672_),
    .X(_12700_));
 sg13g2_nand2_1 _26313_ (.Y(_12701_),
    .A(_00807_),
    .B(net6190));
 sg13g2_o21ai_1 _26314_ (.B1(_12701_),
    .Y(_12702_),
    .A1(net5834),
    .A2(net6070));
 sg13g2_nand2_1 _26315_ (.Y(_12703_),
    .A(_00806_),
    .B(net6190));
 sg13g2_o21ai_1 _26316_ (.B1(_12703_),
    .Y(_12704_),
    .A1(net5903),
    .A2(net6070));
 sg13g2_nand2_1 _26317_ (.Y(_12705_),
    .A(_00805_),
    .B(net6190));
 sg13g2_o21ai_1 _26318_ (.B1(_12705_),
    .Y(_12706_),
    .A1(net5899),
    .A2(net6070));
 sg13g2_nand2_1 _26319_ (.Y(_12707_),
    .A(_00804_),
    .B(net6193));
 sg13g2_o21ai_1 _26320_ (.B1(_12707_),
    .Y(_12708_),
    .A1(net5889),
    .A2(net6193));
 sg13g2_mux2_1 _26321_ (.A0(net5772),
    .A1(_00803_),
    .S(_12671_),
    .X(_12709_));
 sg13g2_nand2_1 _26322_ (.Y(_12710_),
    .A(_00802_),
    .B(net6191));
 sg13g2_o21ai_1 _26323_ (.B1(_12710_),
    .Y(_12711_),
    .A1(net5884),
    .A2(net6191));
 sg13g2_nand2_1 _26324_ (.Y(_12712_),
    .A(_00801_),
    .B(net6188));
 sg13g2_o21ai_1 _26325_ (.B1(_12712_),
    .Y(_12713_),
    .A1(net5926),
    .A2(net6188));
 sg13g2_nand2_1 _26326_ (.Y(_12714_),
    .A(_00800_),
    .B(net6192));
 sg13g2_o21ai_1 _26327_ (.B1(_12714_),
    .Y(_12715_),
    .A1(net5964),
    .A2(net6192));
 sg13g2_nand2_1 _26328_ (.Y(_12716_),
    .A(_00799_),
    .B(net6192));
 sg13g2_o21ai_1 _26329_ (.B1(_12716_),
    .Y(_12717_),
    .A1(net6015),
    .A2(net6192));
 sg13g2_nand2_1 _26330_ (.Y(_12718_),
    .A(_00798_),
    .B(net6190));
 sg13g2_o21ai_1 _26331_ (.B1(_12718_),
    .Y(_12719_),
    .A1(net5959),
    .A2(_12672_));
 sg13g2_nand2_1 _26332_ (.Y(_12720_),
    .A(_00797_),
    .B(net6192));
 sg13g2_o21ai_1 _26333_ (.B1(_12720_),
    .Y(_12721_),
    .A1(net6011),
    .A2(net6192));
 sg13g2_nand2_1 _26334_ (.Y(_12722_),
    .A(_00796_),
    .B(net6191));
 sg13g2_o21ai_1 _26335_ (.B1(_12722_),
    .Y(_12723_),
    .A1(net6001),
    .A2(net6191));
 sg13g2_nand2_1 _26336_ (.Y(_12724_),
    .A(_00795_),
    .B(net6189));
 sg13g2_o21ai_1 _26337_ (.B1(_12724_),
    .Y(_12725_),
    .A1(net6118),
    .A2(net6189));
 sg13g2_nand2_1 _26338_ (.Y(_12726_),
    .A(_00794_),
    .B(net6192));
 sg13g2_o21ai_1 _26339_ (.B1(_12726_),
    .Y(_12727_),
    .A1(net6031),
    .A2(net6192));
 sg13g2_nand2_1 _26340_ (.Y(_12728_),
    .A(_00793_),
    .B(net6187));
 sg13g2_o21ai_1 _26341_ (.B1(_12728_),
    .Y(_12729_),
    .A1(net6112),
    .A2(net6187));
 sg13g2_nand2_1 _26342_ (.Y(_12730_),
    .A(_00792_),
    .B(net6189));
 sg13g2_mux4_1 _26343_ (.S0(net7791),
    .A0(_01067_),
    .A1(_01102_),
    .A2(_01138_),
    .A3(_01173_),
    .S1(net7741),
    .X(_12731_));
 sg13g2_o21ai_1 _26344_ (.B1(_12730_),
    .Y(_12732_),
    .A1(net6023),
    .A2(net6189));
 sg13g2_nand2_1 _26345_ (.Y(_12733_),
    .A(_00791_),
    .B(net6191));
 sg13g2_o21ai_1 _26346_ (.B1(_12733_),
    .Y(_12734_),
    .A1(net6051),
    .A2(net6191));
 sg13g2_nor2b_1 _26347_ (.A(net7709),
    .B_N(_12731_),
    .Y(_12735_));
 sg13g2_nand2_1 _26348_ (.Y(_12736_),
    .A(_00790_),
    .B(net6193));
 sg13g2_o21ai_1 _26349_ (.B1(_12736_),
    .Y(_12737_),
    .A1(net6022),
    .A2(net6193));
 sg13g2_nand2_1 _26350_ (.Y(_12738_),
    .A(_00789_),
    .B(net6191));
 sg13g2_o21ai_1 _26351_ (.B1(_12738_),
    .Y(_12739_),
    .A1(net6107),
    .A2(net6191));
 sg13g2_nand2_1 _26352_ (.Y(_12740_),
    .A(_00788_),
    .B(net6190));
 sg13g2_o21ai_1 _26353_ (.B1(_12740_),
    .Y(_12741_),
    .A1(_10088_),
    .A2(_12672_));
 sg13g2_nor2_1 _26354_ (.A(_09609_),
    .B(_11478_),
    .Y(_12742_));
 sg13g2_nand2_1 _26355_ (.Y(_12743_),
    .A(_09608_),
    .B(net7446));
 sg13g2_nand2_1 _26356_ (.Y(_12744_),
    .A(_00787_),
    .B(net5976));
 sg13g2_o21ai_1 _26357_ (.B1(_12744_),
    .Y(_12745_),
    .A1(net8286),
    .A2(net5976));
 sg13g2_nand2_1 _26358_ (.Y(_12746_),
    .A(net6382),
    .B(_12742_));
 sg13g2_nand2_1 _26359_ (.Y(_12747_),
    .A(_00786_),
    .B(net5976));
 sg13g2_o21ai_1 _26360_ (.B1(_12747_),
    .Y(_12748_),
    .A1(net5853),
    .A2(_12746_));
 sg13g2_nand2_1 _26361_ (.Y(_12749_),
    .A(_00785_),
    .B(net5980));
 sg13g2_o21ai_1 _26362_ (.B1(_12749_),
    .Y(_12750_),
    .A1(net5804),
    .A2(net5980));
 sg13g2_nand2_1 _26363_ (.Y(_12751_),
    .A(_00784_),
    .B(net5978));
 sg13g2_o21ai_1 _26364_ (.B1(_12751_),
    .Y(_12752_),
    .A1(net5847),
    .A2(net5978));
 sg13g2_nand2_1 _26365_ (.Y(_12753_),
    .A(_00783_),
    .B(net5977));
 sg13g2_o21ai_1 _26366_ (.B1(_12753_),
    .Y(_12754_),
    .A1(net5803),
    .A2(net5977));
 sg13g2_nand2_1 _26367_ (.Y(_12755_),
    .A(_00782_),
    .B(net5972));
 sg13g2_o21ai_1 _26368_ (.B1(_12755_),
    .Y(_12756_),
    .A1(net5792),
    .A2(net5972));
 sg13g2_nand2_1 _26369_ (.Y(_12757_),
    .A(net6377),
    .B(_12742_));
 sg13g2_nand2_1 _26370_ (.Y(_12758_),
    .A(_00781_),
    .B(net5976));
 sg13g2_o21ai_1 _26371_ (.B1(_12758_),
    .Y(_12759_),
    .A1(net5917),
    .A2(_12757_));
 sg13g2_nand2_1 _26372_ (.Y(_12760_),
    .A(_00780_),
    .B(net5972));
 sg13g2_o21ai_1 _26373_ (.B1(_12760_),
    .Y(_12761_),
    .A1(net5786),
    .A2(net5972));
 sg13g2_nand2_1 _26374_ (.Y(_12762_),
    .A(net6370),
    .B(_12742_));
 sg13g2_nand2_1 _26375_ (.Y(_12763_),
    .A(_00779_),
    .B(net5976));
 sg13g2_o21ai_1 _26376_ (.B1(_12763_),
    .Y(_12764_),
    .A1(net5915),
    .A2(_12762_));
 sg13g2_nand2_1 _26377_ (.Y(_12765_),
    .A(_00778_),
    .B(net5980));
 sg13g2_o21ai_1 _26378_ (.B1(_12765_),
    .Y(_12766_),
    .A1(net5783),
    .A2(net5980));
 sg13g2_nand2_1 _26379_ (.Y(_12767_),
    .A(net6365),
    .B(_12742_));
 sg13g2_nand2_1 _26380_ (.Y(_12768_),
    .A(_00777_),
    .B(net5976));
 sg13g2_o21ai_1 _26381_ (.B1(_12768_),
    .Y(_12769_),
    .A1(net5908),
    .A2(_12767_));
 sg13g2_mux2_1 _26382_ (.A0(_00776_),
    .A1(net5838),
    .S(_12742_),
    .X(_12770_));
 sg13g2_nand2_1 _26383_ (.Y(_12771_),
    .A(_00775_),
    .B(net5972));
 sg13g2_o21ai_1 _26384_ (.B1(_12771_),
    .Y(_12772_),
    .A1(net5836),
    .A2(net5972));
 sg13g2_a21oi_1 _26385_ (.A1(net7709),
    .A2(_12699_),
    .Y(_12773_),
    .B1(_12735_));
 sg13g2_nand2_1 _26386_ (.Y(_12774_),
    .A(_00774_),
    .B(_12743_));
 sg13g2_o21ai_1 _26387_ (.B1(_12774_),
    .Y(_12775_),
    .A1(net5902),
    .A2(_12743_));
 sg13g2_nand2_1 _26388_ (.Y(_12776_),
    .A(_00773_),
    .B(net5980));
 sg13g2_o21ai_1 _26389_ (.B1(_12776_),
    .Y(_12777_),
    .A1(net5897),
    .A2(net5980));
 sg13g2_nand2_1 _26390_ (.Y(_12778_),
    .A(_00772_),
    .B(net5972));
 sg13g2_o21ai_1 _26391_ (.B1(_12778_),
    .Y(_12779_),
    .A1(net5888),
    .A2(net5979));
 sg13g2_mux2_1 _26392_ (.A0(_00771_),
    .A1(net5772),
    .S(_12742_),
    .X(_12780_));
 sg13g2_a21oi_1 _26393_ (.A1(net7592),
    .A2(_12773_),
    .Y(_12781_),
    .B1(_12669_));
 sg13g2_nand2_1 _26394_ (.Y(_12782_),
    .A(_00770_),
    .B(net5973));
 sg13g2_o21ai_1 _26395_ (.B1(_12782_),
    .Y(_12783_),
    .A1(net5885),
    .A2(net5973));
 sg13g2_nand2_1 _26396_ (.Y(_12784_),
    .A(_00769_),
    .B(net5977));
 sg13g2_o21ai_1 _26397_ (.B1(_12784_),
    .Y(_12785_),
    .A1(net5929),
    .A2(net5977));
 sg13g2_nand2_1 _26398_ (.Y(_12786_),
    .A(_00768_),
    .B(net5975));
 sg13g2_o21ai_1 _26399_ (.B1(_12786_),
    .Y(_12787_),
    .A1(net5962),
    .A2(net5975));
 sg13g2_a221oi_1 _26400_ (.B2(net7592),
    .C1(_12669_),
    .B1(_12773_),
    .A1(_12429_),
    .Y(_12788_),
    .A2(_12553_));
 sg13g2_nand2_1 _26401_ (.Y(_12789_),
    .A(_00767_),
    .B(net5975));
 sg13g2_o21ai_1 _26402_ (.B1(_12789_),
    .Y(_12790_),
    .A1(net6014),
    .A2(net5975));
 sg13g2_nand2_1 _26403_ (.Y(_12791_),
    .A(_12558_),
    .B(_12781_));
 sg13g2_nand2_1 _26404_ (.Y(_12792_),
    .A(_00766_),
    .B(_12743_));
 sg13g2_o21ai_1 _26405_ (.B1(_12792_),
    .Y(_12793_),
    .A1(net5957),
    .A2(_12743_));
 sg13g2_nand2_1 _26406_ (.Y(_12794_),
    .A(_00765_),
    .B(net5975));
 sg13g2_o21ai_1 _26407_ (.B1(_12794_),
    .Y(_12795_),
    .A1(net6010),
    .A2(net5975));
 sg13g2_nor2_1 _26408_ (.A(_08616_),
    .B(net7281),
    .Y(_12796_));
 sg13g2_nand2_1 _26409_ (.Y(_12797_),
    .A(_00764_),
    .B(net5974));
 sg13g2_o21ai_1 _26410_ (.B1(_12797_),
    .Y(_12798_),
    .A1(net6006),
    .A2(net5974));
 sg13g2_nand2_1 _26411_ (.Y(_12799_),
    .A(_00763_),
    .B(net5978));
 sg13g2_o21ai_1 _26412_ (.B1(_12799_),
    .Y(_12800_),
    .A1(net6117),
    .A2(net5978));
 sg13g2_nand2_1 _26413_ (.Y(_12801_),
    .A(_00762_),
    .B(net5975));
 sg13g2_o21ai_1 _26414_ (.B1(_12801_),
    .Y(_12802_),
    .A1(net6033),
    .A2(net5975));
 sg13g2_nand2_1 _26415_ (.Y(_12803_),
    .A(_00761_),
    .B(net5977));
 sg13g2_o21ai_1 _26416_ (.B1(_12803_),
    .Y(_12804_),
    .A1(net6114),
    .A2(net5977));
 sg13g2_nand2_1 _26417_ (.Y(_12805_),
    .A(_00760_),
    .B(net5978));
 sg13g2_o21ai_1 _26418_ (.B1(_12805_),
    .Y(_12806_),
    .A1(_09902_),
    .A2(net5978));
 sg13g2_nand2_1 _26419_ (.Y(_12807_),
    .A(_00759_),
    .B(net5973));
 sg13g2_o21ai_1 _26420_ (.B1(_12807_),
    .Y(_12808_),
    .A1(net6055),
    .A2(net5973));
 sg13g2_nand2_1 _26421_ (.Y(_12809_),
    .A(_00758_),
    .B(net5973));
 sg13g2_o21ai_1 _26422_ (.B1(_12809_),
    .Y(_12810_),
    .A1(net6022),
    .A2(net5973));
 sg13g2_nand2_1 _26423_ (.Y(_12811_),
    .A(_00757_),
    .B(net5973));
 sg13g2_o21ai_1 _26424_ (.B1(_12811_),
    .Y(_12812_),
    .A1(net6108),
    .A2(net5973));
 sg13g2_nand2_1 _26425_ (.Y(_12813_),
    .A(_00756_),
    .B(net5980));
 sg13g2_o21ai_1 _26426_ (.B1(_12813_),
    .Y(_12814_),
    .A1(net5864),
    .A2(net5980));
 sg13g2_nand4_1 _26427_ (.B(_06621_),
    .C(_09604_),
    .A(net7670),
    .Y(_12815_),
    .D(_11477_));
 sg13g2_nand2_1 _26428_ (.Y(_12816_),
    .A(_10985_),
    .B(net7446));
 sg13g2_nand2_1 _26429_ (.Y(_12817_),
    .A(_00755_),
    .B(net6184));
 sg13g2_o21ai_1 _26430_ (.B1(_12817_),
    .Y(_12818_),
    .A1(net5861),
    .A2(net6184));
 sg13g2_nor3_1 _26431_ (.A(net7360),
    .B(_12331_),
    .C(_12796_),
    .Y(_12819_));
 sg13g2_nand2_1 _26432_ (.Y(_12820_),
    .A(_00754_),
    .B(net6184));
 sg13g2_nand2b_1 _26433_ (.Y(_12821_),
    .B(net6382),
    .A_N(net6184));
 sg13g2_or3_1 _26434_ (.A(net7360),
    .B(_12331_),
    .C(_12796_),
    .X(_12822_));
 sg13g2_o21ai_1 _26435_ (.B1(_12820_),
    .Y(_12823_),
    .A1(net5858),
    .A2(_12821_));
 sg13g2_nand2_1 _26436_ (.Y(_12824_),
    .A(_00753_),
    .B(net6177));
 sg13g2_o21ai_1 _26437_ (.B1(_12824_),
    .Y(_12825_),
    .A1(net5804),
    .A2(net5971));
 sg13g2_nand2_1 _26438_ (.Y(_12826_),
    .A(_00752_),
    .B(net6183));
 sg13g2_o21ai_1 _26439_ (.B1(_12826_),
    .Y(_12827_),
    .A1(net5847),
    .A2(net6183));
 sg13g2_nand2_1 _26440_ (.Y(_12828_),
    .A(_00751_),
    .B(net6182));
 sg13g2_o21ai_1 _26441_ (.B1(_12828_),
    .Y(_12829_),
    .A1(net5803),
    .A2(net6182));
 sg13g2_nand2_1 _26442_ (.Y(_12830_),
    .A(_00750_),
    .B(_12815_));
 sg13g2_o21ai_1 _26443_ (.B1(_12830_),
    .Y(_12831_),
    .A1(net5792),
    .A2(net5971));
 sg13g2_nand2_1 _26444_ (.Y(_12832_),
    .A(_00749_),
    .B(net6184));
 sg13g2_nand2b_1 _26445_ (.Y(_12833_),
    .B(net6378),
    .A_N(net6185));
 sg13g2_o21ai_1 _26446_ (.B1(_12832_),
    .Y(_12834_),
    .A1(net5920),
    .A2(_12833_));
 sg13g2_nand2_1 _26447_ (.Y(_12835_),
    .A(_00748_),
    .B(_12815_));
 sg13g2_o21ai_1 _26448_ (.B1(_12835_),
    .Y(_12836_),
    .A1(net5786),
    .A2(net5971));
 sg13g2_nand2b_1 _26449_ (.Y(_12837_),
    .B(net6369),
    .A_N(net6178));
 sg13g2_nand2_1 _26450_ (.Y(_12838_),
    .A(_00747_),
    .B(net6178));
 sg13g2_o21ai_1 _26451_ (.B1(_12838_),
    .Y(_12839_),
    .A1(net5915),
    .A2(_12837_));
 sg13g2_nand2_1 _26452_ (.Y(_12840_),
    .A(_00746_),
    .B(net6177));
 sg13g2_o21ai_1 _26453_ (.B1(_12840_),
    .Y(_12841_),
    .A1(net5783),
    .A2(net5971));
 sg13g2_nand2b_1 _26454_ (.Y(_12842_),
    .B(net6364),
    .A_N(net6178));
 sg13g2_nand2_1 _26455_ (.Y(_12843_),
    .A(_00745_),
    .B(net6178));
 sg13g2_o21ai_1 _26456_ (.B1(_12843_),
    .Y(_12844_),
    .A1(net5907),
    .A2(_12842_));
 sg13g2_mux2_1 _26457_ (.A0(net5838),
    .A1(_00744_),
    .S(_12816_),
    .X(_12845_));
 sg13g2_nand2_1 _26458_ (.Y(_12846_),
    .A(_00743_),
    .B(_12815_));
 sg13g2_nand2_1 _26459_ (.Y(_12847_),
    .A(net7883),
    .B(_01595_));
 sg13g2_o21ai_1 _26460_ (.B1(_12846_),
    .Y(_12848_),
    .A1(net5836),
    .A2(net5971));
 sg13g2_nand2_1 _26461_ (.Y(_12849_),
    .A(_00742_),
    .B(net6177));
 sg13g2_o21ai_1 _26462_ (.B1(_12849_),
    .Y(_12850_),
    .A1(net5902),
    .A2(net5971));
 sg13g2_nand2b_1 _26463_ (.Y(_12851_),
    .B(_01560_),
    .A_N(net7883));
 sg13g2_nand2_1 _26464_ (.Y(_12852_),
    .A(_00741_),
    .B(net6177));
 sg13g2_o21ai_1 _26465_ (.B1(_12852_),
    .Y(_12853_),
    .A1(net5897),
    .A2(net5971));
 sg13g2_nand2_1 _26466_ (.Y(_12854_),
    .A(_00740_),
    .B(net6179));
 sg13g2_o21ai_1 _26467_ (.B1(_12854_),
    .Y(_12855_),
    .A1(net5888),
    .A2(net6179));
 sg13g2_mux2_1 _26468_ (.A0(net5773),
    .A1(_00739_),
    .S(net6178),
    .X(_12856_));
 sg13g2_nand2_1 _26469_ (.Y(_12857_),
    .A(_00738_),
    .B(net6179));
 sg13g2_o21ai_1 _26470_ (.B1(_12857_),
    .Y(_12858_),
    .A1(net5885),
    .A2(net6179));
 sg13g2_nand2_1 _26471_ (.Y(_12859_),
    .A(_00737_),
    .B(net6182));
 sg13g2_o21ai_1 _26472_ (.B1(_12859_),
    .Y(_12860_),
    .A1(net5925),
    .A2(net6182));
 sg13g2_nand2_1 _26473_ (.Y(_12861_),
    .A(_00736_),
    .B(net6180));
 sg13g2_o21ai_1 _26474_ (.B1(_12861_),
    .Y(_12862_),
    .A1(net5962),
    .A2(net6180));
 sg13g2_nand2_1 _26475_ (.Y(_12863_),
    .A(_00735_),
    .B(net6180));
 sg13g2_o21ai_1 _26476_ (.B1(_12863_),
    .Y(_12864_),
    .A1(net6014),
    .A2(net6180));
 sg13g2_nand2_1 _26477_ (.Y(_12865_),
    .A(_00734_),
    .B(net6177));
 sg13g2_o21ai_1 _26478_ (.B1(_12865_),
    .Y(_12866_),
    .A1(net5957),
    .A2(_12816_));
 sg13g2_nand2_1 _26479_ (.Y(_12867_),
    .A(_00733_),
    .B(net6180));
 sg13g2_nand3_1 _26480_ (.B(_12847_),
    .C(_12851_),
    .A(net7450),
    .Y(_12868_));
 sg13g2_o21ai_1 _26481_ (.B1(_12867_),
    .Y(_12869_),
    .A1(net6010),
    .A2(net6180));
 sg13g2_nand2_1 _26482_ (.Y(_12870_),
    .A(_00732_),
    .B(net6181));
 sg13g2_o21ai_1 _26483_ (.B1(_12870_),
    .Y(_12871_),
    .A1(net6007),
    .A2(net6181));
 sg13g2_nand2_1 _26484_ (.Y(_12872_),
    .A(net7849),
    .B(_01525_));
 sg13g2_nand2_1 _26485_ (.Y(_12873_),
    .A(_00731_),
    .B(net6183));
 sg13g2_o21ai_1 _26486_ (.B1(_12873_),
    .Y(_12874_),
    .A1(net6117),
    .A2(net6183));
 sg13g2_nand2_1 _26487_ (.Y(_12875_),
    .A(_00730_),
    .B(net6180));
 sg13g2_nand2b_1 _26488_ (.Y(_12876_),
    .B(_01490_),
    .A_N(net7849));
 sg13g2_o21ai_1 _26489_ (.B1(_12875_),
    .Y(_12877_),
    .A1(net6033),
    .A2(net6180));
 sg13g2_nand2_1 _26490_ (.Y(_12878_),
    .A(_00729_),
    .B(net6183));
 sg13g2_o21ai_1 _26491_ (.B1(_12878_),
    .Y(_12879_),
    .A1(net6109),
    .A2(net6184));
 sg13g2_nand2_1 _26492_ (.Y(_12880_),
    .A(_00728_),
    .B(net6183));
 sg13g2_o21ai_1 _26493_ (.B1(_12880_),
    .Y(_12881_),
    .A1(_09902_),
    .A2(net6183));
 sg13g2_nand2_1 _26494_ (.Y(_12882_),
    .A(_00727_),
    .B(net6181));
 sg13g2_o21ai_1 _26495_ (.B1(_12882_),
    .Y(_12883_),
    .A1(net6055),
    .A2(net6179));
 sg13g2_nand2_1 _26496_ (.Y(_12884_),
    .A(_00726_),
    .B(net6181));
 sg13g2_o21ai_1 _26497_ (.B1(_12884_),
    .Y(_12885_),
    .A1(net6022),
    .A2(net6181));
 sg13g2_nand2_1 _26498_ (.Y(_12886_),
    .A(_00725_),
    .B(net6181));
 sg13g2_o21ai_1 _26499_ (.B1(_12886_),
    .Y(_12887_),
    .A1(net6108),
    .A2(net6179));
 sg13g2_nand2_1 _26500_ (.Y(_12888_),
    .A(_00724_),
    .B(net6177));
 sg13g2_o21ai_1 _26501_ (.B1(_12888_),
    .Y(_12889_),
    .A1(net5864),
    .A2(_12816_));
 sg13g2_or4_1 _26502_ (.A(net7667),
    .B(net6468),
    .C(_09606_),
    .D(_11478_),
    .X(_12890_));
 sg13g2_nand2_1 _26503_ (.Y(_12891_),
    .A(net7446),
    .B(_11799_));
 sg13g2_nand2_1 _26504_ (.Y(_12892_),
    .A(_00723_),
    .B(net6176));
 sg13g2_o21ai_1 _26505_ (.B1(_12892_),
    .Y(_12893_),
    .A1(net5861),
    .A2(net6176));
 sg13g2_nand2_1 _26506_ (.Y(_12894_),
    .A(_00722_),
    .B(net6176));
 sg13g2_nand4_1 _26507_ (.B(net7494),
    .C(_12872_),
    .A(net7512),
    .Y(_12895_),
    .D(_12876_));
 sg13g2_nand2b_1 _26508_ (.Y(_12896_),
    .B(net6381),
    .A_N(net6176));
 sg13g2_o21ai_1 _26509_ (.B1(_12894_),
    .Y(_12897_),
    .A1(net5855),
    .A2(_12896_));
 sg13g2_nand2_1 _26510_ (.Y(_12898_),
    .A(_00721_),
    .B(net6169));
 sg13g2_o21ai_1 _26511_ (.B1(_12898_),
    .Y(_12899_),
    .A1(net5804),
    .A2(net6069));
 sg13g2_nand2_1 _26512_ (.Y(_12900_),
    .A(_00720_),
    .B(net6174));
 sg13g2_o21ai_1 _26513_ (.B1(_12900_),
    .Y(_12901_),
    .A1(net5847),
    .A2(net6174));
 sg13g2_nand2_1 _26514_ (.Y(_12902_),
    .A(net7846),
    .B(_00824_));
 sg13g2_nand2_1 _26515_ (.Y(_12903_),
    .A(_00719_),
    .B(net6175));
 sg13g2_o21ai_1 _26516_ (.B1(_12903_),
    .Y(_12904_),
    .A1(net5798),
    .A2(net6172));
 sg13g2_nand2_1 _26517_ (.Y(_12905_),
    .A(_00718_),
    .B(_12890_));
 sg13g2_o21ai_1 _26518_ (.B1(_12905_),
    .Y(_12906_),
    .A1(net5792),
    .A2(net6069));
 sg13g2_nand2b_1 _26519_ (.Y(_12907_),
    .B(_00792_),
    .A_N(net7846));
 sg13g2_nand2_1 _26520_ (.Y(_12908_),
    .A(_00717_),
    .B(net6171));
 sg13g2_nand2b_1 _26521_ (.Y(_12909_),
    .B(net6378),
    .A_N(net6171));
 sg13g2_o21ai_1 _26522_ (.B1(_12908_),
    .Y(_12910_),
    .A1(net5920),
    .A2(_12909_));
 sg13g2_nand2_1 _26523_ (.Y(_12911_),
    .A(_00716_),
    .B(_12890_));
 sg13g2_o21ai_1 _26524_ (.B1(_12911_),
    .Y(_12912_),
    .A1(net5785),
    .A2(_12891_));
 sg13g2_nand2b_1 _26525_ (.Y(_12913_),
    .B(_10415_),
    .A_N(net6171));
 sg13g2_nand2_1 _26526_ (.Y(_12914_),
    .A(_00715_),
    .B(net6171));
 sg13g2_o21ai_1 _26527_ (.B1(_12914_),
    .Y(_12915_),
    .A1(net5915),
    .A2(_12913_));
 sg13g2_nand2_1 _26528_ (.Y(_12916_),
    .A(_00714_),
    .B(net6169));
 sg13g2_o21ai_1 _26529_ (.B1(_12916_),
    .Y(_12917_),
    .A1(net5783),
    .A2(net6069));
 sg13g2_nand2b_1 _26530_ (.Y(_12918_),
    .B(_10493_),
    .A_N(net6171));
 sg13g2_nand2_1 _26531_ (.Y(_12919_),
    .A(_00713_),
    .B(net6171));
 sg13g2_o21ai_1 _26532_ (.B1(_12919_),
    .Y(_12920_),
    .A1(net5908),
    .A2(_12918_));
 sg13g2_mux2_1 _26533_ (.A0(net5838),
    .A1(_00712_),
    .S(net6069),
    .X(_12921_));
 sg13g2_nand2_1 _26534_ (.Y(_12922_),
    .A(_00711_),
    .B(_12890_));
 sg13g2_o21ai_1 _26535_ (.B1(_12922_),
    .Y(_12923_),
    .A1(net5836),
    .A2(_12891_));
 sg13g2_nand2_1 _26536_ (.Y(_12924_),
    .A(_00710_),
    .B(net6169));
 sg13g2_nand4_1 _26537_ (.B(net7471),
    .C(_12902_),
    .A(net7548),
    .Y(_12925_),
    .D(_12907_));
 sg13g2_o21ai_1 _26538_ (.B1(_12924_),
    .Y(_12926_),
    .A1(net5902),
    .A2(net6069));
 sg13g2_nand2_1 _26539_ (.Y(_12927_),
    .A(_00709_),
    .B(net6169));
 sg13g2_o21ai_1 _26540_ (.B1(_12927_),
    .Y(_12928_),
    .A1(net5897),
    .A2(net6069));
 sg13g2_nand2_1 _26541_ (.Y(_12929_),
    .A(net7846),
    .B(_00891_));
 sg13g2_nand2_1 _26542_ (.Y(_12930_),
    .A(_00708_),
    .B(net6170));
 sg13g2_o21ai_1 _26543_ (.B1(_12930_),
    .Y(_12931_),
    .A1(net5888),
    .A2(net6170));
 sg13g2_mux2_1 _26544_ (.A0(net5772),
    .A1(_00707_),
    .S(net6171),
    .X(_12932_));
 sg13g2_nand2b_1 _26545_ (.Y(_12933_),
    .B(_00856_),
    .A_N(net7846));
 sg13g2_nand2_1 _26546_ (.Y(_12934_),
    .A(_00706_),
    .B(net6170));
 sg13g2_o21ai_1 _26547_ (.B1(_12934_),
    .Y(_12935_),
    .A1(net5885),
    .A2(net6170));
 sg13g2_nand2_1 _26548_ (.Y(_12936_),
    .A(_00705_),
    .B(net6174));
 sg13g2_o21ai_1 _26549_ (.B1(_12936_),
    .Y(_12937_),
    .A1(net5925),
    .A2(net6175));
 sg13g2_nand2_1 _26550_ (.Y(_12938_),
    .A(_00704_),
    .B(net6172));
 sg13g2_o21ai_1 _26551_ (.B1(_12938_),
    .Y(_12939_),
    .A1(net5962),
    .A2(net6172));
 sg13g2_nand2_1 _26552_ (.Y(_12940_),
    .A(_00703_),
    .B(net6172));
 sg13g2_o21ai_1 _26553_ (.B1(_12940_),
    .Y(_12941_),
    .A1(net6014),
    .A2(net6172));
 sg13g2_nand2_1 _26554_ (.Y(_12942_),
    .A(_00702_),
    .B(net6169));
 sg13g2_o21ai_1 _26555_ (.B1(_12942_),
    .Y(_12943_),
    .A1(net5957),
    .A2(net6069));
 sg13g2_nand2_1 _26556_ (.Y(_12944_),
    .A(_00701_),
    .B(net6173));
 sg13g2_o21ai_1 _26557_ (.B1(_12944_),
    .Y(_12945_),
    .A1(net6010),
    .A2(net6173));
 sg13g2_nand2_1 _26558_ (.Y(_12946_),
    .A(_00700_),
    .B(net6173));
 sg13g2_o21ai_1 _26559_ (.B1(_12946_),
    .Y(_12947_),
    .A1(net6006),
    .A2(net6173));
 sg13g2_nand2_1 _26560_ (.Y(_12948_),
    .A(_00699_),
    .B(net6174));
 sg13g2_o21ai_1 _26561_ (.B1(_12948_),
    .Y(_12949_),
    .A1(_09678_),
    .A2(net6174));
 sg13g2_nand2_1 _26562_ (.Y(_12950_),
    .A(_00698_),
    .B(net6172));
 sg13g2_o21ai_1 _26563_ (.B1(_12950_),
    .Y(_12951_),
    .A1(net6033),
    .A2(net6172));
 sg13g2_nand4_1 _26564_ (.B(net7462),
    .C(_12929_),
    .A(net7548),
    .Y(_12952_),
    .D(_12933_));
 sg13g2_nand2_1 _26565_ (.Y(_12953_),
    .A(_00697_),
    .B(net6175));
 sg13g2_o21ai_1 _26566_ (.B1(_12953_),
    .Y(_12954_),
    .A1(net6109),
    .A2(net6175));
 sg13g2_nand2_1 _26567_ (.Y(_12955_),
    .A(_00696_),
    .B(net6174));
 sg13g2_o21ai_1 _26568_ (.B1(_12955_),
    .Y(_12956_),
    .A1(_09902_),
    .A2(net6174));
 sg13g2_nand2_1 _26569_ (.Y(_12957_),
    .A(_00695_),
    .B(net6170));
 sg13g2_o21ai_1 _26570_ (.B1(_12957_),
    .Y(_12958_),
    .A1(net6055),
    .A2(net6170));
 sg13g2_nand2_1 _26571_ (.Y(_12959_),
    .A(_00694_),
    .B(net6173));
 sg13g2_o21ai_1 _26572_ (.B1(_12959_),
    .Y(_12960_),
    .A1(net6022),
    .A2(net6173));
 sg13g2_nand2_1 _26573_ (.Y(_12961_),
    .A(_00693_),
    .B(net6170));
 sg13g2_o21ai_1 _26574_ (.B1(_12961_),
    .Y(_12962_),
    .A1(net6108),
    .A2(net6170));
 sg13g2_nand2_1 _26575_ (.Y(_12963_),
    .A(_00692_),
    .B(net6169));
 sg13g2_nand2_1 _26576_ (.Y(_12964_),
    .A(net7846),
    .B(_01032_));
 sg13g2_o21ai_1 _26577_ (.B1(_12963_),
    .Y(_12965_),
    .A1(net5864),
    .A2(net6069));
 sg13g2_or4_1 _26578_ (.A(net7668),
    .B(_06622_),
    .C(net6468),
    .D(_11478_),
    .X(_12966_));
 sg13g2_nand3_1 _26579_ (.B(_10990_),
    .C(net7446),
    .A(_06621_),
    .Y(_12967_));
 sg13g2_nand2_1 _26580_ (.Y(_12968_),
    .A(_00691_),
    .B(net6167));
 sg13g2_nand2b_1 _26581_ (.Y(_12969_),
    .B(_00997_),
    .A_N(net7847));
 sg13g2_o21ai_1 _26582_ (.B1(_12968_),
    .Y(_12970_),
    .A1(net5861),
    .A2(net6167));
 sg13g2_nand2_1 _26583_ (.Y(_12971_),
    .A(_00690_),
    .B(net6168));
 sg13g2_nand2b_1 _26584_ (.Y(_12972_),
    .B(net6381),
    .A_N(net6168));
 sg13g2_o21ai_1 _26585_ (.B1(_12971_),
    .Y(_12973_),
    .A1(net5855),
    .A2(_12972_));
 sg13g2_nand2_1 _26586_ (.Y(_12974_),
    .A(_00689_),
    .B(net6164));
 sg13g2_o21ai_1 _26587_ (.B1(_12974_),
    .Y(_12975_),
    .A1(net5804),
    .A2(net6068));
 sg13g2_nand2_1 _26588_ (.Y(_12976_),
    .A(_00688_),
    .B(net6167));
 sg13g2_o21ai_1 _26589_ (.B1(_12976_),
    .Y(_12977_),
    .A1(net5847),
    .A2(net6167));
 sg13g2_nand2_1 _26590_ (.Y(_12978_),
    .A(_00687_),
    .B(net6166));
 sg13g2_o21ai_1 _26591_ (.B1(_12978_),
    .Y(_12979_),
    .A1(net5798),
    .A2(net6166));
 sg13g2_nand2_1 _26592_ (.Y(_12980_),
    .A(_00686_),
    .B(net6160));
 sg13g2_o21ai_1 _26593_ (.B1(_12980_),
    .Y(_12981_),
    .A1(net5792),
    .A2(net6068));
 sg13g2_nand2_1 _26594_ (.Y(_12982_),
    .A(_00685_),
    .B(net6166));
 sg13g2_nand2b_1 _26595_ (.Y(_12983_),
    .B(net6377),
    .A_N(_12966_));
 sg13g2_o21ai_1 _26596_ (.B1(_12982_),
    .Y(_12984_),
    .A1(net5920),
    .A2(_12983_));
 sg13g2_nand2_1 _26597_ (.Y(_12985_),
    .A(_00684_),
    .B(net6160));
 sg13g2_o21ai_1 _26598_ (.B1(_12985_),
    .Y(_12986_),
    .A1(net5785),
    .A2(net6068));
 sg13g2_nand4_1 _26599_ (.B(net7525),
    .C(_12964_),
    .A(net7548),
    .Y(_12987_),
    .D(_12969_));
 sg13g2_nand2_1 _26600_ (.Y(_12988_),
    .A(_00683_),
    .B(_12966_));
 sg13g2_nand2b_1 _26601_ (.Y(_12989_),
    .B(_10415_),
    .A_N(_12966_));
 sg13g2_o21ai_1 _26602_ (.B1(_12988_),
    .Y(_12990_),
    .A1(net5915),
    .A2(_12989_));
 sg13g2_nand2_1 _26603_ (.Y(_12991_),
    .A(_00682_),
    .B(net6164));
 sg13g2_nand2_1 _26604_ (.Y(_12992_),
    .A(net7846),
    .B(_00962_));
 sg13g2_o21ai_1 _26605_ (.B1(_12991_),
    .Y(_12993_),
    .A1(net5783),
    .A2(net6068));
 sg13g2_nand2_1 _26606_ (.Y(_12994_),
    .A(_00681_),
    .B(_12966_));
 sg13g2_nand2b_1 _26607_ (.Y(_12995_),
    .B(net6364),
    .A_N(_12966_));
 sg13g2_o21ai_1 _26608_ (.B1(_12994_),
    .Y(_12996_),
    .A1(net5908),
    .A2(_12995_));
 sg13g2_nand2b_1 _26609_ (.Y(_12997_),
    .B(_00926_),
    .A_N(net7846));
 sg13g2_mux2_1 _26610_ (.A0(net5838),
    .A1(_00680_),
    .S(_12967_),
    .X(_12998_));
 sg13g2_nand2_1 _26611_ (.Y(_12999_),
    .A(_00679_),
    .B(net6160));
 sg13g2_o21ai_1 _26612_ (.B1(_12999_),
    .Y(_13000_),
    .A1(net5836),
    .A2(net6068));
 sg13g2_nand2_1 _26613_ (.Y(_13001_),
    .A(_00678_),
    .B(net6164));
 sg13g2_o21ai_1 _26614_ (.B1(_13001_),
    .Y(_13002_),
    .A1(net5902),
    .A2(net6068));
 sg13g2_nand2_1 _26615_ (.Y(_13003_),
    .A(_00677_),
    .B(net6164));
 sg13g2_o21ai_1 _26616_ (.B1(_13003_),
    .Y(_13004_),
    .A1(net5897),
    .A2(net6068));
 sg13g2_nand2_1 _26617_ (.Y(_13005_),
    .A(_00676_),
    .B(net6165));
 sg13g2_o21ai_1 _26618_ (.B1(_13005_),
    .Y(_13006_),
    .A1(net5888),
    .A2(net6165));
 sg13g2_mux2_1 _26619_ (.A0(net5772),
    .A1(_00675_),
    .S(_12966_),
    .X(_13007_));
 sg13g2_nand2_1 _26620_ (.Y(_13008_),
    .A(_00674_),
    .B(net6161));
 sg13g2_o21ai_1 _26621_ (.B1(_13008_),
    .Y(_13009_),
    .A1(net5885),
    .A2(net6161));
 sg13g2_nand2_1 _26622_ (.Y(_13010_),
    .A(_00673_),
    .B(net6168));
 sg13g2_nand4_1 _26623_ (.B(net7512),
    .C(_12992_),
    .A(net7548),
    .Y(_13011_),
    .D(_12997_));
 sg13g2_o21ai_1 _26624_ (.B1(_13010_),
    .Y(_13012_),
    .A1(net5929),
    .A2(net6168));
 sg13g2_nand2_1 _26625_ (.Y(_13013_),
    .A(_00672_),
    .B(net6163));
 sg13g2_o21ai_1 _26626_ (.B1(_13013_),
    .Y(_13014_),
    .A1(net5962),
    .A2(net6163));
 sg13g2_nand2_1 _26627_ (.Y(_13015_),
    .A(_00671_),
    .B(net6163));
 sg13g2_o21ai_1 _26628_ (.B1(_13015_),
    .Y(_13016_),
    .A1(net6014),
    .A2(net6163));
 sg13g2_nand2_1 _26629_ (.Y(_13017_),
    .A(_00670_),
    .B(net6165));
 sg13g2_nand2_1 _26630_ (.Y(_13018_),
    .A(net7849),
    .B(_01384_));
 sg13g2_o21ai_1 _26631_ (.B1(_13017_),
    .Y(_13019_),
    .A1(net5957),
    .A2(_12967_));
 sg13g2_nand2_1 _26632_ (.Y(_13020_),
    .A(_00669_),
    .B(net6162));
 sg13g2_o21ai_1 _26633_ (.B1(_13020_),
    .Y(_13021_),
    .A1(net6010),
    .A2(net6162));
 sg13g2_nand2_1 _26634_ (.Y(_13022_),
    .A(_00668_),
    .B(net6162));
 sg13g2_nand2b_1 _26635_ (.Y(_13023_),
    .B(_01349_),
    .A_N(net7849));
 sg13g2_o21ai_1 _26636_ (.B1(_13022_),
    .Y(_13024_),
    .A1(net6006),
    .A2(net6162));
 sg13g2_nand2_1 _26637_ (.Y(_13025_),
    .A(_00667_),
    .B(net6167));
 sg13g2_o21ai_1 _26638_ (.B1(_13025_),
    .Y(_13026_),
    .A1(_09678_),
    .A2(net6167));
 sg13g2_nand2_1 _26639_ (.Y(_13027_),
    .A(_00666_),
    .B(net6163));
 sg13g2_o21ai_1 _26640_ (.B1(_13027_),
    .Y(_13028_),
    .A1(net6033),
    .A2(net6163));
 sg13g2_nand2_1 _26641_ (.Y(_13029_),
    .A(_00665_),
    .B(net6168));
 sg13g2_o21ai_1 _26642_ (.B1(_13029_),
    .Y(_13030_),
    .A1(net6109),
    .A2(net6168));
 sg13g2_nand2_1 _26643_ (.Y(_13031_),
    .A(_00664_),
    .B(net6167));
 sg13g2_o21ai_1 _26644_ (.B1(_13031_),
    .Y(_13032_),
    .A1(_09902_),
    .A2(net6167));
 sg13g2_nand2_1 _26645_ (.Y(_13033_),
    .A(_00663_),
    .B(net6161));
 sg13g2_o21ai_1 _26646_ (.B1(_13033_),
    .Y(_13034_),
    .A1(net6055),
    .A2(net6161));
 sg13g2_nand2_1 _26647_ (.Y(_13035_),
    .A(_00662_),
    .B(net6161));
 sg13g2_o21ai_1 _26648_ (.B1(_13035_),
    .Y(_13036_),
    .A1(net6022),
    .A2(net6161));
 sg13g2_nand2_1 _26649_ (.Y(_13037_),
    .A(_00661_),
    .B(net6161));
 sg13g2_o21ai_1 _26650_ (.B1(_13037_),
    .Y(_13038_),
    .A1(net6108),
    .A2(net6161));
 sg13g2_nand2_1 _26651_ (.Y(_13039_),
    .A(_00660_),
    .B(net6164));
 sg13g2_nand4_1 _26652_ (.B(net7471),
    .C(_13018_),
    .A(net7494),
    .Y(_13040_),
    .D(_13023_));
 sg13g2_o21ai_1 _26653_ (.B1(_13039_),
    .Y(_13041_),
    .A1(net5864),
    .A2(net6068));
 sg13g2_nand2_1 _26654_ (.Y(_13042_),
    .A(_00659_),
    .B(net6045));
 sg13g2_o21ai_1 _26655_ (.B1(_13042_),
    .Y(_13043_),
    .A1(net6045),
    .A2(net8286));
 sg13g2_nand2_1 _26656_ (.Y(_13044_),
    .A(_09610_),
    .B(net6382));
 sg13g2_nand2_1 _26657_ (.Y(_13045_),
    .A(_00658_),
    .B(net6045));
 sg13g2_o21ai_1 _26658_ (.B1(_13045_),
    .Y(_13046_),
    .A1(net5854),
    .A2(_13044_));
 sg13g2_nand2_1 _26659_ (.Y(_13047_),
    .A(net7849),
    .B(_01454_));
 sg13g2_nand2_1 _26660_ (.Y(_13048_),
    .A(_00657_),
    .B(net6043));
 sg13g2_o21ai_1 _26661_ (.B1(_13048_),
    .Y(_13049_),
    .A1(net6043),
    .A2(net5804));
 sg13g2_nand2_1 _26662_ (.Y(_13050_),
    .A(_00656_),
    .B(net6046));
 sg13g2_o21ai_1 _26663_ (.B1(_13050_),
    .Y(_13051_),
    .A1(net6046),
    .A2(net5847));
 sg13g2_nand2_1 _26664_ (.Y(_13052_),
    .A(_00655_),
    .B(net6045));
 sg13g2_nand2b_1 _26665_ (.Y(_13053_),
    .B(_01419_),
    .A_N(net7849));
 sg13g2_o21ai_1 _26666_ (.B1(_13052_),
    .Y(_13054_),
    .A1(net6045),
    .A2(net5803));
 sg13g2_nand2_1 _26667_ (.Y(_13055_),
    .A(_00654_),
    .B(net6044));
 sg13g2_o21ai_1 _26668_ (.B1(_13055_),
    .Y(_13056_),
    .A1(net6044),
    .A2(net5792));
 sg13g2_nand2_1 _26669_ (.Y(_13057_),
    .A(_09610_),
    .B(net6377));
 sg13g2_nand2_1 _26670_ (.Y(_13058_),
    .A(_00653_),
    .B(net6045));
 sg13g2_o21ai_1 _26671_ (.B1(_13058_),
    .Y(_13059_),
    .A1(net5917),
    .A2(_13057_));
 sg13g2_nand2_1 _26672_ (.Y(_13060_),
    .A(_00652_),
    .B(net6048));
 sg13g2_o21ai_1 _26673_ (.B1(_13060_),
    .Y(_13061_),
    .A1(net6048),
    .A2(net5786));
 sg13g2_nand2_1 _26674_ (.Y(_13062_),
    .A(_09610_),
    .B(net6370));
 sg13g2_nand2_1 _26675_ (.Y(_13063_),
    .A(_00651_),
    .B(net6044));
 sg13g2_o21ai_1 _26676_ (.B1(_13063_),
    .Y(_13064_),
    .A1(net5915),
    .A2(_13062_));
 sg13g2_nand2_1 _26677_ (.Y(_13065_),
    .A(_00650_),
    .B(net6043));
 sg13g2_o21ai_1 _26678_ (.B1(_13065_),
    .Y(_13066_),
    .A1(net6043),
    .A2(net5783));
 sg13g2_nand2_1 _26679_ (.Y(_13067_),
    .A(_09610_),
    .B(net6365));
 sg13g2_nand2_1 _26680_ (.Y(_13068_),
    .A(_00649_),
    .B(net6044));
 sg13g2_o21ai_1 _26681_ (.B1(_13068_),
    .Y(_13069_),
    .A1(net5911),
    .A2(_13067_));
 sg13g2_mux2_1 _26682_ (.A0(_00648_),
    .A1(net5838),
    .S(_09610_),
    .X(_13070_));
 sg13g2_nand2_1 _26683_ (.Y(_13071_),
    .A(_00647_),
    .B(net6048));
 sg13g2_o21ai_1 _26684_ (.B1(_13071_),
    .Y(_13072_),
    .A1(net6048),
    .A2(net5836));
 sg13g2_nand2_1 _26685_ (.Y(_13073_),
    .A(_00646_),
    .B(_09611_));
 sg13g2_o21ai_1 _26686_ (.B1(_13073_),
    .Y(_13074_),
    .A1(_09611_),
    .A2(net5902));
 sg13g2_nand2_1 _26687_ (.Y(_13075_),
    .A(_00645_),
    .B(_09611_));
 sg13g2_nand4_1 _26688_ (.B(net7462),
    .C(_13047_),
    .A(net7494),
    .Y(_13076_),
    .D(_13053_));
 sg13g2_o21ai_1 _26689_ (.B1(_13075_),
    .Y(_13077_),
    .A1(_09611_),
    .A2(net5897));
 sg13g2_nand2_1 _26690_ (.Y(_13078_),
    .A(_00644_),
    .B(net6044));
 sg13g2_o21ai_1 _26691_ (.B1(_13078_),
    .Y(_13079_),
    .A1(net6044),
    .A2(net5894));
 sg13g2_mux2_1 _26692_ (.A0(_00643_),
    .A1(net5772),
    .S(_09610_),
    .X(_13080_));
 sg13g2_nand2_1 _26693_ (.Y(_13081_),
    .A(_00642_),
    .B(net6048));
 sg13g2_o21ai_1 _26694_ (.B1(_13081_),
    .Y(_13082_),
    .A1(net6048),
    .A2(net5885));
 sg13g2_nand2_1 _26695_ (.Y(_13083_),
    .A(_00641_),
    .B(net6046));
 sg13g2_o21ai_1 _26696_ (.B1(_13083_),
    .Y(_13084_),
    .A1(net6046),
    .A2(net5925));
 sg13g2_nand2_1 _26697_ (.Y(_13085_),
    .A(_00640_),
    .B(net6049));
 sg13g2_o21ai_1 _26698_ (.B1(_13085_),
    .Y(_13086_),
    .A1(net6049),
    .A2(net5962));
 sg13g2_nand2_1 _26699_ (.Y(_13087_),
    .A(_00639_),
    .B(net6049));
 sg13g2_o21ai_1 _26700_ (.B1(_13087_),
    .Y(_13088_),
    .A1(net6049),
    .A2(net6014));
 sg13g2_nand2_1 _26701_ (.Y(_13089_),
    .A(_00638_),
    .B(net6043));
 sg13g2_o21ai_1 _26702_ (.B1(_13089_),
    .Y(_13090_),
    .A1(net6043),
    .A2(net5957));
 sg13g2_nand2_1 _26703_ (.Y(_13091_),
    .A(_00637_),
    .B(net6049));
 sg13g2_o21ai_1 _26704_ (.B1(_13091_),
    .Y(_13092_),
    .A1(net6049),
    .A2(net6010));
 sg13g2_nand2_1 _26705_ (.Y(_13093_),
    .A(_00636_),
    .B(net6050));
 sg13g2_o21ai_1 _26706_ (.B1(_13093_),
    .Y(_13094_),
    .A1(net6050),
    .A2(net6006));
 sg13g2_nand2_1 _26707_ (.Y(_13095_),
    .A(_00635_),
    .B(net6046));
 sg13g2_o21ai_1 _26708_ (.B1(_13095_),
    .Y(_13096_),
    .A1(net6046),
    .A2(net6117));
 sg13g2_nand2_1 _26709_ (.Y(_13097_),
    .A(_00634_),
    .B(net6049));
 sg13g2_o21ai_1 _26710_ (.B1(_13097_),
    .Y(_13098_),
    .A1(net6049),
    .A2(net6033));
 sg13g2_nand2_1 _26711_ (.Y(_13099_),
    .A(_00633_),
    .B(net6036));
 sg13g2_o21ai_1 _26712_ (.B1(_13099_),
    .Y(_13100_),
    .A1(net6036),
    .A2(net5860));
 sg13g2_nand2_1 _26713_ (.Y(_13101_),
    .A(net6116),
    .B(_10162_));
 sg13g2_nand2_1 _26714_ (.Y(_13102_),
    .A(_00632_),
    .B(net6036));
 sg13g2_o21ai_1 _26715_ (.B1(_13102_),
    .Y(_13103_),
    .A1(net5854),
    .A2(_13101_));
 sg13g2_nand2_1 _26716_ (.Y(_13104_),
    .A(_00631_),
    .B(net6038));
 sg13g2_o21ai_1 _26717_ (.B1(_13104_),
    .Y(_13105_),
    .A1(net6038),
    .A2(net5808));
 sg13g2_nand2_1 _26718_ (.Y(_13106_),
    .A(_00630_),
    .B(net6034));
 sg13g2_o21ai_1 _26719_ (.B1(_13106_),
    .Y(_13107_),
    .A1(net6035),
    .A2(net5849));
 sg13g2_nand2_1 _26720_ (.Y(_13108_),
    .A(_00629_),
    .B(net6045));
 sg13g2_o21ai_1 _26721_ (.B1(_13108_),
    .Y(_13109_),
    .A1(net6045),
    .A2(net6110));
 sg13g2_nand2_1 _26722_ (.Y(_13110_),
    .A(_00628_),
    .B(net6035));
 sg13g2_o21ai_1 _26723_ (.B1(_13110_),
    .Y(_13111_),
    .A1(net6035),
    .A2(net5800));
 sg13g2_nand4_1 _26724_ (.B(_12987_),
    .C(_13040_),
    .A(_12925_),
    .Y(_13112_),
    .D(_13076_));
 sg13g2_nand2_1 _26725_ (.Y(_13113_),
    .A(_00627_),
    .B(net6037));
 sg13g2_o21ai_1 _26726_ (.B1(_13113_),
    .Y(_13114_),
    .A1(net6037),
    .A2(net5795));
 sg13g2_nand2_1 _26727_ (.Y(_13115_),
    .A(net6116),
    .B(_10341_));
 sg13g2_nand2_1 _26728_ (.Y(_13116_),
    .A(_00626_),
    .B(net6036));
 sg13g2_o21ai_1 _26729_ (.B1(_13116_),
    .Y(_13117_),
    .A1(net5921),
    .A2(_13115_));
 sg13g2_nand2_1 _26730_ (.Y(_13118_),
    .A(_00625_),
    .B(net6037));
 sg13g2_o21ai_1 _26731_ (.B1(_13118_),
    .Y(_13119_),
    .A1(net6037),
    .A2(net5789));
 sg13g2_nand2_1 _26732_ (.Y(_13120_),
    .A(net6116),
    .B(net6373));
 sg13g2_nand2_1 _26733_ (.Y(_13121_),
    .A(_00624_),
    .B(net6036));
 sg13g2_o21ai_1 _26734_ (.B1(_13121_),
    .Y(_13122_),
    .A1(net5914),
    .A2(_13120_));
 sg13g2_nand2_1 _26735_ (.Y(_13123_),
    .A(_00623_),
    .B(net6039));
 sg13g2_o21ai_1 _26736_ (.B1(_13123_),
    .Y(_13124_),
    .A1(net6039),
    .A2(net5778));
 sg13g2_nand2_1 _26737_ (.Y(_13125_),
    .A(net6116),
    .B(net6366));
 sg13g2_nand2_1 _26738_ (.Y(_13126_),
    .A(_00622_),
    .B(net6036));
 sg13g2_o21ai_1 _26739_ (.B1(_13126_),
    .Y(_13127_),
    .A1(net5910),
    .A2(_13125_));
 sg13g2_nand4_1 _26740_ (.B(_12895_),
    .C(_12952_),
    .A(_12868_),
    .Y(_13128_),
    .D(_13011_));
 sg13g2_mux2_1 _26741_ (.A0(_00621_),
    .A1(net5843),
    .S(net6116),
    .X(_13129_));
 sg13g2_nand2_1 _26742_ (.Y(_13130_),
    .A(_00620_),
    .B(net6042));
 sg13g2_o21ai_1 _26743_ (.B1(_13130_),
    .Y(_13131_),
    .A1(net6042),
    .A2(net5833));
 sg13g2_nand2_1 _26744_ (.Y(_13132_),
    .A(_00619_),
    .B(net6039));
 sg13g2_o21ai_1 _26745_ (.B1(_13132_),
    .Y(_13133_),
    .A1(net6038),
    .A2(net5900));
 sg13g2_nand2_1 _26746_ (.Y(_13134_),
    .A(_00618_),
    .B(net6046));
 sg13g2_o21ai_1 _26747_ (.B1(_13134_),
    .Y(_13135_),
    .A1(net6046),
    .A2(_09902_));
 sg13g2_nand2_1 _26748_ (.Y(_13136_),
    .A(_00617_),
    .B(net6038));
 sg13g2_o21ai_1 _26749_ (.B1(_13136_),
    .Y(_13137_),
    .A1(net6038),
    .A2(net5895));
 sg13g2_nand2_1 _26750_ (.Y(_13138_),
    .A(_00616_),
    .B(net6040));
 sg13g2_o21ai_1 _26751_ (.B1(_13138_),
    .Y(_13139_),
    .A1(net6040),
    .A2(net5891));
 sg13g2_mux2_1 _26752_ (.A0(_00615_),
    .A1(net5775),
    .S(net6116),
    .X(_13140_));
 sg13g2_nand2_1 _26753_ (.Y(_13141_),
    .A(_00614_),
    .B(net6040));
 sg13g2_o21ai_1 _26754_ (.B1(_13141_),
    .Y(_13142_),
    .A1(net6040),
    .A2(net5882));
 sg13g2_nand2_1 _26755_ (.Y(_13143_),
    .A(_00613_),
    .B(net6035));
 sg13g2_o21ai_1 _26756_ (.B1(_13143_),
    .Y(_13144_),
    .A1(net6035),
    .A2(net5928));
 sg13g2_nand2_1 _26757_ (.Y(_13145_),
    .A(_00612_),
    .B(net6035));
 sg13g2_o21ai_1 _26758_ (.B1(_13145_),
    .Y(_13146_),
    .A1(net6035),
    .A2(net5966));
 sg13g2_nand2_1 _26759_ (.Y(_13147_),
    .A(_00611_),
    .B(net6041));
 sg13g2_mux2_1 _26760_ (.A0(_01258_),
    .A1(_00618_),
    .S(net7852),
    .X(_13148_));
 sg13g2_o21ai_1 _26761_ (.B1(_13147_),
    .Y(_13149_),
    .A1(net6041),
    .A2(net6012));
 sg13g2_nand2_1 _26762_ (.Y(_13150_),
    .A(_00610_),
    .B(net6037));
 sg13g2_o21ai_1 _26763_ (.B1(_13150_),
    .Y(_13151_),
    .A1(net6037),
    .A2(net5958));
 sg13g2_nand2_1 _26764_ (.Y(_13152_),
    .A(_00609_),
    .B(net6041));
 sg13g2_o21ai_1 _26765_ (.B1(_13152_),
    .Y(_13153_),
    .A1(net6041),
    .A2(net6009));
 sg13g2_nand2_1 _26766_ (.Y(_13154_),
    .A(_00608_),
    .B(net6040));
 sg13g2_o21ai_1 _26767_ (.B1(_13154_),
    .Y(_13155_),
    .A1(net6040),
    .A2(net6002));
 sg13g2_or2_1 _26768_ (.X(_13156_),
    .B(fetch_enable_q),
    .A(net350));
 sg13g2_nor2_1 _26769_ (.A(_05162_),
    .B(_08659_),
    .Y(_13157_));
 sg13g2_nand2_1 _26770_ (.Y(_13158_),
    .A(_00543_),
    .B(_08663_));
 sg13g2_nor2_1 _26771_ (.A(_08791_),
    .B(_13158_),
    .Y(_13159_));
 sg13g2_a21oi_1 _26772_ (.A1(_08986_),
    .A2(_13159_),
    .Y(_13160_),
    .B1(_00607_));
 sg13g2_nand2_1 _26773_ (.Y(_13161_),
    .A(net8003),
    .B(_08658_));
 sg13g2_nor2_1 _26774_ (.A(_13157_),
    .B(_13161_),
    .Y(_13162_));
 sg13g2_nand3_1 _26775_ (.B(net8003),
    .C(_08658_),
    .A(_05162_),
    .Y(_13163_));
 sg13g2_and2_1 _26776_ (.A(net7852),
    .B(_00906_),
    .X(_13164_));
 sg13g2_nor2_1 _26777_ (.A(_13160_),
    .B(net6750),
    .Y(_13165_));
 sg13g2_a21oi_1 _26778_ (.A1(_08999_),
    .A2(_13159_),
    .Y(_13166_),
    .B1(_00606_));
 sg13g2_nor2_1 _26779_ (.A(net6751),
    .B(_13166_),
    .Y(_13167_));
 sg13g2_and3_1 _26780_ (.X(_13168_),
    .A(_00543_),
    .B(_08663_),
    .C(_08850_));
 sg13g2_a21oi_1 _26781_ (.A1(_08957_),
    .A2(_13168_),
    .Y(_13169_),
    .B1(_00605_));
 sg13g2_nor2_1 _26782_ (.A(net6750),
    .B(_13169_),
    .Y(_13170_));
 sg13g2_a21oi_1 _26783_ (.A1(_08972_),
    .A2(_13168_),
    .Y(_13171_),
    .B1(_00604_));
 sg13g2_nor2_1 _26784_ (.A(net6750),
    .B(_13171_),
    .Y(_13172_));
 sg13g2_a21oi_1 _26785_ (.A1(_08986_),
    .A2(_13168_),
    .Y(_13173_),
    .B1(_00603_));
 sg13g2_nor2_1 _26786_ (.A(net6750),
    .B(_13173_),
    .Y(_13174_));
 sg13g2_a22oi_1 _26787_ (.Y(_13175_),
    .B1(_13168_),
    .B2(_08999_),
    .A2(_13163_),
    .A1(_00602_));
 sg13g2_inv_1 _26788_ (.Y(_13176_),
    .A(_13175_));
 sg13g2_nor2_1 _26789_ (.A(_08902_),
    .B(_13158_),
    .Y(_13177_));
 sg13g2_a21oi_1 _26790_ (.A1(_08957_),
    .A2(_13177_),
    .Y(_13178_),
    .B1(_00601_));
 sg13g2_nor2_1 _26791_ (.A(net6751),
    .B(_13178_),
    .Y(_13179_));
 sg13g2_and3_1 _26792_ (.X(_13180_),
    .A(_00543_),
    .B(_08663_),
    .C(net7431));
 sg13g2_a21oi_1 _26793_ (.A1(_08731_),
    .A2(_13180_),
    .Y(_13181_),
    .B1(_00600_));
 sg13g2_nor2_1 _26794_ (.A(net6752),
    .B(_13181_),
    .Y(_13182_));
 sg13g2_a21oi_1 _26795_ (.A1(_08744_),
    .A2(_13180_),
    .Y(_13183_),
    .B1(_00599_));
 sg13g2_nor2_1 _26796_ (.A(net6752),
    .B(_13183_),
    .Y(_13184_));
 sg13g2_a21oi_1 _26797_ (.A1(_08972_),
    .A2(_13177_),
    .Y(_13185_),
    .B1(_00598_));
 sg13g2_nor2_1 _26798_ (.A(net6751),
    .B(_13185_),
    .Y(_13186_));
 sg13g2_mux2_1 _26799_ (.A0(_00664_),
    .A1(_00696_),
    .S(net7852),
    .X(_13187_));
 sg13g2_a21oi_1 _26800_ (.A1(_08760_),
    .A2(_13180_),
    .Y(_13188_),
    .B1(_00597_));
 sg13g2_nor2_1 _26801_ (.A(net6749),
    .B(_13188_),
    .Y(_13189_));
 sg13g2_a22oi_1 _26802_ (.Y(_13190_),
    .B1(_13180_),
    .B2(_08774_),
    .A2(_13163_),
    .A1(_00596_));
 sg13g2_inv_1 _26803_ (.Y(_13191_),
    .A(_13190_));
 sg13g2_a21oi_1 _26804_ (.A1(_08731_),
    .A2(_13159_),
    .Y(_13192_),
    .B1(_00595_));
 sg13g2_nor2_1 _26805_ (.A(net6752),
    .B(_13192_),
    .Y(_13193_));
 sg13g2_a21oi_1 _26806_ (.A1(_08744_),
    .A2(_13159_),
    .Y(_13194_),
    .B1(_00594_));
 sg13g2_nor2_1 _26807_ (.A(net6752),
    .B(_13194_),
    .Y(_13195_));
 sg13g2_a21oi_1 _26808_ (.A1(_08760_),
    .A2(_13159_),
    .Y(_13196_),
    .B1(_00593_));
 sg13g2_nor2_1 _26809_ (.A(net6749),
    .B(_13196_),
    .Y(_13197_));
 sg13g2_a21oi_1 _26810_ (.A1(_08774_),
    .A2(_13159_),
    .Y(_13198_),
    .B1(_00592_));
 sg13g2_nor2_1 _26811_ (.A(net6752),
    .B(_13198_),
    .Y(_13199_));
 sg13g2_a21oi_1 _26812_ (.A1(_08731_),
    .A2(_13168_),
    .Y(_13200_),
    .B1(_00591_));
 sg13g2_nor2_1 _26813_ (.A(net6749),
    .B(_13200_),
    .Y(_13201_));
 sg13g2_mux2_1 _26814_ (.A0(_00728_),
    .A1(_00760_),
    .S(net7852),
    .X(_13202_));
 sg13g2_a21oi_1 _26815_ (.A1(_08744_),
    .A2(_13168_),
    .Y(_13203_),
    .B1(_00590_));
 sg13g2_nor2_1 _26816_ (.A(net6749),
    .B(_13203_),
    .Y(_13204_));
 sg13g2_a21oi_1 _26817_ (.A1(_08760_),
    .A2(_13168_),
    .Y(_13205_),
    .B1(_00589_));
 sg13g2_nor2_1 _26818_ (.A(net6749),
    .B(_13205_),
    .Y(_13206_));
 sg13g2_a22oi_1 _26819_ (.Y(_13207_),
    .B1(_13168_),
    .B2(_08774_),
    .A2(_13163_),
    .A1(_00588_));
 sg13g2_inv_1 _26820_ (.Y(_13208_),
    .A(_13207_));
 sg13g2_nand2_1 _26821_ (.Y(_13209_),
    .A(_00587_),
    .B(net6789));
 sg13g2_o21ai_1 _26822_ (.B1(_13209_),
    .Y(_13210_),
    .A1(_09130_),
    .A2(_13158_));
 sg13g2_a21oi_1 _26823_ (.A1(_08731_),
    .A2(_13177_),
    .Y(_13211_),
    .B1(_00586_));
 sg13g2_nor2_1 _26824_ (.A(net6749),
    .B(_13211_),
    .Y(_13212_));
 sg13g2_a21oi_1 _26825_ (.A1(_08744_),
    .A2(_13177_),
    .Y(_13213_),
    .B1(_00585_));
 sg13g2_nor2_1 _26826_ (.A(net6749),
    .B(_13213_),
    .Y(_13214_));
 sg13g2_a21oi_1 _26827_ (.A1(_08760_),
    .A2(_13177_),
    .Y(_13215_),
    .B1(_00584_));
 sg13g2_nor2_1 _26828_ (.A(net6749),
    .B(_13215_),
    .Y(_13216_));
 sg13g2_a21oi_1 _26829_ (.A1(_08939_),
    .A2(_13157_),
    .Y(_13217_),
    .B1(_00583_));
 sg13g2_nor2_1 _26830_ (.A(_13162_),
    .B(_13217_),
    .Y(_13218_));
 sg13g2_a21oi_1 _26831_ (.A1(_08957_),
    .A2(_13180_),
    .Y(_13219_),
    .B1(_00582_));
 sg13g2_nor2_1 _26832_ (.A(net6750),
    .B(_13219_),
    .Y(_13220_));
 sg13g2_a21oi_1 _26833_ (.A1(_08972_),
    .A2(_13180_),
    .Y(_13221_),
    .B1(_00581_));
 sg13g2_nor2_1 _26834_ (.A(net6750),
    .B(_13221_),
    .Y(_13222_));
 sg13g2_a21oi_1 _26835_ (.A1(_08986_),
    .A2(_13180_),
    .Y(_13223_),
    .B1(_00580_));
 sg13g2_nor2_1 _26836_ (.A(net6750),
    .B(_13223_),
    .Y(_13224_));
 sg13g2_a21oi_1 _26837_ (.A1(_08999_),
    .A2(_13180_),
    .Y(_13225_),
    .B1(_00579_));
 sg13g2_nor2_1 _26838_ (.A(net6751),
    .B(_13225_),
    .Y(_13226_));
 sg13g2_a21oi_1 _26839_ (.A1(_08957_),
    .A2(_13159_),
    .Y(_13227_),
    .B1(_00578_));
 sg13g2_nor2_1 _26840_ (.A(net6750),
    .B(_13227_),
    .Y(_13228_));
 sg13g2_a21oi_1 _26841_ (.A1(_08972_),
    .A2(_13159_),
    .Y(_13229_),
    .B1(_00577_));
 sg13g2_nor2_1 _26842_ (.A(net6752),
    .B(_13229_),
    .Y(_13230_));
 sg13g2_a21oi_1 _26843_ (.A1(_09144_),
    .A2(_13157_),
    .Y(_13231_),
    .B1(_00576_));
 sg13g2_nor2_1 _26844_ (.A(_13162_),
    .B(_13231_),
    .Y(_13232_));
 sg13g2_nand2_1 _26845_ (.Y(_13233_),
    .A(_00575_),
    .B(net6784));
 sg13g2_nand2_1 _26846_ (.Y(_13234_),
    .A(net7349),
    .B(_04796_));
 sg13g2_o21ai_1 _26847_ (.B1(_13234_),
    .Y(_13235_),
    .A1(net6625),
    .A2(_08688_));
 sg13g2_o21ai_1 _26848_ (.B1(_13233_),
    .Y(_13236_),
    .A1(net6784),
    .A2(_13235_));
 sg13g2_nand2_1 _26849_ (.Y(_13237_),
    .A(_00574_),
    .B(net6786));
 sg13g2_nor2_1 _26850_ (.A(_02067_),
    .B(net7043),
    .Y(_13238_));
 sg13g2_a21oi_1 _26851_ (.A1(net6626),
    .A2(net7040),
    .Y(_13239_),
    .B1(_13238_));
 sg13g2_o21ai_1 _26852_ (.B1(_13237_),
    .Y(_13240_),
    .A1(net6787),
    .A2(_13239_));
 sg13g2_nand2_1 _26853_ (.Y(_13241_),
    .A(_00573_),
    .B(net6786));
 sg13g2_nor2_1 _26854_ (.A(_15563_),
    .B(net7042),
    .Y(_13242_));
 sg13g2_a21oi_1 _26855_ (.A1(net6627),
    .A2(net7042),
    .Y(_13243_),
    .B1(_13242_));
 sg13g2_o21ai_1 _26856_ (.B1(_13241_),
    .Y(_13244_),
    .A1(net6787),
    .A2(_13243_));
 sg13g2_nand2_1 _26857_ (.Y(_13245_),
    .A(_00572_),
    .B(net6793));
 sg13g2_nand2_1 _26858_ (.Y(_13246_),
    .A(net7273),
    .B(net7318));
 sg13g2_o21ai_1 _26859_ (.B1(_13246_),
    .Y(_13247_),
    .A1(net6628),
    .A2(net7102));
 sg13g2_o21ai_1 _26860_ (.B1(_13245_),
    .Y(_13248_),
    .A1(net6790),
    .A2(_13247_));
 sg13g2_nand2_1 _26861_ (.Y(_13249_),
    .A(_00571_),
    .B(net6786));
 sg13g2_nand2_1 _26862_ (.Y(_13250_),
    .A(net7275),
    .B(net7318));
 sg13g2_o21ai_1 _26863_ (.B1(_13250_),
    .Y(_13251_),
    .A1(net6636),
    .A2(net7102));
 sg13g2_mux4_1 _26864_ (.S0(net7811),
    .A0(_13164_),
    .A1(_13187_),
    .A2(_13148_),
    .A3(_13202_),
    .S1(net7826),
    .X(_13252_));
 sg13g2_o21ai_1 _26865_ (.B1(_13249_),
    .Y(_13253_),
    .A1(net6788),
    .A2(_13251_));
 sg13g2_nor2_1 _26866_ (.A(net7529),
    .B(_13252_),
    .Y(_13254_));
 sg13g2_nand2_1 _26867_ (.Y(_13255_),
    .A(_00570_),
    .B(net6793));
 sg13g2_nor2_1 _26868_ (.A(_13358_),
    .B(net7044),
    .Y(_13256_));
 sg13g2_a21oi_1 _26869_ (.A1(net6638),
    .A2(net7044),
    .Y(_13257_),
    .B1(_13256_));
 sg13g2_o21ai_1 _26870_ (.B1(_13255_),
    .Y(_13258_),
    .A1(net6793),
    .A2(_13257_));
 sg13g2_nand2_1 _26871_ (.Y(_13259_),
    .A(_00569_),
    .B(net6786));
 sg13g2_nor2_1 _26872_ (.A(net7282),
    .B(net7042),
    .Y(_13260_));
 sg13g2_a21oi_1 _26873_ (.A1(net6639),
    .A2(net7043),
    .Y(_13261_),
    .B1(_13260_));
 sg13g2_o21ai_1 _26874_ (.B1(_13259_),
    .Y(_13262_),
    .A1(net6786),
    .A2(_13261_));
 sg13g2_nand2_1 _26875_ (.Y(_13263_),
    .A(_00568_),
    .B(net6790));
 sg13g2_o21ai_1 _26876_ (.B1(_03629_),
    .Y(_13264_),
    .A1(net6568),
    .A2(_04792_));
 sg13g2_o21ai_1 _26877_ (.B1(_13263_),
    .Y(_13265_),
    .A1(net6790),
    .A2(_13264_));
 sg13g2_nand2_1 _26878_ (.Y(_13266_),
    .A(_00567_),
    .B(net6789));
 sg13g2_nand2_1 _26879_ (.Y(_13267_),
    .A(net7328),
    .B(net7318));
 sg13g2_o21ai_1 _26880_ (.B1(_13267_),
    .Y(_13268_),
    .A1(net6569),
    .A2(net7102));
 sg13g2_o21ai_1 _26881_ (.B1(_13266_),
    .Y(_13269_),
    .A1(net6789),
    .A2(_13268_));
 sg13g2_nand2_1 _26882_ (.Y(_13270_),
    .A(_00566_),
    .B(net6792));
 sg13g2_nand2_1 _26883_ (.Y(_13271_),
    .A(net7283),
    .B(net7318));
 sg13g2_o21ai_1 _26884_ (.B1(_13271_),
    .Y(_13272_),
    .A1(net6640),
    .A2(net7102));
 sg13g2_o21ai_1 _26885_ (.B1(_13270_),
    .Y(_13273_),
    .A1(net6792),
    .A2(_13272_));
 sg13g2_nand2_1 _26886_ (.Y(_13274_),
    .A(_00565_),
    .B(net6784));
 sg13g2_nor2_1 _26887_ (.A(net7329),
    .B(_08687_),
    .Y(_13275_));
 sg13g2_a21oi_1 _26888_ (.A1(net6571),
    .A2(net7040),
    .Y(_13276_),
    .B1(_13275_));
 sg13g2_o21ai_1 _26889_ (.B1(_13274_),
    .Y(_13277_),
    .A1(net6784),
    .A2(_13276_));
 sg13g2_nand2_1 _26890_ (.Y(_13278_),
    .A(_00564_),
    .B(net6793));
 sg13g2_nor2_1 _26891_ (.A(net7331),
    .B(net7045),
    .Y(_13279_));
 sg13g2_a21oi_1 _26892_ (.A1(net6572),
    .A2(net7045),
    .Y(_13280_),
    .B1(_13279_));
 sg13g2_o21ai_1 _26893_ (.B1(_13278_),
    .Y(_13281_),
    .A1(net6789),
    .A2(_13280_));
 sg13g2_nand2_1 _26894_ (.Y(_13282_),
    .A(_00563_),
    .B(net6785));
 sg13g2_nor2_1 _26895_ (.A(_03367_),
    .B(net7043),
    .Y(_13283_));
 sg13g2_a21oi_1 _26896_ (.A1(net6575),
    .A2(net7041),
    .Y(_13284_),
    .B1(_13283_));
 sg13g2_o21ai_1 _26897_ (.B1(_13282_),
    .Y(_13285_),
    .A1(net6785),
    .A2(_13284_));
 sg13g2_nand2_1 _26898_ (.Y(_13286_),
    .A(_00562_),
    .B(net6785));
 sg13g2_nand2_1 _26899_ (.Y(_13287_),
    .A(net7332),
    .B(net7318));
 sg13g2_o21ai_1 _26900_ (.B1(_13287_),
    .Y(_13288_),
    .A1(net6576),
    .A2(net7102));
 sg13g2_o21ai_1 _26901_ (.B1(_13286_),
    .Y(_13289_),
    .A1(net6785),
    .A2(_13288_));
 sg13g2_mux4_1 _26902_ (.S0(net7892),
    .A0(_01067_),
    .A1(_01102_),
    .A2(_01138_),
    .A3(_01173_),
    .S1(net7825),
    .X(_13290_));
 sg13g2_nand2_1 _26903_ (.Y(_13291_),
    .A(_00561_),
    .B(net6785));
 sg13g2_nor2_1 _26904_ (.A(net7333),
    .B(net7043),
    .Y(_13292_));
 sg13g2_a21oi_1 _26905_ (.A1(net6579),
    .A2(net7041),
    .Y(_13293_),
    .B1(_13292_));
 sg13g2_o21ai_1 _26906_ (.B1(_13291_),
    .Y(_13294_),
    .A1(net6785),
    .A2(_13293_));
 sg13g2_nand2_1 _26907_ (.Y(_13295_),
    .A(_00560_),
    .B(net6785));
 sg13g2_nand2_1 _26908_ (.Y(_13296_),
    .A(net7334),
    .B(net7318));
 sg13g2_o21ai_1 _26909_ (.B1(_13296_),
    .Y(_13297_),
    .A1(net6582),
    .A2(net7102));
 sg13g2_o21ai_1 _26910_ (.B1(_13295_),
    .Y(_13298_),
    .A1(net6785),
    .A2(_13297_));
 sg13g2_nand2_1 _26911_ (.Y(_13299_),
    .A(_00559_),
    .B(net6786));
 sg13g2_nor2_1 _26912_ (.A(net7336),
    .B(net7040),
    .Y(_13300_));
 sg13g2_a21oi_1 _26913_ (.A1(net6603),
    .A2(net7040),
    .Y(_13301_),
    .B1(_13300_));
 sg13g2_o21ai_1 _26914_ (.B1(_13299_),
    .Y(_13302_),
    .A1(net6786),
    .A2(_13301_));
 sg13g2_nand2_1 _26915_ (.Y(_13303_),
    .A(_00558_),
    .B(net6787));
 sg13g2_nor2_1 _26916_ (.A(net7338),
    .B(net7041),
    .Y(_13304_));
 sg13g2_a21oi_1 _26917_ (.A1(net6605),
    .A2(net7041),
    .Y(_13305_),
    .B1(_13304_));
 sg13g2_o21ai_1 _26918_ (.B1(_13303_),
    .Y(_13306_),
    .A1(net6788),
    .A2(_13305_));
 sg13g2_nand2_1 _26919_ (.Y(_13307_),
    .A(_00557_),
    .B(net6787));
 sg13g2_nor2_1 _26920_ (.A(net7340),
    .B(net7041),
    .Y(_13308_));
 sg13g2_a21oi_1 _26921_ (.A1(net6584),
    .A2(net7041),
    .Y(_13309_),
    .B1(_13308_));
 sg13g2_o21ai_1 _26922_ (.B1(_13307_),
    .Y(_13310_),
    .A1(net6788),
    .A2(_13309_));
 sg13g2_nand2_1 _26923_ (.Y(_13311_),
    .A(_00556_),
    .B(net6787));
 sg13g2_nor2_1 _26924_ (.A(net7341),
    .B(net7041),
    .Y(_13312_));
 sg13g2_a21oi_1 _26925_ (.A1(net6586),
    .A2(net7041),
    .Y(_13313_),
    .B1(_13312_));
 sg13g2_o21ai_1 _26926_ (.B1(_13311_),
    .Y(_13314_),
    .A1(net6788),
    .A2(_13313_));
 sg13g2_nand2_1 _26927_ (.Y(_13315_),
    .A(_00555_),
    .B(net6790));
 sg13g2_nor2_1 _26928_ (.A(net7076),
    .B(net7044),
    .Y(_13316_));
 sg13g2_a21oi_1 _26929_ (.A1(net6717),
    .A2(net7044),
    .Y(_13317_),
    .B1(_13316_));
 sg13g2_o21ai_1 _26930_ (.B1(_13315_),
    .Y(_13318_),
    .A1(net6790),
    .A2(_13317_));
 sg13g2_nand2_1 _26931_ (.Y(_13319_),
    .A(_00554_),
    .B(net6788));
 sg13g2_nor2_1 _26932_ (.A(_02818_),
    .B(net7040),
    .Y(_13320_));
 sg13g2_a21oi_1 _26933_ (.A1(net6607),
    .A2(net7040),
    .Y(_13321_),
    .B1(_13320_));
 sg13g2_o21ai_1 _26934_ (.B1(_13319_),
    .Y(_13322_),
    .A1(net6783),
    .A2(_13321_));
 sg13g2_nand2_1 _26935_ (.Y(_13323_),
    .A(_00553_),
    .B(net6788));
 sg13g2_nor2_1 _26936_ (.A(net7343),
    .B(net7040),
    .Y(_13324_));
 sg13g2_a21oi_1 _26937_ (.A1(net6608),
    .A2(net7043),
    .Y(_13325_),
    .B1(_13324_));
 sg13g2_mux4_1 _26938_ (.S0(net7892),
    .A0(_01208_),
    .A1(_01243_),
    .A2(_01278_),
    .A3(_01314_),
    .S1(net7825),
    .X(_13326_));
 sg13g2_o21ai_1 _26939_ (.B1(_13323_),
    .Y(_13327_),
    .A1(net6783),
    .A2(_13325_));
 sg13g2_nand2_1 _26940_ (.Y(_13328_),
    .A(_00552_),
    .B(net6788));
 sg13g2_nand2_1 _26941_ (.Y(_13329_),
    .A(net7344),
    .B(net7318));
 sg13g2_o21ai_1 _26942_ (.B1(_13329_),
    .Y(_13330_),
    .A1(net6609),
    .A2(net7102));
 sg13g2_or2_1 _26943_ (.X(_13331_),
    .B(_13326_),
    .A(net7443));
 sg13g2_o21ai_1 _26944_ (.B1(_13328_),
    .Y(_13332_),
    .A1(net6784),
    .A2(_13330_));
 sg13g2_nand2_1 _26945_ (.Y(_13333_),
    .A(_00551_),
    .B(net6783));
 sg13g2_nand2_1 _26946_ (.Y(_13334_),
    .A(net7346),
    .B(net7318));
 sg13g2_o21ai_1 _26947_ (.B1(_13334_),
    .Y(_13335_),
    .A1(net6611),
    .A2(net7102));
 sg13g2_o21ai_1 _26948_ (.B1(_13333_),
    .Y(_13336_),
    .A1(net6784),
    .A2(_13335_));
 sg13g2_nand2_1 _26949_ (.Y(_13337_),
    .A(_00550_),
    .B(net6786));
 sg13g2_nor2_1 _26950_ (.A(_02549_),
    .B(net7042),
    .Y(_13338_));
 sg13g2_a21oi_1 _26951_ (.A1(net6612),
    .A2(net7042),
    .Y(_13339_),
    .B1(_13338_));
 sg13g2_o21ai_1 _26952_ (.B1(_13337_),
    .Y(_13340_),
    .A1(net6787),
    .A2(_13339_));
 sg13g2_nand2_1 _26953_ (.Y(_13341_),
    .A(_00549_),
    .B(net6791));
 sg13g2_nor2_1 _26954_ (.A(net7347),
    .B(net7044),
    .Y(_13342_));
 sg13g2_a21oi_1 _26955_ (.A1(net6614),
    .A2(net7044),
    .Y(_13343_),
    .B1(_13342_));
 sg13g2_o21ai_1 _26956_ (.B1(_13341_),
    .Y(_13344_),
    .A1(net6791),
    .A2(_13343_));
 sg13g2_nand2_1 _26957_ (.Y(_13345_),
    .A(_00548_),
    .B(net6791));
 sg13g2_nor2_1 _26958_ (.A(_02439_),
    .B(net7045),
    .Y(_13346_));
 sg13g2_a21oi_1 _26959_ (.A1(net6599),
    .A2(net7045),
    .Y(_13347_),
    .B1(_13346_));
 sg13g2_o21ai_1 _26960_ (.B1(_13345_),
    .Y(_13348_),
    .A1(net6791),
    .A2(_13347_));
 sg13g2_nand2_1 _26961_ (.Y(_13349_),
    .A(_00547_),
    .B(net6791));
 sg13g2_nand2_1 _26962_ (.Y(_13350_),
    .A(_02361_),
    .B(_04796_));
 sg13g2_o21ai_1 _26963_ (.B1(_13350_),
    .Y(_13351_),
    .A1(net6602),
    .A2(_08688_));
 sg13g2_o21ai_1 _26964_ (.B1(_13331_),
    .Y(_13352_),
    .A1(net7421),
    .A2(_13290_));
 sg13g2_o21ai_1 _26965_ (.B1(_13349_),
    .Y(_13353_),
    .A1(net6791),
    .A2(_13351_));
 sg13g2_nand2_1 _26966_ (.Y(_13354_),
    .A(_00546_),
    .B(net6791));
 sg13g2_nor2_1 _26967_ (.A(_02283_),
    .B(net7045),
    .Y(_13355_));
 sg13g2_nor4_1 _26968_ (.A(_13112_),
    .B(_13128_),
    .C(_13254_),
    .D(_13352_),
    .Y(_13356_));
 sg13g2_a21oi_1 _26969_ (.A1(net6621),
    .A2(net7045),
    .Y(_13357_),
    .B1(_13355_));
 sg13g2_or4_1 _26970_ (.A(_13112_),
    .B(_13128_),
    .C(_13254_),
    .D(_13352_),
    .X(_13358_));
 sg13g2_o21ai_1 _26971_ (.B1(_13354_),
    .Y(_13359_),
    .A1(net6791),
    .A2(_13357_));
 sg13g2_nand2_1 _26972_ (.Y(_13360_),
    .A(_00545_),
    .B(net6783));
 sg13g2_nor2_1 _26973_ (.A(net7348),
    .B(net7042),
    .Y(_13361_));
 sg13g2_a21oi_1 _26974_ (.A1(net6623),
    .A2(net7042),
    .Y(_13362_),
    .B1(_13361_));
 sg13g2_o21ai_1 _26975_ (.B1(_13360_),
    .Y(_13363_),
    .A1(net6783),
    .A2(_13362_));
 sg13g2_nand2_1 _26976_ (.Y(_13364_),
    .A(_00544_),
    .B(net6792));
 sg13g2_nand2_1 _26977_ (.Y(_13365_),
    .A(_09252_),
    .B(_04796_));
 sg13g2_o21ai_1 _26978_ (.B1(_13365_),
    .Y(_13366_),
    .A1(net6743),
    .A2(_08688_));
 sg13g2_nand2b_1 _26979_ (.Y(_13367_),
    .B(net8002),
    .A_N(_01636_));
 sg13g2_o21ai_1 _26980_ (.B1(_13364_),
    .Y(_13368_),
    .A1(net6792),
    .A2(_13366_));
 sg13g2_nor4_1 _26981_ (.A(net8017),
    .B(_08659_),
    .C(_08759_),
    .D(_08902_),
    .Y(_13369_));
 sg13g2_o21ai_1 _26982_ (.B1(_13367_),
    .Y(_13370_),
    .A1(_01649_),
    .A2(net7481));
 sg13g2_o21ai_1 _26983_ (.B1(_08660_),
    .Y(_13371_),
    .A1(_05162_),
    .A2(_13369_));
 sg13g2_mux2_1 _26984_ (.A0(net7997),
    .A1(net8010),
    .S(_08658_),
    .X(_13372_));
 sg13g2_nor3_1 _26985_ (.A(net8015),
    .B(net6395),
    .C(net6852),
    .Y(_13373_));
 sg13g2_a21o_1 _26986_ (.A2(net6852),
    .A1(net8003),
    .B1(_13373_),
    .X(_13374_));
 sg13g2_nand2_1 _26987_ (.Y(_13375_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_valid ),
    .B(net6852));
 sg13g2_a21oi_1 _26988_ (.A1(net7629),
    .A2(net6395),
    .Y(_13376_),
    .B1(net7993));
 sg13g2_a221oi_1 _26989_ (.B2(_00541_),
    .C1(_13370_),
    .B1(_13358_),
    .A1(_09275_),
    .Y(_13377_),
    .A2(_12791_));
 sg13g2_o21ai_1 _26990_ (.B1(_13375_),
    .Y(_13378_),
    .A1(net6852),
    .A2(_13376_));
 sg13g2_o21ai_1 _26991_ (.B1(net6784),
    .Y(_13379_),
    .A1(_05174_),
    .A2(_08658_));
 sg13g2_nor4_1 _26992_ (.A(_05162_),
    .B(net8017),
    .C(_08759_),
    .D(_08902_),
    .Y(_13380_));
 sg13g2_mux2_1 _26993_ (.A0(net8010),
    .A1(_13380_),
    .S(_08658_),
    .X(_13381_));
 sg13g2_nand2_1 _26994_ (.Y(_13382_),
    .A(net8015),
    .B(net6852));
 sg13g2_o21ai_1 _26995_ (.B1(_13382_),
    .Y(_13383_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.div_valid ),
    .A2(net6852));
 sg13g2_nand2_1 _26996_ (.Y(_13384_),
    .A(_06767_),
    .B(_08706_));
 sg13g2_mux2_1 _26997_ (.A0(_03818_),
    .A1(net8016),
    .S(_13384_),
    .X(_13385_));
 sg13g2_nand2_1 _26998_ (.Y(_13386_),
    .A(_00537_),
    .B(_13384_));
 sg13g2_nor2_1 _26999_ (.A(net7376),
    .B(_13377_),
    .Y(_13387_));
 sg13g2_o21ai_1 _27000_ (.B1(_13386_),
    .Y(_13388_),
    .A1(_00004_),
    .A2(_13384_));
 sg13g2_mux2_1 _27001_ (.A0(_00537_),
    .A1(_00536_),
    .S(_13384_),
    .X(_13389_));
 sg13g2_a21oi_1 _27002_ (.A1(net6917),
    .A2(_12819_),
    .Y(_13390_),
    .B1(_13387_));
 sg13g2_a21oi_1 _27003_ (.A1(_00536_),
    .A2(_03816_),
    .Y(_13391_),
    .B1(net8016));
 sg13g2_mux2_1 _27004_ (.A0(_13391_),
    .A1(_00004_),
    .S(_13384_),
    .X(_13392_));
 sg13g2_nor2_1 _27005_ (.A(net8003),
    .B(_08685_),
    .Y(_13393_));
 sg13g2_a21oi_1 _27006_ (.A1(_08938_),
    .A2(_13393_),
    .Y(_13394_),
    .B1(_08659_));
 sg13g2_and2_1 _27007_ (.A(_08663_),
    .B(_13393_),
    .X(_13395_));
 sg13g2_nand4_1 _27008_ (.B(_08772_),
    .C(_08901_),
    .A(net8017),
    .Y(_13396_),
    .D(_13395_));
 sg13g2_o21ai_1 _27009_ (.B1(_13396_),
    .Y(_13397_),
    .A1(net8017),
    .A2(_13394_));
 sg13g2_inv_1 _27010_ (.Y(_13398_),
    .A(_13397_));
 sg13g2_a21o_1 _27011_ (.A2(_13393_),
    .A1(_08937_),
    .B1(_08659_),
    .X(_13399_));
 sg13g2_a22oi_1 _27012_ (.Y(_13400_),
    .B1(_13399_),
    .B2(_05199_),
    .A2(_13395_),
    .A1(_09168_));
 sg13g2_a21oi_1 _27013_ (.A1(_08773_),
    .A2(_13393_),
    .Y(_13401_),
    .B1(_08659_));
 sg13g2_o21ai_1 _27014_ (.B1(_13390_),
    .Y(_13402_),
    .A1(_08228_),
    .A2(_12819_));
 sg13g2_nand3_1 _27015_ (.B(_08772_),
    .C(_13395_),
    .A(_00533_),
    .Y(_13403_));
 sg13g2_inv_1 _27016_ (.Y(_13404_),
    .A(_13405_));
 sg13g2_o21ai_1 _27017_ (.B1(_13403_),
    .Y(_13405_),
    .A1(_00533_),
    .A2(_13401_));
 sg13g2_nand2_1 _27018_ (.Y(_13406_),
    .A(net8021),
    .B(_13393_));
 sg13g2_o21ai_1 _27019_ (.B1(_08777_),
    .Y(_13407_),
    .A1(_08797_),
    .A2(_08819_));
 sg13g2_a21oi_1 _27020_ (.A1(_08658_),
    .A2(_13406_),
    .Y(_13408_),
    .B1(net8019));
 sg13g2_nor2b_1 _27021_ (.A(_08743_),
    .B_N(_13395_),
    .Y(_13409_));
 sg13g2_and2_1 _27022_ (.A(_08851_),
    .B(_13407_),
    .X(_13410_));
 sg13g2_nor2_1 _27023_ (.A(_13408_),
    .B(_13409_),
    .Y(_13411_));
 sg13g2_nor2_1 _27024_ (.A(net8022),
    .B(_08663_),
    .Y(_13412_));
 sg13g2_a21oi_1 _27025_ (.A1(net8022),
    .A2(_13395_),
    .Y(_13413_),
    .B1(_13412_));
 sg13g2_nor3_1 _27026_ (.A(net8015),
    .B(net6852),
    .C(_08690_),
    .Y(_13414_));
 sg13g2_nand2_1 _27027_ (.Y(_13415_),
    .A(net6395),
    .B(_13414_));
 sg13g2_o21ai_1 _27028_ (.B1(_13415_),
    .Y(_13416_),
    .A1(_05213_),
    .A2(_13414_));
 sg13g2_inv_1 _27029_ (.Y(_13417_),
    .A(_13418_));
 sg13g2_nand3b_1 _27030_ (.B(net6768),
    .C(_07660_),
    .Y(_13418_),
    .A_N(_07085_));
 sg13g2_nand4_1 _27031_ (.B(_06890_),
    .C(_06894_),
    .A(_06885_),
    .Y(_13419_),
    .D(_06914_));
 sg13g2_nor2_1 _27032_ (.A(_06887_),
    .B(_13419_),
    .Y(_13420_));
 sg13g2_nor3_1 _27033_ (.A(_06884_),
    .B(_06936_),
    .C(_06937_),
    .Y(_13421_));
 sg13g2_nand2_1 _27034_ (.Y(_13422_),
    .A(_06894_),
    .B(_13421_));
 sg13g2_nor2_1 _27035_ (.A(_06935_),
    .B(_13422_),
    .Y(_13423_));
 sg13g2_and2_1 _27036_ (.A(_10063_),
    .B(_13423_),
    .X(_13424_));
 sg13g2_nand4_1 _27037_ (.B(_06885_),
    .C(_06911_),
    .A(net6932),
    .Y(_13425_),
    .D(_06913_));
 sg13g2_a21oi_1 _27038_ (.A1(_06889_),
    .A2(_06953_),
    .Y(_13426_),
    .B1(_13425_));
 sg13g2_nor2_1 _27039_ (.A(_13417_),
    .B(_13424_),
    .Y(_13427_));
 sg13g2_nand2b_1 _27040_ (.Y(_13428_),
    .B(_13427_),
    .A_N(_00530_));
 sg13g2_o21ai_1 _27041_ (.B1(_13428_),
    .Y(_13429_),
    .A1(net313),
    .A2(_13418_));
 sg13g2_nor3_1 _27042_ (.A(net7021),
    .B(net7415),
    .C(_10917_),
    .Y(_13430_));
 sg13g2_a21oi_1 _27043_ (.A1(net7021),
    .A2(net7310),
    .Y(_13431_),
    .B1(_13430_));
 sg13g2_a21oi_1 _27044_ (.A1(net6546),
    .A2(net6459),
    .Y(_13432_),
    .B1(_13429_));
 sg13g2_nand2b_1 _27045_ (.Y(_13433_),
    .B(net6461),
    .A_N(_00529_));
 sg13g2_o21ai_1 _27046_ (.B1(_13433_),
    .Y(_13434_),
    .A1(net312),
    .A2(_13418_));
 sg13g2_nor3_1 _27047_ (.A(_03695_),
    .B(_06968_),
    .C(_10954_),
    .Y(_13435_));
 sg13g2_a21oi_1 _27048_ (.A1(_03695_),
    .A2(_06970_),
    .Y(_13436_),
    .B1(_13435_));
 sg13g2_a21oi_1 _27049_ (.A1(net6546),
    .A2(_13436_),
    .Y(_13437_),
    .B1(_13434_));
 sg13g2_nand2b_1 _27050_ (.Y(_13438_),
    .B(net6462),
    .A_N(_00528_));
 sg13g2_o21ai_1 _27051_ (.B1(_13438_),
    .Y(_13439_),
    .A1(net311),
    .A2(net6729));
 sg13g2_nor3_1 _27052_ (.A(_03812_),
    .B(net7414),
    .C(_10125_),
    .Y(_13440_));
 sg13g2_a21oi_1 _27053_ (.A1(_03812_),
    .A2(net7312),
    .Y(_13441_),
    .B1(_13440_));
 sg13g2_a21oi_1 _27054_ (.A1(net6545),
    .A2(net6158),
    .Y(_13442_),
    .B1(_13439_));
 sg13g2_nand2b_1 _27055_ (.Y(_13443_),
    .B(net6462),
    .A_N(_00527_));
 sg13g2_o21ai_1 _27056_ (.B1(_13443_),
    .Y(_13444_),
    .A1(net310),
    .A2(net6729));
 sg13g2_nor3_1 _27057_ (.A(net7006),
    .B(net7414),
    .C(_10151_),
    .Y(_13445_));
 sg13g2_a21oi_1 _27058_ (.A1(net7006),
    .A2(net7309),
    .Y(_13446_),
    .B1(_13445_));
 sg13g2_a21oi_1 _27059_ (.A1(net6545),
    .A2(net6157),
    .Y(_13447_),
    .B1(_13444_));
 sg13g2_nand2b_1 _27060_ (.Y(_13448_),
    .B(net6462),
    .A_N(_00526_));
 sg13g2_o21ai_1 _27061_ (.B1(_13448_),
    .Y(_13449_),
    .A1(net309),
    .A2(net6729));
 sg13g2_nor3_1 _27062_ (.A(net7007),
    .B(net7414),
    .C(_10195_),
    .Y(_13450_));
 sg13g2_a21oi_1 _27063_ (.A1(net7007),
    .A2(net7309),
    .Y(_13451_),
    .B1(_13450_));
 sg13g2_mux4_1 _27064_ (.S0(net7792),
    .A0(_00793_),
    .A1(_00825_),
    .A2(_00857_),
    .A3(_00892_),
    .S1(net7741),
    .X(_13452_));
 sg13g2_a21oi_1 _27065_ (.A1(net6545),
    .A2(net6154),
    .Y(_13453_),
    .B1(_13449_));
 sg13g2_nand2b_1 _27066_ (.Y(_13454_),
    .B(net6462),
    .A_N(_00525_));
 sg13g2_and2_1 _27067_ (.A(net7604),
    .B(_13452_),
    .X(_13455_));
 sg13g2_o21ai_1 _27068_ (.B1(_13454_),
    .Y(_13456_),
    .A1(net308),
    .A2(net6729));
 sg13g2_nor2_1 _27069_ (.A(_03796_),
    .B(net7414),
    .Y(_13457_));
 sg13g2_a22oi_1 _27070_ (.Y(_13458_),
    .B1(_10230_),
    .B2(_13457_),
    .A2(net7312),
    .A1(_03796_));
 sg13g2_nand2_1 _27071_ (.Y(_13459_),
    .A(net7710),
    .B(_00761_));
 sg13g2_a21oi_1 _27072_ (.A1(net6545),
    .A2(net6458),
    .Y(_13460_),
    .B1(_13456_));
 sg13g2_nand2b_1 _27073_ (.Y(_13461_),
    .B(net6460),
    .A_N(_00524_));
 sg13g2_o21ai_1 _27074_ (.B1(_13461_),
    .Y(_13462_),
    .A1(net307),
    .A2(net6730));
 sg13g2_nor3_1 _27075_ (.A(net7008),
    .B(net7414),
    .C(_10263_),
    .Y(_13463_));
 sg13g2_nand2b_1 _27076_ (.Y(_13464_),
    .B(_00629_),
    .A_N(net7710));
 sg13g2_a21oi_1 _27077_ (.A1(net7008),
    .A2(net7309),
    .Y(_13465_),
    .B1(_13463_));
 sg13g2_a21oi_1 _27078_ (.A1(net6544),
    .A2(net6153),
    .Y(_13466_),
    .B1(_13462_));
 sg13g2_nand2b_1 _27079_ (.Y(_13467_),
    .B(net6460),
    .A_N(_00523_));
 sg13g2_a21oi_1 _27080_ (.A1(_13459_),
    .A2(_13464_),
    .Y(_13468_),
    .B1(net7600));
 sg13g2_o21ai_1 _27081_ (.B1(_13467_),
    .Y(_13469_),
    .A1(net306),
    .A2(net6730));
 sg13g2_nor3_1 _27082_ (.A(_03785_),
    .B(net7414),
    .C(_10290_),
    .Y(_13470_));
 sg13g2_a21oi_1 _27083_ (.A1(_03785_),
    .A2(net7309),
    .Y(_13471_),
    .B1(_13470_));
 sg13g2_a21oi_1 _27084_ (.A1(net6544),
    .A2(net6150),
    .Y(_13472_),
    .B1(_13469_));
 sg13g2_nand2b_1 _27085_ (.Y(_13473_),
    .B(net6460),
    .A_N(_00522_));
 sg13g2_o21ai_1 _27086_ (.B1(_13473_),
    .Y(_13474_),
    .A1(net305),
    .A2(net6730));
 sg13g2_nor3_1 _27087_ (.A(_03780_),
    .B(net7414),
    .C(_10327_),
    .Y(_13475_));
 sg13g2_nand3b_1 _27088_ (.B(net7792),
    .C(_00917_),
    .Y(_13476_),
    .A_N(net7742));
 sg13g2_a21oi_1 _27089_ (.A1(_03780_),
    .A2(net7309),
    .Y(_13477_),
    .B1(_13475_));
 sg13g2_nand3b_1 _27090_ (.B(_01269_),
    .C(net7741),
    .Y(_13478_),
    .A_N(net7792));
 sg13g2_a21oi_1 _27091_ (.A1(net6544),
    .A2(net6149),
    .Y(_13479_),
    .B1(_13474_));
 sg13g2_nand2b_1 _27092_ (.Y(_13480_),
    .B(net6460),
    .A_N(_00521_));
 sg13g2_o21ai_1 _27093_ (.B1(_13480_),
    .Y(_13481_),
    .A1(net304),
    .A2(net6730));
 sg13g2_nor3_1 _27094_ (.A(net7010),
    .B(net7416),
    .C(_10361_),
    .Y(_13482_));
 sg13g2_a21oi_1 _27095_ (.A1(_13476_),
    .A2(_13478_),
    .Y(_13483_),
    .B1(net7598));
 sg13g2_a21oi_1 _27096_ (.A1(net7010),
    .A2(net7311),
    .Y(_13484_),
    .B1(_13482_));
 sg13g2_a21oi_1 _27097_ (.A1(net6544),
    .A2(net6147),
    .Y(_13485_),
    .B1(_13481_));
 sg13g2_nand2b_1 _27098_ (.Y(_13486_),
    .B(net6461),
    .A_N(_00520_));
 sg13g2_o21ai_1 _27099_ (.B1(_13486_),
    .Y(_13487_),
    .A1(net303),
    .A2(net6731));
 sg13g2_nor3_1 _27100_ (.A(net7011),
    .B(net7416),
    .C(_10406_),
    .Y(_13488_));
 sg13g2_nor4_1 _27101_ (.A(net7690),
    .B(_13455_),
    .C(_13468_),
    .D(_13483_),
    .Y(_13489_));
 sg13g2_a21oi_1 _27102_ (.A1(net7011),
    .A2(net7311),
    .Y(_13490_),
    .B1(_13488_));
 sg13g2_a21oi_1 _27103_ (.A1(_13424_),
    .A2(net6145),
    .Y(_13491_),
    .B1(_13487_));
 sg13g2_nand2b_1 _27104_ (.Y(_13492_),
    .B(net6461),
    .A_N(_00519_));
 sg13g2_o21ai_1 _27105_ (.B1(_13492_),
    .Y(_13493_),
    .A1(net302),
    .A2(net6731));
 sg13g2_nor3_1 _27106_ (.A(_03765_),
    .B(net7414),
    .C(_10441_),
    .Y(_13494_));
 sg13g2_a21oi_1 _27107_ (.A1(_03765_),
    .A2(net7309),
    .Y(_13495_),
    .B1(_13494_));
 sg13g2_a21oi_1 _27108_ (.A1(_13424_),
    .A2(net6144),
    .Y(_13496_),
    .B1(_13493_));
 sg13g2_nand2b_1 _27109_ (.Y(_13497_),
    .B(net6460),
    .A_N(_00518_));
 sg13g2_o21ai_1 _27110_ (.B1(_13497_),
    .Y(_13498_),
    .A1(net301),
    .A2(net6730));
 sg13g2_nor3_1 _27111_ (.A(_03760_),
    .B(net7416),
    .C(_10485_),
    .Y(_13499_));
 sg13g2_mux2_1 _27112_ (.A0(_00665_),
    .A1(_00697_),
    .S(net7792),
    .X(_13500_));
 sg13g2_a21oi_1 _27113_ (.A1(_03760_),
    .A2(net7311),
    .Y(_13501_),
    .B1(_13499_));
 sg13g2_a21oi_1 _27114_ (.A1(net6544),
    .A2(net6143),
    .Y(_13502_),
    .B1(_13498_));
 sg13g2_nand2b_1 _27115_ (.Y(_13503_),
    .B(net6460),
    .A_N(_00517_));
 sg13g2_o21ai_1 _27116_ (.B1(_13503_),
    .Y(_13504_),
    .A1(net300),
    .A2(net6730));
 sg13g2_nor3_1 _27117_ (.A(_03755_),
    .B(net7417),
    .C(_10517_),
    .Y(_13505_));
 sg13g2_a21oi_1 _27118_ (.A1(_03755_),
    .A2(net7311),
    .Y(_13506_),
    .B1(_13505_));
 sg13g2_a21oi_1 _27119_ (.A1(net6544),
    .A2(_13506_),
    .Y(_13507_),
    .B1(_13504_));
 sg13g2_nand2b_1 _27120_ (.Y(_13508_),
    .B(net6460),
    .A_N(_00516_));
 sg13g2_o21ai_1 _27121_ (.B1(_13508_),
    .Y(_13509_),
    .A1(net299),
    .A2(net6730));
 sg13g2_nor3_1 _27122_ (.A(net7012),
    .B(net7415),
    .C(_10562_),
    .Y(_13510_));
 sg13g2_a21oi_1 _27123_ (.A1(net7012),
    .A2(net7310),
    .Y(_13511_),
    .B1(_13510_));
 sg13g2_a21oi_1 _27124_ (.A1(net6544),
    .A2(net6141),
    .Y(_13512_),
    .B1(_13509_));
 sg13g2_nand2b_1 _27125_ (.Y(_13513_),
    .B(net6462),
    .A_N(_00515_));
 sg13g2_o21ai_1 _27126_ (.B1(_13513_),
    .Y(_13514_),
    .A1(net298),
    .A2(net6729));
 sg13g2_nor3_1 _27127_ (.A(net7013),
    .B(net7415),
    .C(_10604_),
    .Y(_13515_));
 sg13g2_a21oi_1 _27128_ (.A1(net7013),
    .A2(net7310),
    .Y(_13516_),
    .B1(_13515_));
 sg13g2_a21oi_1 _27129_ (.A1(net6545),
    .A2(net6140),
    .Y(_13517_),
    .B1(_13514_));
 sg13g2_nand2b_1 _27130_ (.Y(_13518_),
    .B(net6460),
    .A_N(_00514_));
 sg13g2_a221oi_1 _27131_ (.B2(net7516),
    .C1(net7694),
    .B1(_13500_),
    .A1(_00729_),
    .Y(_13519_),
    .A2(net7595));
 sg13g2_o21ai_1 _27132_ (.B1(_13518_),
    .Y(_13520_),
    .A1(net297),
    .A2(net6730));
 sg13g2_nor3_1 _27133_ (.A(net7014),
    .B(net7415),
    .C(_10641_),
    .Y(_13521_));
 sg13g2_a21oi_1 _27134_ (.A1(net7014),
    .A2(net7310),
    .Y(_13522_),
    .B1(_13521_));
 sg13g2_a21oi_1 _27135_ (.A1(net6544),
    .A2(net6138),
    .Y(_13523_),
    .B1(_13520_));
 sg13g2_nand2b_1 _27136_ (.Y(_13524_),
    .B(net6461),
    .A_N(_00513_));
 sg13g2_o21ai_1 _27137_ (.B1(_13524_),
    .Y(_13525_),
    .A1(net296),
    .A2(net6731));
 sg13g2_nor3_1 _27138_ (.A(net7015),
    .B(net7416),
    .C(_10679_),
    .Y(_13526_));
 sg13g2_a21oi_1 _27139_ (.A1(net7015),
    .A2(net7311),
    .Y(_13527_),
    .B1(_13526_));
 sg13g2_a21oi_1 _27140_ (.A1(net6546),
    .A2(_13527_),
    .Y(_13528_),
    .B1(_13525_));
 sg13g2_nand2b_1 _27141_ (.Y(_13529_),
    .B(net6461),
    .A_N(_00512_));
 sg13g2_o21ai_1 _27142_ (.B1(_13529_),
    .Y(_13530_),
    .A1(net295),
    .A2(net6731));
 sg13g2_o21ai_1 _27143_ (.B1(_03729_),
    .Y(_13531_),
    .A1(net7417),
    .A2(_10722_));
 sg13g2_o21ai_1 _27144_ (.B1(_13531_),
    .Y(_13532_),
    .A1(_03729_),
    .A2(net7312));
 sg13g2_a21oi_1 _27145_ (.A1(_13424_),
    .A2(net6543),
    .Y(_13533_),
    .B1(_13530_));
 sg13g2_nand2b_1 _27146_ (.Y(_13534_),
    .B(net6461),
    .A_N(_00511_));
 sg13g2_o21ai_1 _27147_ (.B1(_13534_),
    .Y(_13535_),
    .A1(net294),
    .A2(_13418_));
 sg13g2_nor2_1 _27148_ (.A(net7016),
    .B(net7415),
    .Y(_13536_));
 sg13g2_a22oi_1 _27149_ (.Y(_13537_),
    .B1(_10754_),
    .B2(_13536_),
    .A2(net7310),
    .A1(net7016));
 sg13g2_a21oi_1 _27150_ (.A1(net6546),
    .A2(net6542),
    .Y(_13538_),
    .B1(_13535_));
 sg13g2_nand2b_1 _27151_ (.Y(_13539_),
    .B(net6462),
    .A_N(_00510_));
 sg13g2_o21ai_1 _27152_ (.B1(_13539_),
    .Y(_13540_),
    .A1(net293),
    .A2(net6729));
 sg13g2_nor3_1 _27153_ (.A(net7017),
    .B(net7415),
    .C(_10783_),
    .Y(_13541_));
 sg13g2_a21oi_1 _27154_ (.A1(net7017),
    .A2(net7310),
    .Y(_13542_),
    .B1(_13541_));
 sg13g2_a21oi_1 _27155_ (.A1(net6545),
    .A2(net6136),
    .Y(_13543_),
    .B1(_13540_));
 sg13g2_nand2b_1 _27156_ (.Y(_13544_),
    .B(net6462),
    .A_N(_00509_));
 sg13g2_o21ai_1 _27157_ (.B1(_13544_),
    .Y(_13545_),
    .A1(net292),
    .A2(net6729));
 sg13g2_nor3_1 _27158_ (.A(net7018),
    .B(net7415),
    .C(_10817_),
    .Y(_13546_));
 sg13g2_a21oi_1 _27159_ (.A1(net7018),
    .A2(net7310),
    .Y(_13547_),
    .B1(_13546_));
 sg13g2_a21oi_1 _27160_ (.A1(net6545),
    .A2(net6456),
    .Y(_13548_),
    .B1(_13545_));
 sg13g2_nand2b_1 _27161_ (.Y(_13549_),
    .B(net6462),
    .A_N(_00508_));
 sg13g2_mux4_1 _27162_ (.S0(net7792),
    .A0(_00927_),
    .A1(_00963_),
    .A2(_00998_),
    .A3(_01033_),
    .S1(net7741),
    .X(_13550_));
 sg13g2_o21ai_1 _27163_ (.B1(_13549_),
    .Y(_13551_),
    .A1(net291),
    .A2(net6729));
 sg13g2_nor3_1 _27164_ (.A(net7019),
    .B(net7415),
    .C(_10848_),
    .Y(_13552_));
 sg13g2_a21oi_1 _27165_ (.A1(net7019),
    .A2(net7310),
    .Y(_13553_),
    .B1(_13552_));
 sg13g2_a21oi_1 _27166_ (.A1(net6545),
    .A2(net6134),
    .Y(_13554_),
    .B1(_13551_));
 sg13g2_nand2b_1 _27167_ (.Y(_13555_),
    .B(net6461),
    .A_N(_00507_));
 sg13g2_o21ai_1 _27168_ (.B1(_13555_),
    .Y(_13556_),
    .A1(net290),
    .A2(_13418_));
 sg13g2_nor3_1 _27169_ (.A(net7020),
    .B(_06968_),
    .C(_10873_),
    .Y(_13557_));
 sg13g2_o21ai_1 _27170_ (.B1(net7707),
    .Y(_13558_),
    .A1(net7531),
    .A2(_13550_));
 sg13g2_a21oi_1 _27171_ (.A1(net7020),
    .A2(net7309),
    .Y(_13559_),
    .B1(_13557_));
 sg13g2_a21oi_1 _27172_ (.A1(net6546),
    .A2(net6455),
    .Y(_13560_),
    .B1(_13556_));
 sg13g2_nand2_1 _27173_ (.Y(_13561_),
    .A(_06899_),
    .B(net7437));
 sg13g2_o21ai_1 _27174_ (.B1(_13561_),
    .Y(_13562_),
    .A1(_02235_),
    .A2(_06899_));
 sg13g2_a21oi_1 _27175_ (.A1(_06906_),
    .A2(net7437),
    .Y(_13563_),
    .B1(_07089_));
 sg13g2_inv_1 _27176_ (.Y(_13564_),
    .A(_13563_));
 sg13g2_a21oi_1 _27177_ (.A1(_02226_),
    .A2(_13562_),
    .Y(_13565_),
    .B1(_13564_));
 sg13g2_a21o_1 _27178_ (.A2(_13562_),
    .A1(_02226_),
    .B1(_13564_),
    .X(_13566_));
 sg13g2_nor3_1 _27179_ (.A(net7984),
    .B(_02235_),
    .C(_06899_),
    .Y(_13567_));
 sg13g2_inv_1 _27180_ (.Y(_13568_),
    .A(_13569_));
 sg13g2_or2_1 _27181_ (.X(_13569_),
    .B(_13567_),
    .A(_06909_));
 sg13g2_nor2_1 _27182_ (.A(\cs_registers_i.debug_mode_i ),
    .B(_13569_),
    .Y(_13570_));
 sg13g2_nand2_1 _27183_ (.Y(_13571_),
    .A(_02226_),
    .B(_13568_));
 sg13g2_nor2_1 _27184_ (.A(_13565_),
    .B(_13571_),
    .Y(_13572_));
 sg13g2_nand2_1 _27185_ (.Y(_13573_),
    .A(_13566_),
    .B(_13570_));
 sg13g2_nand2_1 _27186_ (.Y(_13574_),
    .A(net6675),
    .B(_13420_));
 sg13g2_nand3_1 _27187_ (.B(_09551_),
    .C(_13423_),
    .A(_09549_),
    .Y(_13575_));
 sg13g2_a21oi_1 _27188_ (.A1(net6675),
    .A2(_13420_),
    .Y(_13576_),
    .B1(net6668));
 sg13g2_o21ai_1 _27189_ (.B1(_06903_),
    .Y(_13577_),
    .A1(_06782_),
    .A2(_06895_));
 sg13g2_and3_1 _27190_ (.X(_13578_),
    .A(net7437),
    .B(_13572_),
    .C(_13577_));
 sg13g2_and2_1 _27191_ (.A(\id_stage_i.controller_i.illegal_insn_q ),
    .B(_06902_),
    .X(_13579_));
 sg13g2_o21ai_1 _27192_ (.B1(_13489_),
    .Y(_13580_),
    .A1(_13519_),
    .A2(_13558_));
 sg13g2_mux2_1 _27193_ (.A0(net7666),
    .A1(_01885_),
    .S(net7933),
    .X(_13581_));
 sg13g2_a22oi_1 _27194_ (.Y(_13582_),
    .B1(_13579_),
    .B2(_13581_),
    .A2(_07762_),
    .A1(_01980_));
 sg13g2_nand3_1 _27195_ (.B(_01928_),
    .C(\id_stage_i.controller_i.instr_fetch_err_plus2_i ),
    .A(_01939_),
    .Y(_13583_));
 sg13g2_nor2_1 _27196_ (.A(_07622_),
    .B(_13583_),
    .Y(_13584_));
 sg13g2_and2_1 _27197_ (.A(_01943_),
    .B(_13584_),
    .X(_13585_));
 sg13g2_nand2_1 _27198_ (.Y(_13586_),
    .A(_01944_),
    .B(_13585_));
 sg13g2_nand3_1 _27199_ (.B(_01944_),
    .C(_13585_),
    .A(_01945_),
    .Y(_13587_));
 sg13g2_nor2_1 _27200_ (.A(_07450_),
    .B(_13587_),
    .Y(_13588_));
 sg13g2_nand2_1 _27201_ (.Y(_13589_),
    .A(_01947_),
    .B(_13588_));
 sg13g2_xor2_1 _27202_ (.B(_13589_),
    .A(_01948_),
    .X(_13590_));
 sg13g2_o21ai_1 _27203_ (.B1(_13582_),
    .Y(_13591_),
    .A1(net7624),
    .A2(_13590_));
 sg13g2_nand2b_1 _27204_ (.Y(_13592_),
    .B(_13431_),
    .A_N(_13574_));
 sg13g2_a22oi_1 _27205_ (.Y(_13593_),
    .B1(_13592_),
    .B2(net6655),
    .A2(_13591_),
    .A1(net6643));
 sg13g2_a21oi_1 _27206_ (.A1(_05288_),
    .A2(_13576_),
    .Y(_13594_),
    .B1(_13593_));
 sg13g2_mux2_1 _27207_ (.A0(net7671),
    .A1(_01884_),
    .S(net7933),
    .X(_13595_));
 sg13g2_nand2_1 _27208_ (.Y(_13596_),
    .A(_01979_),
    .B(net6988));
 sg13g2_xor2_1 _27209_ (.B(_13588_),
    .A(_01947_),
    .X(_13597_));
 sg13g2_a22oi_1 _27210_ (.Y(_13598_),
    .B1(_13597_),
    .B2(_06901_),
    .A2(_13595_),
    .A1(net7419));
 sg13g2_nand2_1 _27211_ (.Y(_13599_),
    .A(_13596_),
    .B(_13598_));
 sg13g2_nand2b_1 _27212_ (.Y(_13600_),
    .B(net6159),
    .A_N(_13574_));
 sg13g2_a22oi_1 _27213_ (.Y(_13601_),
    .B1(_13600_),
    .B2(net6653),
    .A2(_13599_),
    .A1(net6644));
 sg13g2_a21oi_1 _27214_ (.A1(_05289_),
    .A2(net6536),
    .Y(_13602_),
    .B1(_13601_));
 sg13g2_nand2_1 _27215_ (.Y(_13603_),
    .A(_01978_),
    .B(net6988));
 sg13g2_xnor2_1 _27216_ (.Y(_13604_),
    .A(_01946_),
    .B(_13587_));
 sg13g2_nand2_1 _27217_ (.Y(_13605_),
    .A(_01883_),
    .B(net7933));
 sg13g2_o21ai_1 _27218_ (.B1(_13605_),
    .Y(_13606_),
    .A1(_08510_),
    .A2(net7936));
 sg13g2_a22oi_1 _27219_ (.Y(_13607_),
    .B1(_13606_),
    .B2(net7419),
    .A2(_13604_),
    .A1(_06901_));
 sg13g2_nand2_1 _27220_ (.Y(_13608_),
    .A(_13603_),
    .B(_13607_));
 sg13g2_nor3_1 _27221_ (.A(net7023),
    .B(net7416),
    .C(_09670_),
    .Y(_13609_));
 sg13g2_a21oi_1 _27222_ (.A1(net7023),
    .A2(net7311),
    .Y(_13610_),
    .B1(_13609_));
 sg13g2_nand2b_1 _27223_ (.Y(_13611_),
    .B(_13610_),
    .A_N(net6539));
 sg13g2_a22oi_1 _27224_ (.Y(_13612_),
    .B1(_13611_),
    .B2(net6656),
    .A2(_13608_),
    .A1(net6641));
 sg13g2_a21oi_1 _27225_ (.A1(_05292_),
    .A2(net6536),
    .Y(_13613_),
    .B1(_13612_));
 sg13g2_nand2_1 _27226_ (.Y(_13614_),
    .A(_01977_),
    .B(net6988));
 sg13g2_nand2_1 _27227_ (.Y(_13615_),
    .A(_01882_),
    .B(net7933));
 sg13g2_o21ai_1 _27228_ (.B1(_13615_),
    .Y(_13616_),
    .A1(_08533_),
    .A2(net7936));
 sg13g2_xnor2_1 _27229_ (.Y(_13617_),
    .A(_01945_),
    .B(_13586_));
 sg13g2_a22oi_1 _27230_ (.Y(_13618_),
    .B1(_13617_),
    .B2(_06901_),
    .A2(_13616_),
    .A1(net7420));
 sg13g2_nand2_1 _27231_ (.Y(_13619_),
    .A(_13614_),
    .B(_13618_));
 sg13g2_nor3_1 _27232_ (.A(net7024),
    .B(net7416),
    .C(_09769_),
    .Y(_13620_));
 sg13g2_a21oi_1 _27233_ (.A1(net7024),
    .A2(net7312),
    .Y(_13621_),
    .B1(_13620_));
 sg13g2_nand2b_1 _27234_ (.Y(_13622_),
    .B(_13621_),
    .A_N(net6540));
 sg13g2_mux4_1 _27235_ (.S0(net7799),
    .A0(_01068_),
    .A1(_01103_),
    .A2(_01139_),
    .A3(_01174_),
    .S1(net7746),
    .X(_13623_));
 sg13g2_a22oi_1 _27236_ (.Y(_13624_),
    .B1(_13622_),
    .B2(net6656),
    .A2(_13619_),
    .A1(net6641));
 sg13g2_a21oi_1 _27237_ (.A1(_05296_),
    .A2(net6536),
    .Y(_13625_),
    .B1(_13624_));
 sg13g2_nand2_1 _27238_ (.Y(_13626_),
    .A(_01976_),
    .B(net6987));
 sg13g2_xor2_1 _27239_ (.B(_13585_),
    .A(_01944_),
    .X(_13627_));
 sg13g2_nand2_1 _27240_ (.Y(_13628_),
    .A(_01881_),
    .B(net7934));
 sg13g2_nand2b_1 _27241_ (.Y(_13629_),
    .B(_08387_),
    .A_N(_13623_));
 sg13g2_o21ai_1 _27242_ (.B1(_13628_),
    .Y(_13630_),
    .A1(_08563_),
    .A2(net7935));
 sg13g2_a22oi_1 _27243_ (.Y(_13631_),
    .B1(_13630_),
    .B2(net7420),
    .A2(_13627_),
    .A1(_06901_));
 sg13g2_nand2_1 _27244_ (.Y(_13632_),
    .A(_13626_),
    .B(_13631_));
 sg13g2_nor3_1 _27245_ (.A(net7025),
    .B(net7417),
    .C(_09826_),
    .Y(_13633_));
 sg13g2_a21oi_1 _27246_ (.A1(net7025),
    .A2(net7312),
    .Y(_13634_),
    .B1(_13633_));
 sg13g2_nand2b_1 _27247_ (.Y(_13635_),
    .B(net6533),
    .A_N(net6540));
 sg13g2_a22oi_1 _27248_ (.Y(_13636_),
    .B1(_13635_),
    .B2(net6653),
    .A2(_13632_),
    .A1(net6644));
 sg13g2_a21oi_1 _27249_ (.A1(_05301_),
    .A2(net6535),
    .Y(_13637_),
    .B1(_13636_));
 sg13g2_nand2_1 _27250_ (.Y(_13638_),
    .A(_01975_),
    .B(net6985));
 sg13g2_xor2_1 _27251_ (.B(_13584_),
    .A(_01943_),
    .X(_13639_));
 sg13g2_mux2_1 _27252_ (.A0(_01912_),
    .A1(_01880_),
    .S(net7934),
    .X(_13640_));
 sg13g2_a22oi_1 _27253_ (.Y(_13641_),
    .B1(_13640_),
    .B2(net7420),
    .A2(_13639_),
    .A1(_06901_));
 sg13g2_nand2_1 _27254_ (.Y(_13642_),
    .A(_13638_),
    .B(_13641_));
 sg13g2_nand2_1 _27255_ (.Y(_13643_),
    .A(_13578_),
    .B(_13642_));
 sg13g2_nor3_1 _27256_ (.A(net7026),
    .B(_06968_),
    .C(_09899_),
    .Y(_13644_));
 sg13g2_inv_1 _27257_ (.Y(_13645_),
    .A(_13646_));
 sg13g2_a21o_1 _27258_ (.A2(_06970_),
    .A1(net7026),
    .B1(_13644_),
    .X(_13646_));
 sg13g2_o21ai_1 _27259_ (.B1(net6656),
    .Y(_13647_),
    .A1(net6539),
    .A2(_13646_));
 sg13g2_a22oi_1 _27260_ (.Y(_13648_),
    .B1(_13643_),
    .B2(_13647_),
    .A2(net6536),
    .A1(_05306_));
 sg13g2_and2_1 _27261_ (.A(_07622_),
    .B(_13583_),
    .X(_13649_));
 sg13g2_nor3_1 _27262_ (.A(net7625),
    .B(_13584_),
    .C(_13649_),
    .Y(_13650_));
 sg13g2_nand2_1 _27263_ (.Y(_13651_),
    .A(_01879_),
    .B(net7934));
 sg13g2_o21ai_1 _27264_ (.B1(_13651_),
    .Y(_13652_),
    .A1(_08622_),
    .A2(net7936));
 sg13g2_a221oi_1 _27265_ (.B2(_13652_),
    .C1(_13650_),
    .B1(net7420),
    .A1(_01974_),
    .Y(_13653_),
    .A2(net6985));
 sg13g2_nand2b_1 _27266_ (.Y(_13654_),
    .B(_13578_),
    .A_N(_13653_));
 sg13g2_nor3_1 _27267_ (.A(net7027),
    .B(_06968_),
    .C(_09599_),
    .Y(_13655_));
 sg13g2_inv_1 _27268_ (.Y(_13656_),
    .A(_13657_));
 sg13g2_a21o_1 _27269_ (.A2(_06970_),
    .A1(net7027),
    .B1(_13655_),
    .X(_13657_));
 sg13g2_o21ai_1 _27270_ (.B1(net6657),
    .Y(_13658_),
    .A1(net6539),
    .A2(_13657_));
 sg13g2_a22oi_1 _27271_ (.Y(_13659_),
    .B1(_13654_),
    .B2(_13658_),
    .A2(net6536),
    .A1(_05308_));
 sg13g2_nor2b_1 _27272_ (.A(net7935),
    .B_N(_13579_),
    .Y(_13660_));
 sg13g2_a22oi_1 _27273_ (.Y(_13661_),
    .B1(net7350),
    .B2(net7677),
    .A2(net6988),
    .A1(_01973_));
 sg13g2_nand3_1 _27274_ (.B(_01947_),
    .C(_13588_),
    .A(_01948_),
    .Y(_13662_));
 sg13g2_nor2_1 _27275_ (.A(_08414_),
    .B(_13662_),
    .Y(_13663_));
 sg13g2_and4_1 _27276_ (.A(_01921_),
    .B(_01920_),
    .C(_01919_),
    .D(_13663_),
    .X(_13664_));
 sg13g2_mux4_1 _27277_ (.S0(net7799),
    .A0(_01209_),
    .A1(_01244_),
    .A2(_01279_),
    .A3(_01315_),
    .S1(net7747),
    .X(_13665_));
 sg13g2_nand2_1 _27278_ (.Y(_13666_),
    .A(_01922_),
    .B(_13664_));
 sg13g2_and3_1 _27279_ (.X(_13667_),
    .A(_01923_),
    .B(_01922_),
    .C(_13664_));
 sg13g2_nand2_1 _27280_ (.Y(_13668_),
    .A(_01924_),
    .B(_13667_));
 sg13g2_nand3_1 _27281_ (.B(_01924_),
    .C(_13667_),
    .A(_01925_),
    .Y(_13669_));
 sg13g2_nor2_1 _27282_ (.A(_08227_),
    .B(_13669_),
    .Y(_13670_));
 sg13g2_and2_1 _27283_ (.A(_01927_),
    .B(_13670_),
    .X(_13671_));
 sg13g2_nand2_1 _27284_ (.Y(_13672_),
    .A(_01929_),
    .B(_13671_));
 sg13g2_and3_1 _27285_ (.X(_13673_),
    .A(_01930_),
    .B(_01929_),
    .C(_13671_));
 sg13g2_and2_1 _27286_ (.A(_01931_),
    .B(_13673_),
    .X(_13674_));
 sg13g2_nand2_1 _27287_ (.Y(_13675_),
    .A(_01932_),
    .B(_13674_));
 sg13g2_and3_1 _27288_ (.X(_13676_),
    .A(_01933_),
    .B(_01932_),
    .C(_13674_));
 sg13g2_and2_1 _27289_ (.A(_01934_),
    .B(_13676_),
    .X(_13677_));
 sg13g2_nand2_1 _27290_ (.Y(_13678_),
    .A(_01935_),
    .B(_13677_));
 sg13g2_and3_1 _27291_ (.X(_13679_),
    .A(_01936_),
    .B(_01935_),
    .C(_13677_));
 sg13g2_and2_1 _27292_ (.A(_01937_),
    .B(_13679_),
    .X(_13680_));
 sg13g2_or2_1 _27293_ (.X(_13681_),
    .B(_13665_),
    .A(net7588));
 sg13g2_nand2_1 _27294_ (.Y(_13682_),
    .A(_01938_),
    .B(_13680_));
 sg13g2_nand3_1 _27295_ (.B(_01938_),
    .C(_13680_),
    .A(_01940_),
    .Y(_13683_));
 sg13g2_xor2_1 _27296_ (.B(_13683_),
    .A(_01941_),
    .X(_13684_));
 sg13g2_o21ai_1 _27297_ (.B1(_13661_),
    .Y(_13685_),
    .A1(net7622),
    .A2(_13684_));
 sg13g2_nand2b_1 _27298_ (.Y(_13686_),
    .B(_13441_),
    .A_N(_13574_));
 sg13g2_a22oi_1 _27299_ (.Y(_13687_),
    .B1(_13686_),
    .B2(net6653),
    .A2(_13685_),
    .A1(net6644));
 sg13g2_a21oi_1 _27300_ (.A1(_05314_),
    .A2(net6536),
    .Y(_13688_),
    .B1(_13687_));
 sg13g2_a22oi_1 _27301_ (.Y(_13689_),
    .B1(net7350),
    .B2(net7678),
    .A2(net6987),
    .A1(_01972_));
 sg13g2_xor2_1 _27302_ (.B(_13682_),
    .A(_01940_),
    .X(_13690_));
 sg13g2_o21ai_1 _27303_ (.B1(_13689_),
    .Y(_13691_),
    .A1(net7622),
    .A2(_13690_));
 sg13g2_nand2b_1 _27304_ (.Y(_13692_),
    .B(_13446_),
    .A_N(net6541));
 sg13g2_a22oi_1 _27305_ (.Y(_13693_),
    .B1(_13692_),
    .B2(net6655),
    .A2(_13691_),
    .A1(net6643));
 sg13g2_a21oi_1 _27306_ (.A1(_05317_),
    .A2(_13576_),
    .Y(_13694_),
    .B1(_13693_));
 sg13g2_mux2_1 _27307_ (.A0(_01561_),
    .A1(_01596_),
    .S(net7802),
    .X(_13695_));
 sg13g2_a21o_1 _27308_ (.A2(\id_stage_i.controller_i.instr_fetch_err_plus2_i ),
    .A1(_01928_),
    .B1(_01939_),
    .X(_13696_));
 sg13g2_and3_1 _27309_ (.X(_13697_),
    .A(_06901_),
    .B(_13583_),
    .C(_13696_));
 sg13g2_mux2_1 _27310_ (.A0(_01908_),
    .A1(_01878_),
    .S(\id_stage_i.controller_i.instr_is_compressed_i ),
    .X(_13698_));
 sg13g2_nor2_1 _27311_ (.A(net7555),
    .B(_13695_),
    .Y(_13699_));
 sg13g2_a221oi_1 _27312_ (.B2(_13698_),
    .C1(_13697_),
    .B1(net7420),
    .A1(_01971_),
    .Y(_13700_),
    .A2(net6985));
 sg13g2_nand2b_1 _27313_ (.Y(_13701_),
    .B(_13578_),
    .A_N(_13700_));
 sg13g2_nor3_1 _27314_ (.A(net7028),
    .B(net7416),
    .C(_09956_),
    .Y(_13702_));
 sg13g2_a21o_1 _27315_ (.A2(net7312),
    .A1(net7028),
    .B1(_13702_),
    .X(_13703_));
 sg13g2_inv_1 _27316_ (.Y(_13704_),
    .A(_13703_));
 sg13g2_o21ai_1 _27317_ (.B1(net6656),
    .Y(_13705_),
    .A1(_13574_),
    .A2(_13703_));
 sg13g2_a22oi_1 _27318_ (.Y(_13706_),
    .B1(_13701_),
    .B2(_13705_),
    .A2(net6536),
    .A1(_05323_));
 sg13g2_a22oi_1 _27319_ (.Y(_13707_),
    .B1(net7350),
    .B2(net7680),
    .A2(net6987),
    .A1(_01970_));
 sg13g2_xnor2_1 _27320_ (.Y(_13708_),
    .A(_01938_),
    .B(_13680_));
 sg13g2_o21ai_1 _27321_ (.B1(_13707_),
    .Y(_13709_),
    .A1(net7624),
    .A2(_13708_));
 sg13g2_nand2b_1 _27322_ (.Y(_13710_),
    .B(net6155),
    .A_N(net6538));
 sg13g2_a22oi_1 _27323_ (.Y(_13711_),
    .B1(_13710_),
    .B2(net6655),
    .A2(_13709_),
    .A1(net6643));
 sg13g2_a21oi_1 _27324_ (.A1(_05326_),
    .A2(net6535),
    .Y(_13712_),
    .B1(_13711_));
 sg13g2_a22oi_1 _27325_ (.Y(_13713_),
    .B1(net7350),
    .B2(net7681),
    .A2(net6987),
    .A1(_01969_));
 sg13g2_xnor2_1 _27326_ (.Y(_13714_),
    .A(_01937_),
    .B(_13679_));
 sg13g2_mux2_1 _27327_ (.A0(_01491_),
    .A1(_01526_),
    .S(net7791),
    .X(_13715_));
 sg13g2_o21ai_1 _27328_ (.B1(_13713_),
    .Y(_13716_),
    .A1(net7624),
    .A2(_13714_));
 sg13g2_nand2b_1 _27329_ (.Y(_13717_),
    .B(_13458_),
    .A_N(net6538));
 sg13g2_a22oi_1 _27330_ (.Y(_13718_),
    .B1(_13717_),
    .B2(net6655),
    .A2(_13716_),
    .A1(net6643));
 sg13g2_a21oi_1 _27331_ (.A1(_05331_),
    .A2(net6535),
    .Y(_13719_),
    .B1(_13718_));
 sg13g2_nor3_1 _27332_ (.A(net7573),
    .B(net7562),
    .C(_13715_),
    .Y(_13720_));
 sg13g2_a22oi_1 _27333_ (.Y(_13721_),
    .B1(net7351),
    .B2(net7682),
    .A2(net6986),
    .A1(_01968_));
 sg13g2_xor2_1 _27334_ (.B(_13678_),
    .A(_01936_),
    .X(_13722_));
 sg13g2_o21ai_1 _27335_ (.B1(_13721_),
    .Y(_13723_),
    .A1(net7623),
    .A2(_13722_));
 sg13g2_nand2b_1 _27336_ (.Y(_13724_),
    .B(net6152),
    .A_N(net6537));
 sg13g2_a22oi_1 _27337_ (.Y(_13725_),
    .B1(_13724_),
    .B2(net6654),
    .A2(_13723_),
    .A1(net6642));
 sg13g2_a21oi_1 _27338_ (.A1(_05334_),
    .A2(net6534),
    .Y(_13726_),
    .B1(_13725_));
 sg13g2_a22oi_1 _27339_ (.Y(_13727_),
    .B1(net7351),
    .B2(net7683),
    .A2(net6986),
    .A1(_01967_));
 sg13g2_xnor2_1 _27340_ (.Y(_13728_),
    .A(_01935_),
    .B(_13677_));
 sg13g2_o21ai_1 _27341_ (.B1(_13727_),
    .Y(_13729_),
    .A1(net7623),
    .A2(_13728_));
 sg13g2_nand2b_1 _27342_ (.Y(_13730_),
    .B(_13471_),
    .A_N(net6537));
 sg13g2_a22oi_1 _27343_ (.Y(_13731_),
    .B1(_13730_),
    .B2(net6654),
    .A2(_13729_),
    .A1(net6642));
 sg13g2_a21oi_1 _27344_ (.A1(_05339_),
    .A2(net6534),
    .Y(_13732_),
    .B1(_13731_));
 sg13g2_a22oi_1 _27345_ (.Y(_13733_),
    .B1(net7351),
    .B2(net7684),
    .A2(net6986),
    .A1(_01966_));
 sg13g2_xnor2_1 _27346_ (.Y(_13734_),
    .A(_01934_),
    .B(_13676_));
 sg13g2_o21ai_1 _27347_ (.B1(_13733_),
    .Y(_13735_),
    .A1(net7623),
    .A2(_13734_));
 sg13g2_nand2b_1 _27348_ (.Y(_13736_),
    .B(_13477_),
    .A_N(net6537));
 sg13g2_a22oi_1 _27349_ (.Y(_13737_),
    .B1(_13736_),
    .B2(net6654),
    .A2(_13735_),
    .A1(net6642));
 sg13g2_a21oi_1 _27350_ (.A1(_05343_),
    .A2(net6535),
    .Y(_13738_),
    .B1(_13737_));
 sg13g2_a22oi_1 _27351_ (.Y(_13739_),
    .B1(net7351),
    .B2(net7685),
    .A2(net6986),
    .A1(_01965_));
 sg13g2_mux2_1 _27352_ (.A0(_01350_),
    .A1(_01385_),
    .S(net7792),
    .X(_13740_));
 sg13g2_xor2_1 _27353_ (.B(_13675_),
    .A(_01933_),
    .X(_13741_));
 sg13g2_o21ai_1 _27354_ (.B1(_13739_),
    .Y(_13742_),
    .A1(net7623),
    .A2(_13741_));
 sg13g2_nand2b_1 _27355_ (.Y(_13743_),
    .B(net6148),
    .A_N(net6537));
 sg13g2_nor3_1 _27356_ (.A(net7573),
    .B(net7558),
    .C(_13740_),
    .Y(_13744_));
 sg13g2_a22oi_1 _27357_ (.Y(_13745_),
    .B1(_13743_),
    .B2(net6654),
    .A2(_13742_),
    .A1(net6642));
 sg13g2_a21oi_1 _27358_ (.A1(_05348_),
    .A2(net6534),
    .Y(_13746_),
    .B1(_13745_));
 sg13g2_a22oi_1 _27359_ (.Y(_13747_),
    .B1(net7351),
    .B2(net7692),
    .A2(net6986),
    .A1(_01964_));
 sg13g2_xnor2_1 _27360_ (.Y(_13748_),
    .A(_01932_),
    .B(_13674_));
 sg13g2_o21ai_1 _27361_ (.B1(_13747_),
    .Y(_13749_),
    .A1(net7623),
    .A2(_13748_));
 sg13g2_nand2b_1 _27362_ (.Y(_13750_),
    .B(net6146),
    .A_N(net6537));
 sg13g2_a22oi_1 _27363_ (.Y(_13751_),
    .B1(_13750_),
    .B2(net6654),
    .A2(_13749_),
    .A1(net6642));
 sg13g2_a21oi_1 _27364_ (.A1(_05350_),
    .A2(net6535),
    .Y(_13752_),
    .B1(_13751_));
 sg13g2_a22oi_1 _27365_ (.Y(_13753_),
    .B1(net7351),
    .B2(net7699),
    .A2(net6986),
    .A1(_01963_));
 sg13g2_xnor2_1 _27366_ (.Y(_13754_),
    .A(_01931_),
    .B(_13673_));
 sg13g2_o21ai_1 _27367_ (.B1(_13753_),
    .Y(_13755_),
    .A1(net7623),
    .A2(_13754_));
 sg13g2_nand2b_1 _27368_ (.Y(_13756_),
    .B(_13495_),
    .A_N(net6537));
 sg13g2_a22oi_1 _27369_ (.Y(_13757_),
    .B1(_13756_),
    .B2(net6654),
    .A2(_13755_),
    .A1(net6642));
 sg13g2_a21oi_1 _27370_ (.A1(_05354_),
    .A2(net6534),
    .Y(_13758_),
    .B1(_13757_));
 sg13g2_a22oi_1 _27371_ (.Y(_13759_),
    .B1(net7351),
    .B2(net7734),
    .A2(net6986),
    .A1(_01962_));
 sg13g2_xor2_1 _27372_ (.B(_13672_),
    .A(_01930_),
    .X(_13760_));
 sg13g2_o21ai_1 _27373_ (.B1(_13759_),
    .Y(_13761_),
    .A1(net7623),
    .A2(_13760_));
 sg13g2_nand2b_1 _27374_ (.Y(_13762_),
    .B(_13501_),
    .A_N(_13574_));
 sg13g2_mux2_1 _27375_ (.A0(_01420_),
    .A1(_01455_),
    .S(net7791),
    .X(_13763_));
 sg13g2_a22oi_1 _27376_ (.Y(_13764_),
    .B1(_13762_),
    .B2(net6653),
    .A2(_13761_),
    .A1(net6644));
 sg13g2_a21oi_1 _27377_ (.A1(_05358_),
    .A2(_13576_),
    .Y(_13765_),
    .B1(_13764_));
 sg13g2_nor3_1 _27378_ (.A(net7574),
    .B(net7571),
    .C(_13763_),
    .Y(_13766_));
 sg13g2_xnor2_1 _27379_ (.Y(_13767_),
    .A(_01929_),
    .B(_13671_));
 sg13g2_a22oi_1 _27380_ (.Y(_13768_),
    .B1(net7351),
    .B2(net7748),
    .A2(net6986),
    .A1(_01961_));
 sg13g2_o21ai_1 _27381_ (.B1(_13768_),
    .Y(_13769_),
    .A1(net7624),
    .A2(_13767_));
 sg13g2_nand2b_1 _27382_ (.Y(_13770_),
    .B(net6142),
    .A_N(net6537));
 sg13g2_a22oi_1 _27383_ (.Y(_13771_),
    .B1(_13770_),
    .B2(net6654),
    .A2(_13769_),
    .A1(net6642));
 sg13g2_a21oi_1 _27384_ (.A1(_05364_),
    .A2(net6534),
    .Y(_13772_),
    .B1(_13771_));
 sg13g2_mux2_1 _27385_ (.A0(_01897_),
    .A1(_01877_),
    .S(\id_stage_i.controller_i.instr_is_compressed_i ),
    .X(_13773_));
 sg13g2_xnor2_1 _27386_ (.Y(_13774_),
    .A(_01928_),
    .B(\id_stage_i.controller_i.instr_fetch_err_plus2_i ));
 sg13g2_nor2_1 _27387_ (.A(net7625),
    .B(_13774_),
    .Y(_13775_));
 sg13g2_a221oi_1 _27388_ (.B2(_13773_),
    .C1(_13775_),
    .B1(net7420),
    .A1(_01960_),
    .Y(_13776_),
    .A2(net6985));
 sg13g2_nand2b_1 _27389_ (.Y(_13777_),
    .B(_13578_),
    .A_N(_13776_));
 sg13g2_nand3b_1 _27390_ (.B(_06967_),
    .C(net7029),
    .Y(_13778_),
    .A_N(_10007_));
 sg13g2_inv_1 _27391_ (.Y(_13779_),
    .A(_13780_));
 sg13g2_o21ai_1 _27392_ (.B1(_13778_),
    .Y(_13780_),
    .A1(net7029),
    .A2(_06969_));
 sg13g2_o21ai_1 _27393_ (.B1(net6657),
    .Y(_13781_),
    .A1(net6539),
    .A2(_13780_));
 sg13g2_a22oi_1 _27394_ (.Y(_13782_),
    .B1(_13777_),
    .B2(_13781_),
    .A2(net6536),
    .A1(_05371_));
 sg13g2_nor4_1 _27395_ (.A(_13699_),
    .B(_13720_),
    .C(_13744_),
    .D(_13766_),
    .Y(_13783_));
 sg13g2_xnor2_1 _27396_ (.Y(_13784_),
    .A(_01927_),
    .B(_13670_));
 sg13g2_a22oi_1 _27397_ (.Y(_13785_),
    .B1(net7350),
    .B2(net7805),
    .A2(net6987),
    .A1(_01959_));
 sg13g2_o21ai_1 _27398_ (.B1(_13785_),
    .Y(_13786_),
    .A1(net7624),
    .A2(_13784_));
 sg13g2_nand2b_1 _27399_ (.Y(_13787_),
    .B(_13511_),
    .A_N(net6537));
 sg13g2_a22oi_1 _27400_ (.Y(_13788_),
    .B1(_13787_),
    .B2(net6654),
    .A2(_13786_),
    .A1(net6642));
 sg13g2_a21oi_1 _27401_ (.A1(_05382_),
    .A2(net6534),
    .Y(_13789_),
    .B1(_13788_));
 sg13g2_a22oi_1 _27402_ (.Y(_13790_),
    .B1(net7350),
    .B2(net7807),
    .A2(net6987),
    .A1(_01958_));
 sg13g2_xnor2_1 _27403_ (.Y(_13791_),
    .A(_08227_),
    .B(_13669_));
 sg13g2_o21ai_1 _27404_ (.B1(_13790_),
    .Y(_13792_),
    .A1(net7622),
    .A2(_13791_));
 sg13g2_nand2b_1 _27405_ (.Y(_13793_),
    .B(net6140),
    .A_N(net6538));
 sg13g2_a22oi_1 _27406_ (.Y(_13794_),
    .B1(_13793_),
    .B2(net6655),
    .A2(_13792_),
    .A1(net6643));
 sg13g2_a21oi_1 _27407_ (.A1(_05388_),
    .A2(net6535),
    .Y(_13795_),
    .B1(_13794_));
 sg13g2_a22oi_1 _27408_ (.Y(_13796_),
    .B1(net7350),
    .B2(net7810),
    .A2(net6988),
    .A1(_01957_));
 sg13g2_xor2_1 _27409_ (.B(_13668_),
    .A(_01925_),
    .X(_13797_));
 sg13g2_o21ai_1 _27410_ (.B1(_13796_),
    .Y(_13798_),
    .A1(net7622),
    .A2(_13797_));
 sg13g2_nand2_1 _27411_ (.Y(_13799_),
    .A(net6643),
    .B(_13798_));
 sg13g2_nor2_1 _27412_ (.A(_13522_),
    .B(net6538),
    .Y(_13800_));
 sg13g2_a21oi_1 _27413_ (.A1(_00483_),
    .A2(net6538),
    .Y(_13801_),
    .B1(_13800_));
 sg13g2_o21ai_1 _27414_ (.B1(_13799_),
    .Y(_13802_),
    .A1(net6668),
    .A2(_13801_));
 sg13g2_nand4_1 _27415_ (.B(_13629_),
    .C(_13681_),
    .A(_13580_),
    .Y(_13803_),
    .D(_13783_));
 sg13g2_a22oi_1 _27416_ (.Y(_13804_),
    .B1(net7350),
    .B2(net7820),
    .A2(net6987),
    .A1(_01956_));
 sg13g2_nor2_1 _27417_ (.A(net7291),
    .B(net7074),
    .Y(_13805_));
 sg13g2_xnor2_1 _27418_ (.Y(_13806_),
    .A(_01924_),
    .B(_13667_));
 sg13g2_o21ai_1 _27419_ (.B1(_13804_),
    .Y(_13807_),
    .A1(net7622),
    .A2(_13806_));
 sg13g2_nand2_1 _27420_ (.Y(_13808_),
    .A(net6641),
    .B(_13807_));
 sg13g2_nor2_1 _27421_ (.A(_13527_),
    .B(net6540),
    .Y(_13809_));
 sg13g2_a21oi_1 _27422_ (.A1(_00482_),
    .A2(net6540),
    .Y(_13810_),
    .B1(_13809_));
 sg13g2_o21ai_1 _27423_ (.B1(_13808_),
    .Y(_13811_),
    .A1(net6658),
    .A2(_13810_));
 sg13g2_mux2_1 _27424_ (.A0(net7838),
    .A1(_01876_),
    .S(net7935),
    .X(_13812_));
 sg13g2_a22oi_1 _27425_ (.Y(_13813_),
    .B1(net7419),
    .B2(_13812_),
    .A2(_07762_),
    .A1(_01955_));
 sg13g2_xor2_1 _27426_ (.B(_13666_),
    .A(_01923_),
    .X(_13814_));
 sg13g2_o21ai_1 _27427_ (.B1(_13813_),
    .Y(_13815_),
    .A1(net7622),
    .A2(_13814_));
 sg13g2_nand2_1 _27428_ (.Y(_13816_),
    .A(_13578_),
    .B(_13815_));
 sg13g2_nor2_1 _27429_ (.A(_13532_),
    .B(net6539),
    .Y(_13817_));
 sg13g2_a21oi_1 _27430_ (.A1(_00481_),
    .A2(net6539),
    .Y(_13818_),
    .B1(_13817_));
 sg13g2_o21ai_1 _27431_ (.B1(_13816_),
    .Y(_13819_),
    .A1(_13572_),
    .A2(_13818_));
 sg13g2_nand2_1 _27432_ (.Y(_13820_),
    .A(_01875_),
    .B(net7936));
 sg13g2_o21ai_1 _27433_ (.B1(_13820_),
    .Y(_13821_),
    .A1(_09244_),
    .A2(net7935));
 sg13g2_a22oi_1 _27434_ (.Y(_13822_),
    .B1(net7419),
    .B2(_13821_),
    .A2(_07762_),
    .A1(_01954_));
 sg13g2_xnor2_1 _27435_ (.Y(_13823_),
    .A(_01922_),
    .B(_13664_));
 sg13g2_o21ai_1 _27436_ (.B1(_13822_),
    .Y(_13824_),
    .A1(net7625),
    .A2(_13823_));
 sg13g2_nand2_1 _27437_ (.Y(_13825_),
    .A(_13578_),
    .B(_13824_));
 sg13g2_nor2_1 _27438_ (.A(net6542),
    .B(net6541),
    .Y(_13826_));
 sg13g2_a21oi_1 _27439_ (.A1(_00480_),
    .A2(net6541),
    .Y(_13827_),
    .B1(_13826_));
 sg13g2_o21ai_1 _27440_ (.B1(_13825_),
    .Y(_13828_),
    .A1(net6662),
    .A2(_13827_));
 sg13g2_nand2_1 _27441_ (.Y(_13829_),
    .A(_01874_),
    .B(net7934));
 sg13g2_o21ai_1 _27442_ (.B1(_13829_),
    .Y(_13830_),
    .A1(_09282_),
    .A2(net7935));
 sg13g2_a22oi_1 _27443_ (.Y(_13831_),
    .B1(net7419),
    .B2(_13830_),
    .A2(net6985),
    .A1(_01953_));
 sg13g2_nand2_1 _27444_ (.Y(_13832_),
    .A(_01919_),
    .B(_13663_));
 sg13g2_nand3_1 _27445_ (.B(_01919_),
    .C(_13663_),
    .A(_01920_),
    .Y(_13833_));
 sg13g2_xor2_1 _27446_ (.B(_13833_),
    .A(_01921_),
    .X(_13834_));
 sg13g2_o21ai_1 _27447_ (.B1(_13831_),
    .Y(_13835_),
    .A1(net7625),
    .A2(_13834_));
 sg13g2_nand2_1 _27448_ (.Y(_13836_),
    .A(net6641),
    .B(_13835_));
 sg13g2_nor2_1 _27449_ (.A(net6136),
    .B(net6541),
    .Y(_13837_));
 sg13g2_a21o_1 _27450_ (.A2(net7039),
    .A1(net7684),
    .B1(_13805_),
    .X(_13838_));
 sg13g2_a21oi_1 _27451_ (.A1(_00479_),
    .A2(net6541),
    .Y(_13839_),
    .B1(_13837_));
 sg13g2_a21oi_1 _27452_ (.A1(net7684),
    .A2(net7039),
    .Y(_13840_),
    .B1(_13805_));
 sg13g2_o21ai_1 _27453_ (.B1(_13836_),
    .Y(_13841_),
    .A1(net6662),
    .A2(_13839_));
 sg13g2_nand2_1 _27454_ (.Y(_13842_),
    .A(_01873_),
    .B(net7934));
 sg13g2_o21ai_1 _27455_ (.B1(_13842_),
    .Y(_13843_),
    .A1(_09324_),
    .A2(net7935));
 sg13g2_a22oi_1 _27456_ (.Y(_13844_),
    .B1(net7419),
    .B2(_13843_),
    .A2(_07762_),
    .A1(_01952_));
 sg13g2_xor2_1 _27457_ (.B(_13832_),
    .A(_01920_),
    .X(_13845_));
 sg13g2_o21ai_1 _27458_ (.B1(_13844_),
    .Y(_13846_),
    .A1(net7625),
    .A2(_13845_));
 sg13g2_nand2_1 _27459_ (.Y(_13847_),
    .A(net6641),
    .B(_13846_));
 sg13g2_nor2_1 _27460_ (.A(_13547_),
    .B(net6540),
    .Y(_13848_));
 sg13g2_a21oi_1 _27461_ (.A1(_00478_),
    .A2(net6540),
    .Y(_13849_),
    .B1(_13848_));
 sg13g2_o21ai_1 _27462_ (.B1(_13847_),
    .Y(_13850_),
    .A1(net6658),
    .A2(_13849_));
 sg13g2_nand2_1 _27463_ (.Y(_13851_),
    .A(_01872_),
    .B(net7933));
 sg13g2_o21ai_1 _27464_ (.B1(_13851_),
    .Y(_13852_),
    .A1(_09373_),
    .A2(net7933));
 sg13g2_a22oi_1 _27465_ (.Y(_13853_),
    .B1(net7419),
    .B2(_13852_),
    .A2(net6985),
    .A1(_01951_));
 sg13g2_xnor2_1 _27466_ (.Y(_13854_),
    .A(_01919_),
    .B(_13663_));
 sg13g2_o21ai_1 _27467_ (.B1(_13853_),
    .Y(_13855_),
    .A1(net7625),
    .A2(_13854_));
 sg13g2_nand2_1 _27468_ (.Y(_13856_),
    .A(net6641),
    .B(_13855_));
 sg13g2_nor2_1 _27469_ (.A(net6134),
    .B(net6538),
    .Y(_13857_));
 sg13g2_a21oi_1 _27470_ (.A1(_00477_),
    .A2(net6538),
    .Y(_13858_),
    .B1(_13857_));
 sg13g2_o21ai_1 _27471_ (.B1(_13856_),
    .Y(_13859_),
    .A1(net6668),
    .A2(_13858_));
 sg13g2_mux2_1 _27472_ (.A0(net7932),
    .A1(_01871_),
    .S(\id_stage_i.controller_i.instr_is_compressed_i ),
    .X(_13860_));
 sg13g2_a22oi_1 _27473_ (.Y(_13861_),
    .B1(net7419),
    .B2(_13860_),
    .A2(net6985),
    .A1(_01950_));
 sg13g2_xnor2_1 _27474_ (.Y(_13862_),
    .A(_08414_),
    .B(_13662_));
 sg13g2_o21ai_1 _27475_ (.B1(_13861_),
    .Y(_13863_),
    .A1(net7625),
    .A2(_13862_));
 sg13g2_nand2_1 _27476_ (.Y(_13864_),
    .A(net6641),
    .B(_13863_));
 sg13g2_nor2_1 _27477_ (.A(net6455),
    .B(net6541),
    .Y(_13865_));
 sg13g2_a21oi_1 _27478_ (.A1(_00476_),
    .A2(net6541),
    .Y(_13866_),
    .B1(_13865_));
 sg13g2_o21ai_1 _27479_ (.B1(_13864_),
    .Y(_13867_),
    .A1(net6662),
    .A2(_13866_));
 sg13g2_mux2_1 _27480_ (.A0(_01886_),
    .A1(_01870_),
    .S(net7936),
    .X(_13868_));
 sg13g2_a22oi_1 _27481_ (.Y(_13869_),
    .B1(net7420),
    .B2(_13868_),
    .A2(net6985),
    .A1(_01949_));
 sg13g2_nand2b_1 _27482_ (.Y(_13870_),
    .B(_13578_),
    .A_N(_13869_));
 sg13g2_nor2_1 _27483_ (.A(_06968_),
    .B(_10076_),
    .Y(_13871_));
 sg13g2_nor2_1 _27484_ (.A(net7072),
    .B(_13871_),
    .Y(_13872_));
 sg13g2_a21oi_1 _27485_ (.A1(net7072),
    .A2(_06969_),
    .Y(_13873_),
    .B1(_13872_));
 sg13g2_inv_1 _27486_ (.Y(_13874_),
    .A(_13873_));
 sg13g2_mux2_1 _27487_ (.A0(_01269_),
    .A1(_00629_),
    .S(net7885),
    .X(_13875_));
 sg13g2_nand2b_1 _27488_ (.Y(_13876_),
    .B(_13575_),
    .A_N(_00475_));
 sg13g2_o21ai_1 _27489_ (.B1(_13876_),
    .Y(_13877_),
    .A1(_13575_),
    .A2(_13873_));
 sg13g2_o21ai_1 _27490_ (.B1(_13870_),
    .Y(_13878_),
    .A1(_13572_),
    .A2(_13877_));
 sg13g2_a21oi_1 _27491_ (.A1(_09320_),
    .A2(net6728),
    .Y(_13879_),
    .B1(net6668));
 sg13g2_nand2_1 _27492_ (.Y(_13880_),
    .A(_09547_),
    .B(net6592));
 sg13g2_nand2_1 _27493_ (.Y(_13881_),
    .A(\cs_registers_i.csr_mstatus_mie_o ),
    .B(net6532));
 sg13g2_o21ai_1 _27494_ (.B1(_13881_),
    .Y(_13882_),
    .A1(_13656_),
    .A2(net6532));
 sg13g2_nand2_1 _27495_ (.Y(_13883_),
    .A(_13879_),
    .B(_13882_));
 sg13g2_o21ai_1 _27496_ (.B1(_13883_),
    .Y(_13884_),
    .A1(_00003_),
    .A2(net7078));
 sg13g2_nand2_1 _27497_ (.Y(_13885_),
    .A(net7982),
    .B(_00002_));
 sg13g2_a21oi_1 _27498_ (.A1(net7079),
    .A2(_13885_),
    .Y(_13886_),
    .B1(\cs_registers_i.csr_mstatus_mie_o ));
 sg13g2_nand2_1 _27499_ (.Y(_13887_),
    .A(_00003_),
    .B(net6532));
 sg13g2_o21ai_1 _27500_ (.B1(net6653),
    .Y(_13888_),
    .A1(net7079),
    .A2(_13887_));
 sg13g2_o21ai_1 _27501_ (.B1(_13888_),
    .Y(_13889_),
    .A1(net6653),
    .A2(_13886_));
 sg13g2_nand2b_1 _27502_ (.Y(_13890_),
    .B(net6132),
    .A_N(net6532));
 sg13g2_nand3_1 _27503_ (.B(_13887_),
    .C(_13890_),
    .A(_13879_),
    .Y(_13891_));
 sg13g2_o21ai_1 _27504_ (.B1(net6532),
    .Y(_13892_),
    .A1(net7078),
    .A2(_13885_));
 sg13g2_nand3_1 _27505_ (.B(_13891_),
    .C(_13892_),
    .A(net6653),
    .Y(_13893_));
 sg13g2_nand2_1 _27506_ (.Y(_13894_),
    .A(_13889_),
    .B(_13893_));
 sg13g2_nor2_1 _27507_ (.A(_02211_),
    .B(_09321_),
    .Y(_13895_));
 sg13g2_a22oi_1 _27508_ (.Y(_13896_),
    .B1(net7036),
    .B2(_00439_),
    .A2(net6658),
    .A1(_06152_));
 sg13g2_nand2_1 _27509_ (.Y(_13897_),
    .A(_13547_),
    .B(_13553_));
 sg13g2_o21ai_1 _27510_ (.B1(_13879_),
    .Y(_13898_),
    .A1(net6532),
    .A2(_13897_));
 sg13g2_a21oi_1 _27511_ (.A1(_09547_),
    .A2(_13423_),
    .Y(_13899_),
    .B1(_00474_));
 sg13g2_o21ai_1 _27512_ (.B1(_13896_),
    .Y(_13900_),
    .A1(_13898_),
    .A2(_13899_));
 sg13g2_a22oi_1 _27513_ (.Y(_13901_),
    .B1(net7036),
    .B2(_00438_),
    .A2(net6658),
    .A1(_06162_));
 sg13g2_a21oi_1 _27514_ (.A1(_09547_),
    .A2(_13423_),
    .Y(_13902_),
    .B1(_00473_));
 sg13g2_o21ai_1 _27515_ (.B1(_13901_),
    .Y(_13903_),
    .A1(_13898_),
    .A2(_13902_));
 sg13g2_nand2_1 _27516_ (.Y(_13904_),
    .A(_00472_),
    .B(_13880_));
 sg13g2_o21ai_1 _27517_ (.B1(_13904_),
    .Y(_13905_),
    .A1(net6138),
    .A2(_13880_));
 sg13g2_nand2_1 _27518_ (.Y(_13906_),
    .A(\cs_registers_i.csr_mstatus_tw_o ),
    .B(net6532));
 sg13g2_a22oi_1 _27519_ (.Y(_13907_),
    .B1(_13875_),
    .B2(net7824),
    .A2(net7527),
    .A1(_00917_));
 sg13g2_o21ai_1 _27520_ (.B1(_13906_),
    .Y(_13908_),
    .A1(net6143),
    .A2(net6532));
 sg13g2_mux2_1 _27521_ (.A0(_00471_),
    .A1(_00381_),
    .S(net6660),
    .X(_13909_));
 sg13g2_mux2_1 _27522_ (.A0(_00470_),
    .A1(_00380_),
    .S(net6669),
    .X(_13910_));
 sg13g2_mux2_1 _27523_ (.A0(_00469_),
    .A1(_00379_),
    .S(net6661),
    .X(_13911_));
 sg13g2_mux2_1 _27524_ (.A0(_00468_),
    .A1(_00378_),
    .S(net6659),
    .X(_13912_));
 sg13g2_mux2_1 _27525_ (.A0(_00467_),
    .A1(_00377_),
    .S(net6659),
    .X(_13913_));
 sg13g2_nand2_1 _27526_ (.Y(_13914_),
    .A(_00466_),
    .B(_13573_));
 sg13g2_o21ai_1 _27527_ (.B1(_13914_),
    .Y(_13915_),
    .A1(_05742_),
    .A2(_13573_));
 sg13g2_nand2_1 _27528_ (.Y(_13916_),
    .A(_00465_),
    .B(_13573_));
 sg13g2_o21ai_1 _27529_ (.B1(_13916_),
    .Y(_13917_),
    .A1(_05744_),
    .A2(_13573_));
 sg13g2_mux2_1 _27530_ (.A0(_00464_),
    .A1(_00374_),
    .S(net6660),
    .X(_13918_));
 sg13g2_mux2_1 _27531_ (.A0(_00463_),
    .A1(_00373_),
    .S(net6665),
    .X(_13919_));
 sg13g2_nand2_1 _27532_ (.Y(_13920_),
    .A(_00372_),
    .B(net6659));
 sg13g2_o21ai_1 _27533_ (.B1(_13920_),
    .Y(_13921_),
    .A1(_05464_),
    .A2(net6659));
 sg13g2_mux2_1 _27534_ (.A0(_00461_),
    .A1(_00371_),
    .S(net6665),
    .X(_13922_));
 sg13g2_mux2_1 _27535_ (.A0(_00460_),
    .A1(_00370_),
    .S(net6665),
    .X(_13923_));
 sg13g2_mux2_1 _27536_ (.A0(_00459_),
    .A1(_00369_),
    .S(net6663),
    .X(_13924_));
 sg13g2_mux2_1 _27537_ (.A0(_00458_),
    .A1(_00368_),
    .S(net6664),
    .X(_13925_));
 sg13g2_nand2b_1 _27538_ (.Y(_13926_),
    .B(net7885),
    .A_N(_00697_));
 sg13g2_mux2_1 _27539_ (.A0(_00457_),
    .A1(_00367_),
    .S(net6664),
    .X(_13927_));
 sg13g2_mux2_1 _27540_ (.A0(_00456_),
    .A1(_00366_),
    .S(net6664),
    .X(_13928_));
 sg13g2_mux2_1 _27541_ (.A0(_00455_),
    .A1(_00365_),
    .S(net6663),
    .X(_13929_));
 sg13g2_mux2_1 _27542_ (.A0(_00454_),
    .A1(_00364_),
    .S(net6663),
    .X(_13930_));
 sg13g2_mux2_1 _27543_ (.A0(_00453_),
    .A1(_00363_),
    .S(net6663),
    .X(_13931_));
 sg13g2_mux2_1 _27544_ (.A0(_00452_),
    .A1(_00362_),
    .S(net6663),
    .X(_13932_));
 sg13g2_mux2_1 _27545_ (.A0(_00451_),
    .A1(_00361_),
    .S(_13572_),
    .X(_13933_));
 sg13g2_o21ai_1 _27546_ (.B1(_13926_),
    .Y(_13934_),
    .A1(net7885),
    .A2(_00665_));
 sg13g2_mux2_1 _27547_ (.A0(_00450_),
    .A1(_00360_),
    .S(net6666),
    .X(_13935_));
 sg13g2_mux2_1 _27548_ (.A0(_00449_),
    .A1(_00359_),
    .S(net6665),
    .X(_13936_));
 sg13g2_mux2_1 _27549_ (.A0(_00448_),
    .A1(_00358_),
    .S(net6665),
    .X(_13937_));
 sg13g2_mux2_1 _27550_ (.A0(_00447_),
    .A1(_00357_),
    .S(net6661),
    .X(_13938_));
 sg13g2_mux2_1 _27551_ (.A0(_00446_),
    .A1(_00356_),
    .S(net6659),
    .X(_13939_));
 sg13g2_mux2_1 _27552_ (.A0(_00445_),
    .A1(_00355_),
    .S(net6669),
    .X(_13940_));
 sg13g2_mux2_1 _27553_ (.A0(_00444_),
    .A1(_00354_),
    .S(net6669),
    .X(_13941_));
 sg13g2_mux2_1 _27554_ (.A0(_00443_),
    .A1(_00353_),
    .S(net6669),
    .X(_13942_));
 sg13g2_mux2_1 _27555_ (.A0(_00442_),
    .A1(_00352_),
    .S(net6660),
    .X(_13943_));
 sg13g2_mux2_1 _27556_ (.A0(_00441_),
    .A1(_00351_),
    .S(net6669),
    .X(_13944_));
 sg13g2_mux2_1 _27557_ (.A0(_00440_),
    .A1(_00350_),
    .S(net6658),
    .X(_13945_));
 sg13g2_nand2_1 _27558_ (.Y(_13946_),
    .A(_00002_),
    .B(net6655));
 sg13g2_o21ai_1 _27559_ (.B1(_13946_),
    .Y(_13947_),
    .A1(_05419_),
    .A2(net6655));
 sg13g2_mux2_1 _27560_ (.A0(_00474_),
    .A1(_00439_),
    .S(net6657),
    .X(_13948_));
 sg13g2_mux2_1 _27561_ (.A0(_00473_),
    .A1(_00438_),
    .S(net6656),
    .X(_13949_));
 sg13g2_mux2_1 _27562_ (.A0(_00437_),
    .A1(_00349_),
    .S(net6667),
    .X(_13950_));
 sg13g2_nand2_1 _27563_ (.Y(_13951_),
    .A(_00436_),
    .B(net6657));
 sg13g2_o21ai_1 _27564_ (.B1(_13951_),
    .Y(_13952_),
    .A1(_05827_),
    .A2(net6657));
 sg13g2_nand2_1 _27565_ (.Y(_13953_),
    .A(_00435_),
    .B(net6657));
 sg13g2_o21ai_1 _27566_ (.B1(_13953_),
    .Y(_13954_),
    .A1(_05829_),
    .A2(net6657));
 sg13g2_nand2_1 _27567_ (.Y(_13955_),
    .A(_00346_),
    .B(net6662));
 sg13g2_o21ai_1 _27568_ (.B1(_13955_),
    .Y(_13956_),
    .A1(_05552_),
    .A2(net6662));
 sg13g2_mux2_1 _27569_ (.A0(_00433_),
    .A1(_00345_),
    .S(net6658),
    .X(_13957_));
 sg13g2_mux2_1 _27570_ (.A0(_00432_),
    .A1(_00344_),
    .S(net6662),
    .X(_13958_));
 sg13g2_nand2_1 _27571_ (.Y(_13959_),
    .A(net6678),
    .B(_13420_));
 sg13g2_nand2_1 _27572_ (.Y(_13960_),
    .A(_00431_),
    .B(net6525));
 sg13g2_mux2_1 _27573_ (.A0(_00729_),
    .A1(_00761_),
    .S(net7885),
    .X(_13961_));
 sg13g2_o21ai_1 _27574_ (.B1(_13960_),
    .Y(_13962_),
    .A1(_13431_),
    .A2(net6525));
 sg13g2_nand2_1 _27575_ (.Y(_13963_),
    .A(_00430_),
    .B(_13959_));
 sg13g2_o21ai_1 _27576_ (.B1(_13963_),
    .Y(_13964_),
    .A1(net6159),
    .A2(_13959_));
 sg13g2_nand2_1 _27577_ (.Y(_13965_),
    .A(_00429_),
    .B(net6526));
 sg13g2_o21ai_1 _27578_ (.B1(_13965_),
    .Y(_13966_),
    .A1(net6132),
    .A2(net6526));
 sg13g2_nand2_1 _27579_ (.Y(_13967_),
    .A(_00428_),
    .B(net6524));
 sg13g2_o21ai_1 _27580_ (.B1(_13967_),
    .Y(_13968_),
    .A1(_13621_),
    .A2(net6524));
 sg13g2_nand2_1 _27581_ (.Y(_13969_),
    .A(_00427_),
    .B(_13959_));
 sg13g2_o21ai_1 _27582_ (.B1(_13969_),
    .Y(_13970_),
    .A1(net6533),
    .A2(_13959_));
 sg13g2_nand2_1 _27583_ (.Y(_13971_),
    .A(_00426_),
    .B(net6523));
 sg13g2_o21ai_1 _27584_ (.B1(_13971_),
    .Y(_13972_),
    .A1(_13645_),
    .A2(net6523));
 sg13g2_nand2_1 _27585_ (.Y(_13973_),
    .A(_00425_),
    .B(net6524));
 sg13g2_o21ai_1 _27586_ (.B1(_13973_),
    .Y(_13974_),
    .A1(_13656_),
    .A2(net6524));
 sg13g2_nand2_1 _27587_ (.Y(_13975_),
    .A(_00424_),
    .B(net6525));
 sg13g2_o21ai_1 _27588_ (.B1(net7530),
    .Y(_13976_),
    .A1(net7521),
    .A2(_13961_));
 sg13g2_o21ai_1 _27589_ (.B1(_13975_),
    .Y(_13977_),
    .A1(net6158),
    .A2(net6525));
 sg13g2_a221oi_1 _27590_ (.B2(net7512),
    .C1(_13976_),
    .B1(_13934_),
    .A1(net7483),
    .Y(_13978_),
    .A2(_13907_));
 sg13g2_nand2_1 _27591_ (.Y(_13979_),
    .A(_00423_),
    .B(net6530));
 sg13g2_o21ai_1 _27592_ (.B1(_13979_),
    .Y(_13980_),
    .A1(net6156),
    .A2(net6530));
 sg13g2_nand2_1 _27593_ (.Y(_13981_),
    .A(_00422_),
    .B(net6524));
 sg13g2_o21ai_1 _27594_ (.B1(_13981_),
    .Y(_13982_),
    .A1(_13704_),
    .A2(net6524));
 sg13g2_nand2_1 _27595_ (.Y(_13983_),
    .A(_00421_),
    .B(net6530));
 sg13g2_o21ai_1 _27596_ (.B1(_13983_),
    .Y(_13984_),
    .A1(net6155),
    .A2(net6530));
 sg13g2_nand2_1 _27597_ (.Y(_13985_),
    .A(_00420_),
    .B(net6530));
 sg13g2_o21ai_1 _27598_ (.B1(_13985_),
    .Y(_13986_),
    .A1(net6458),
    .A2(net6530));
 sg13g2_nand2_1 _27599_ (.Y(_13987_),
    .A(_00419_),
    .B(net6529));
 sg13g2_o21ai_1 _27600_ (.B1(_13987_),
    .Y(_13988_),
    .A1(net6152),
    .A2(net6529));
 sg13g2_nand2_1 _27601_ (.Y(_13989_),
    .A(_00418_),
    .B(net6529));
 sg13g2_o21ai_1 _27602_ (.B1(_13989_),
    .Y(_13990_),
    .A1(net6151),
    .A2(net6529));
 sg13g2_nand2_1 _27603_ (.Y(_13991_),
    .A(_00417_),
    .B(net6528));
 sg13g2_mux2_1 _27604_ (.A0(_01279_),
    .A1(_01315_),
    .S(net7887),
    .X(_13992_));
 sg13g2_o21ai_1 _27605_ (.B1(_13991_),
    .Y(_13993_),
    .A1(net6149),
    .A2(net6528));
 sg13g2_nand2_1 _27606_ (.Y(_13994_),
    .A(_00416_),
    .B(net6527));
 sg13g2_nor2_1 _27607_ (.A(net7520),
    .B(_13992_),
    .Y(_13995_));
 sg13g2_o21ai_1 _27608_ (.B1(_13994_),
    .Y(_13996_),
    .A1(net6148),
    .A2(net6527));
 sg13g2_nand2_1 _27609_ (.Y(_13997_),
    .A(_00415_),
    .B(net6527));
 sg13g2_o21ai_1 _27610_ (.B1(_13997_),
    .Y(_13998_),
    .A1(net6146),
    .A2(net6527));
 sg13g2_nand2_1 _27611_ (.Y(_13999_),
    .A(_00414_),
    .B(net6527));
 sg13g2_o21ai_1 _27612_ (.B1(_13999_),
    .Y(_14000_),
    .A1(_13495_),
    .A2(net6527));
 sg13g2_nand2_1 _27613_ (.Y(_14001_),
    .A(_00413_),
    .B(net6527));
 sg13g2_o21ai_1 _27614_ (.B1(_14001_),
    .Y(_14002_),
    .A1(net6143),
    .A2(net6527));
 sg13g2_nand2_1 _27615_ (.Y(_14003_),
    .A(_00412_),
    .B(net6528));
 sg13g2_o21ai_1 _27616_ (.B1(_14003_),
    .Y(_14004_),
    .A1(_13506_),
    .A2(net6528));
 sg13g2_nand2_1 _27617_ (.Y(_14005_),
    .A(_00411_),
    .B(net6523));
 sg13g2_o21ai_1 _27618_ (.B1(_14005_),
    .Y(_14006_),
    .A1(net6454),
    .A2(net6523));
 sg13g2_nand2_1 _27619_ (.Y(_14007_),
    .A(_00410_),
    .B(net6528));
 sg13g2_o21ai_1 _27620_ (.B1(_14007_),
    .Y(_14008_),
    .A1(net6141),
    .A2(net6528));
 sg13g2_nand2_1 _27621_ (.Y(_14009_),
    .A(_00409_),
    .B(net6530));
 sg13g2_mux2_1 _27622_ (.A0(_01068_),
    .A1(_01103_),
    .S(net7887),
    .X(_14010_));
 sg13g2_o21ai_1 _27623_ (.B1(_14009_),
    .Y(_14011_),
    .A1(net6139),
    .A2(net6530));
 sg13g2_nand2_1 _27624_ (.Y(_14012_),
    .A(_00408_),
    .B(net6531));
 sg13g2_nor2_1 _27625_ (.A(net7465),
    .B(_14010_),
    .Y(_14013_));
 sg13g2_o21ai_1 _27626_ (.B1(_14012_),
    .Y(_14014_),
    .A1(net6138),
    .A2(net6531));
 sg13g2_nand2_1 _27627_ (.Y(_14015_),
    .A(_00407_),
    .B(net6528));
 sg13g2_o21ai_1 _27628_ (.B1(_14015_),
    .Y(_14016_),
    .A1(net6137),
    .A2(net6528));
 sg13g2_nand2_1 _27629_ (.Y(_14017_),
    .A(_00406_),
    .B(net6523));
 sg13g2_o21ai_1 _27630_ (.B1(_14017_),
    .Y(_14018_),
    .A1(_13532_),
    .A2(net6523));
 sg13g2_nand2_1 _27631_ (.Y(_14019_),
    .A(_00405_),
    .B(net6529));
 sg13g2_o21ai_1 _27632_ (.B1(_14019_),
    .Y(_14020_),
    .A1(net6542),
    .A2(net6531));
 sg13g2_nand2_1 _27633_ (.Y(_14021_),
    .A(_00404_),
    .B(net6525));
 sg13g2_o21ai_1 _27634_ (.B1(_14021_),
    .Y(_14022_),
    .A1(net6135),
    .A2(net6525));
 sg13g2_nand2_1 _27635_ (.Y(_14023_),
    .A(_00403_),
    .B(_13959_));
 sg13g2_o21ai_1 _27636_ (.B1(_14023_),
    .Y(_14024_),
    .A1(net6457),
    .A2(net6526));
 sg13g2_nand2_1 _27637_ (.Y(_14025_),
    .A(_00402_),
    .B(net6526));
 sg13g2_o21ai_1 _27638_ (.B1(_14025_),
    .Y(_14026_),
    .A1(net6133),
    .A2(net6526));
 sg13g2_nand2_1 _27639_ (.Y(_14027_),
    .A(_00401_),
    .B(net6525));
 sg13g2_mux2_1 _27640_ (.A0(_01139_),
    .A1(_01174_),
    .S(net7887),
    .X(_14028_));
 sg13g2_o21ai_1 _27641_ (.B1(_14027_),
    .Y(_14029_),
    .A1(net6455),
    .A2(net6525));
 sg13g2_nand2_1 _27642_ (.Y(_14030_),
    .A(_00400_),
    .B(net6523));
 sg13g2_nor2_1 _27643_ (.A(net7461),
    .B(_14028_),
    .Y(_14031_));
 sg13g2_o21ai_1 _27644_ (.B1(_14030_),
    .Y(_14032_),
    .A1(_13874_),
    .A2(net6523));
 sg13g2_nand2_1 _27645_ (.Y(_14033_),
    .A(_09558_),
    .B(net6592));
 sg13g2_nand2_1 _27646_ (.Y(_14034_),
    .A(_00399_),
    .B(net6519));
 sg13g2_o21ai_1 _27647_ (.B1(_14034_),
    .Y(_14035_),
    .A1(net6149),
    .A2(net6519));
 sg13g2_nand2_1 _27648_ (.Y(_14036_),
    .A(_00398_),
    .B(net6519));
 sg13g2_o21ai_1 _27649_ (.B1(_14036_),
    .Y(_14037_),
    .A1(net6147),
    .A2(net6519));
 sg13g2_nand2_1 _27650_ (.Y(_14038_),
    .A(_00397_),
    .B(net6518));
 sg13g2_o21ai_1 _27651_ (.B1(_14038_),
    .Y(_14039_),
    .A1(net6145),
    .A2(net6518));
 sg13g2_nand2_1 _27652_ (.Y(_14040_),
    .A(_00396_),
    .B(net6518));
 sg13g2_o21ai_1 _27653_ (.B1(_14040_),
    .Y(_14041_),
    .A1(net6144),
    .A2(net6518));
 sg13g2_nand2_1 _27654_ (.Y(_14042_),
    .A(_00395_),
    .B(net6522));
 sg13g2_o21ai_1 _27655_ (.B1(_14042_),
    .Y(_14043_),
    .A1(net6143),
    .A2(net6522));
 sg13g2_nand2_1 _27656_ (.Y(_14044_),
    .A(_00394_),
    .B(net6522));
 sg13g2_o21ai_1 _27657_ (.B1(_14044_),
    .Y(_14045_),
    .A1(_13506_),
    .A2(net6522));
 sg13g2_nand2_1 _27658_ (.Y(_14046_),
    .A(_00393_),
    .B(net6519));
 sg13g2_o21ai_1 _27659_ (.B1(_14046_),
    .Y(_14047_),
    .A1(net6141),
    .A2(net6519));
 sg13g2_nand2_1 _27660_ (.Y(_14048_),
    .A(_00392_),
    .B(net6521));
 sg13g2_o21ai_1 _27661_ (.B1(_14048_),
    .Y(_14049_),
    .A1(net6139),
    .A2(net6521));
 sg13g2_nand2_1 _27662_ (.Y(_14050_),
    .A(_00391_),
    .B(net6519));
 sg13g2_o21ai_1 _27663_ (.B1(_14050_),
    .Y(_14051_),
    .A1(net6138),
    .A2(net6519));
 sg13g2_nand2_1 _27664_ (.Y(_14052_),
    .A(_00390_),
    .B(net6518));
 sg13g2_o21ai_1 _27665_ (.B1(_14052_),
    .Y(_14053_),
    .A1(_13656_),
    .A2(net6518));
 sg13g2_mux2_1 _27666_ (.A0(_01209_),
    .A1(_01244_),
    .S(net7887),
    .X(_14054_));
 sg13g2_nand2_1 _27667_ (.Y(_14055_),
    .A(_00389_),
    .B(_14033_));
 sg13g2_o21ai_1 _27668_ (.B1(_14055_),
    .Y(_14056_),
    .A1(net6132),
    .A2(net6518));
 sg13g2_nand2_1 _27669_ (.Y(_14057_),
    .A(_00388_),
    .B(net6520));
 sg13g2_o21ai_1 _27670_ (.B1(_14057_),
    .Y(_14058_),
    .A1(net6133),
    .A2(net6520));
 sg13g2_nand2_1 _27671_ (.Y(_14059_),
    .A(_00387_),
    .B(net6520));
 sg13g2_o21ai_1 _27672_ (.B1(net7501),
    .Y(_14060_),
    .A1(net7509),
    .A2(_14054_));
 sg13g2_o21ai_1 _27673_ (.B1(_14059_),
    .Y(_14061_),
    .A1(net6156),
    .A2(net6520));
 sg13g2_nand2_1 _27674_ (.Y(_14062_),
    .A(_00386_),
    .B(net6520));
 sg13g2_nor4_1 _27675_ (.A(_13995_),
    .B(_14013_),
    .C(_14031_),
    .D(_14060_),
    .Y(_14063_));
 sg13g2_o21ai_1 _27676_ (.B1(_14062_),
    .Y(_14064_),
    .A1(net6155),
    .A2(net6520));
 sg13g2_nand2_1 _27677_ (.Y(_14065_),
    .A(_00385_),
    .B(net6520));
 sg13g2_o21ai_1 _27678_ (.B1(_14065_),
    .Y(_14066_),
    .A1(net6458),
    .A2(net6520));
 sg13g2_nand2_1 _27679_ (.Y(_14067_),
    .A(_00384_),
    .B(net6521));
 sg13g2_o21ai_1 _27680_ (.B1(_14067_),
    .Y(_14068_),
    .A1(net6153),
    .A2(net6521));
 sg13g2_nand2_1 _27681_ (.Y(_14069_),
    .A(_00383_),
    .B(net6521));
 sg13g2_o21ai_1 _27682_ (.B1(_14069_),
    .Y(_14070_),
    .A1(net6150),
    .A2(net6521));
 sg13g2_nand2_1 _27683_ (.Y(_14071_),
    .A(_00382_),
    .B(net6522));
 sg13g2_mux2_1 _27684_ (.A0(_00793_),
    .A1(_00825_),
    .S(net7883),
    .X(_14072_));
 sg13g2_o21ai_1 _27685_ (.B1(_14071_),
    .Y(_14073_),
    .A1(net6137),
    .A2(net6522));
 sg13g2_nand3_1 _27686_ (.B(net7471),
    .C(_14072_),
    .A(net7547),
    .Y(_14074_));
 sg13g2_a221oi_1 _27687_ (.B2(_13420_),
    .C1(net6668),
    .B1(net6701),
    .A1(\cs_registers_i.nmi_mode_i ),
    .Y(_14075_),
    .A2(net7079));
 sg13g2_a21oi_1 _27688_ (.A1(_02211_),
    .A2(net7079),
    .Y(_14076_),
    .B1(_13879_));
 sg13g2_mux2_1 _27689_ (.A0(_01948_),
    .A1(_01738_),
    .S(net6856),
    .X(_14077_));
 sg13g2_a22oi_1 _27690_ (.Y(_14078_),
    .B1(_14077_),
    .B2(net6660),
    .A2(net7038),
    .A1(_00471_));
 sg13g2_o21ai_1 _27691_ (.B1(_14078_),
    .Y(_14079_),
    .A1(net6459),
    .A2(net6632));
 sg13g2_mux2_1 _27692_ (.A0(_14079_),
    .A1(_00381_),
    .S(net6517),
    .X(_14080_));
 sg13g2_mux2_1 _27693_ (.A0(_01947_),
    .A1(_01737_),
    .S(net6856),
    .X(_14081_));
 sg13g2_a22oi_1 _27694_ (.Y(_14082_),
    .B1(_14081_),
    .B2(_13572_),
    .A2(net7037),
    .A1(_00470_));
 sg13g2_o21ai_1 _27695_ (.B1(_14082_),
    .Y(_14083_),
    .A1(_13436_),
    .A2(net6631));
 sg13g2_mux2_1 _27696_ (.A0(_14083_),
    .A1(_00380_),
    .S(net6516),
    .X(_14084_));
 sg13g2_mux2_1 _27697_ (.A0(_00857_),
    .A1(_00892_),
    .S(net7883),
    .X(_14085_));
 sg13g2_nand2_1 _27698_ (.Y(_14086_),
    .A(_01736_),
    .B(net6857));
 sg13g2_o21ai_1 _27699_ (.B1(_14086_),
    .Y(_14087_),
    .A1(_07450_),
    .A2(net6856));
 sg13g2_a22oi_1 _27700_ (.Y(_14088_),
    .B1(_14087_),
    .B2(net6661),
    .A2(net7038),
    .A1(_00469_));
 sg13g2_o21ai_1 _27701_ (.B1(_14088_),
    .Y(_14089_),
    .A1(net6132),
    .A2(net6632));
 sg13g2_mux2_1 _27702_ (.A0(_14089_),
    .A1(_00379_),
    .S(net6517),
    .X(_14090_));
 sg13g2_nand3_1 _27703_ (.B(net7462),
    .C(_14085_),
    .A(net7547),
    .Y(_14091_));
 sg13g2_mux2_1 _27704_ (.A0(_01945_),
    .A1(_01735_),
    .S(net6857),
    .X(_14092_));
 sg13g2_a22oi_1 _27705_ (.Y(_14093_),
    .B1(_14092_),
    .B2(net6659),
    .A2(_13895_),
    .A1(_00468_));
 sg13g2_o21ai_1 _27706_ (.B1(_14093_),
    .Y(_14094_),
    .A1(_13621_),
    .A2(_14076_));
 sg13g2_mux2_1 _27707_ (.A0(_14094_),
    .A1(_00378_),
    .S(net6515),
    .X(_14095_));
 sg13g2_mux2_1 _27708_ (.A0(_01944_),
    .A1(_01734_),
    .S(net6855),
    .X(_14096_));
 sg13g2_a22oi_1 _27709_ (.Y(_14097_),
    .B1(_14096_),
    .B2(net6659),
    .A2(net7038),
    .A1(_00467_));
 sg13g2_o21ai_1 _27710_ (.B1(_14097_),
    .Y(_14098_),
    .A1(net6533),
    .A2(net6632));
 sg13g2_mux2_1 _27711_ (.A0(_14098_),
    .A1(_00377_),
    .S(net6517),
    .X(_14099_));
 sg13g2_nor2_1 _27712_ (.A(_09320_),
    .B(_13566_),
    .Y(_14100_));
 sg13g2_and2_1 _27713_ (.A(_13646_),
    .B(_14100_),
    .X(_14101_));
 sg13g2_nand2_1 _27714_ (.Y(_14102_),
    .A(_13571_),
    .B(_13646_));
 sg13g2_mux2_1 _27715_ (.A0(_01943_),
    .A1(_01733_),
    .S(net6857),
    .X(_14103_));
 sg13g2_nand2_1 _27716_ (.Y(_14104_),
    .A(net7075),
    .B(_14103_));
 sg13g2_a21oi_1 _27717_ (.A1(_14102_),
    .A2(_14104_),
    .Y(_14105_),
    .B1(net6728));
 sg13g2_nor2_1 _27718_ (.A(_02211_),
    .B(_00466_),
    .Y(_14106_));
 sg13g2_nor2_1 _27719_ (.A(net7983),
    .B(_13646_),
    .Y(_14107_));
 sg13g2_nor3_1 _27720_ (.A(net7078),
    .B(_14106_),
    .C(_14107_),
    .Y(_14108_));
 sg13g2_mux2_1 _27721_ (.A0(_00998_),
    .A1(_01033_),
    .S(net7884),
    .X(_14109_));
 sg13g2_nor4_1 _27722_ (.A(net6513),
    .B(_14101_),
    .C(_14105_),
    .D(_14108_),
    .Y(_14110_));
 sg13g2_a21oi_1 _27723_ (.A1(_05742_),
    .A2(net6513),
    .Y(_14111_),
    .B1(_14110_));
 sg13g2_and2_1 _27724_ (.A(_13657_),
    .B(_14100_),
    .X(_14112_));
 sg13g2_nand2_1 _27725_ (.Y(_14113_),
    .A(_13571_),
    .B(_13657_));
 sg13g2_nand3_1 _27726_ (.B(net7525),
    .C(_14109_),
    .A(net7547),
    .Y(_14114_));
 sg13g2_nand2_1 _27727_ (.Y(_14115_),
    .A(_01732_),
    .B(net6857));
 sg13g2_o21ai_1 _27728_ (.B1(_14115_),
    .Y(_14116_),
    .A1(_07622_),
    .A2(net6857));
 sg13g2_nand2_1 _27729_ (.Y(_14117_),
    .A(net7075),
    .B(_14116_));
 sg13g2_a21oi_1 _27730_ (.A1(_14113_),
    .A2(_14117_),
    .Y(_14118_),
    .B1(net6728));
 sg13g2_nor2_1 _27731_ (.A(net7983),
    .B(_13657_),
    .Y(_14119_));
 sg13g2_nor2_1 _27732_ (.A(net7078),
    .B(_14119_),
    .Y(_14120_));
 sg13g2_o21ai_1 _27733_ (.B1(_14120_),
    .Y(_14121_),
    .A1(_02211_),
    .A2(_00465_));
 sg13g2_nor3_1 _27734_ (.A(net6513),
    .B(_14112_),
    .C(_14118_),
    .Y(_14122_));
 sg13g2_a22oi_1 _27735_ (.Y(_14123_),
    .B1(_14121_),
    .B2(_14122_),
    .A2(net6513),
    .A1(_05744_));
 sg13g2_mux2_1 _27736_ (.A0(_00927_),
    .A1(_00963_),
    .S(net7884),
    .X(_14124_));
 sg13g2_mux2_1 _27737_ (.A0(_01941_),
    .A1(_01731_),
    .S(net6853),
    .X(_14125_));
 sg13g2_a22oi_1 _27738_ (.Y(_14126_),
    .B1(_14125_),
    .B2(net6660),
    .A2(net7038),
    .A1(_00464_));
 sg13g2_o21ai_1 _27739_ (.B1(_14126_),
    .Y(_14127_),
    .A1(net6158),
    .A2(net6632));
 sg13g2_mux2_1 _27740_ (.A0(_14127_),
    .A1(_00374_),
    .S(net6517),
    .X(_14128_));
 sg13g2_nand3_1 _27741_ (.B(net7512),
    .C(_14124_),
    .A(net7547),
    .Y(_14129_));
 sg13g2_mux2_1 _27742_ (.A0(_01940_),
    .A1(_01730_),
    .S(net6853),
    .X(_14130_));
 sg13g2_a22oi_1 _27743_ (.Y(_14131_),
    .B1(_14130_),
    .B2(net6666),
    .A2(net7034),
    .A1(_00463_));
 sg13g2_o21ai_1 _27744_ (.B1(_14131_),
    .Y(_14132_),
    .A1(_13446_),
    .A2(net6629));
 sg13g2_mux2_1 _27745_ (.A0(_14132_),
    .A1(_00373_),
    .S(net6514),
    .X(_14133_));
 sg13g2_inv_1 _27746_ (.Y(_14134_),
    .A(_14135_));
 sg13g2_mux2_1 _27747_ (.A0(_01939_),
    .A1(_01729_),
    .S(net6857),
    .X(_14135_));
 sg13g2_nor2_1 _27748_ (.A(net7075),
    .B(net6131),
    .Y(_14136_));
 sg13g2_a21oi_1 _27749_ (.A1(net7075),
    .A2(_14134_),
    .Y(_14137_),
    .B1(net6728));
 sg13g2_o21ai_1 _27750_ (.B1(_14137_),
    .Y(_14138_),
    .A1(net7075),
    .A2(net6131));
 sg13g2_nor2_1 _27751_ (.A(net7982),
    .B(net6131),
    .Y(_14139_));
 sg13g2_a21oi_1 _27752_ (.A1(net7982),
    .A2(_05464_),
    .Y(_14140_),
    .B1(_14139_));
 sg13g2_a221oi_1 _27753_ (.B2(_09320_),
    .C1(net6513),
    .B1(_14140_),
    .A1(net6131),
    .Y(_14141_),
    .A2(_14100_));
 sg13g2_a22oi_1 _27754_ (.Y(_14142_),
    .B1(_14138_),
    .B2(_14141_),
    .A2(net6513),
    .A1(_05752_));
 sg13g2_mux2_1 _27755_ (.A0(_01938_),
    .A1(_01728_),
    .S(net6853),
    .X(_14143_));
 sg13g2_a22oi_1 _27756_ (.Y(_14144_),
    .B1(_14143_),
    .B2(net6666),
    .A2(net7034),
    .A1(_00461_));
 sg13g2_o21ai_1 _27757_ (.B1(_14144_),
    .Y(_14145_),
    .A1(net6155),
    .A2(net6629));
 sg13g2_mux2_1 _27758_ (.A0(_14145_),
    .A1(_00371_),
    .S(net6514),
    .X(_14146_));
 sg13g2_mux2_1 _27759_ (.A0(_01561_),
    .A1(_01596_),
    .S(net7892),
    .X(_14147_));
 sg13g2_mux2_1 _27760_ (.A0(_01937_),
    .A1(_01727_),
    .S(net6853),
    .X(_14148_));
 sg13g2_a22oi_1 _27761_ (.Y(_14149_),
    .B1(_14148_),
    .B2(net6666),
    .A2(net7034),
    .A1(_00460_));
 sg13g2_o21ai_1 _27762_ (.B1(_14149_),
    .Y(_14150_),
    .A1(_13458_),
    .A2(net6629));
 sg13g2_nand2_1 _27763_ (.Y(_14151_),
    .A(net7450),
    .B(_14147_));
 sg13g2_mux2_1 _27764_ (.A0(_14150_),
    .A1(_00370_),
    .S(net6514),
    .X(_14152_));
 sg13g2_mux2_1 _27765_ (.A0(_01936_),
    .A1(_01726_),
    .S(net6854),
    .X(_14153_));
 sg13g2_a22oi_1 _27766_ (.Y(_14154_),
    .B1(_14153_),
    .B2(net6664),
    .A2(net7035),
    .A1(_00459_));
 sg13g2_o21ai_1 _27767_ (.B1(_14154_),
    .Y(_14155_),
    .A1(net6153),
    .A2(net6630));
 sg13g2_mux2_1 _27768_ (.A0(_14155_),
    .A1(_00369_),
    .S(net6515),
    .X(_14156_));
 sg13g2_mux2_1 _27769_ (.A0(_01935_),
    .A1(_01725_),
    .S(net6854),
    .X(_14157_));
 sg13g2_a22oi_1 _27770_ (.Y(_14158_),
    .B1(_14157_),
    .B2(net6664),
    .A2(net7034),
    .A1(_00458_));
 sg13g2_o21ai_1 _27771_ (.B1(_14158_),
    .Y(_14159_),
    .A1(net6150),
    .A2(net6629));
 sg13g2_mux2_1 _27772_ (.A0(_14159_),
    .A1(_00368_),
    .S(net6514),
    .X(_14160_));
 sg13g2_mux2_1 _27773_ (.A0(_01934_),
    .A1(_01724_),
    .S(net6855),
    .X(_14161_));
 sg13g2_mux2_1 _27774_ (.A0(_01491_),
    .A1(_01526_),
    .S(net7892),
    .X(_14162_));
 sg13g2_a22oi_1 _27775_ (.Y(_14163_),
    .B1(_14161_),
    .B2(net6664),
    .A2(net7034),
    .A1(_00457_));
 sg13g2_o21ai_1 _27776_ (.B1(_14163_),
    .Y(_14164_),
    .A1(_13477_),
    .A2(net6629));
 sg13g2_mux2_1 _27777_ (.A0(_14164_),
    .A1(_00367_),
    .S(net6514),
    .X(_14165_));
 sg13g2_mux2_1 _27778_ (.A0(_01933_),
    .A1(_01723_),
    .S(net6854),
    .X(_14166_));
 sg13g2_nand3_1 _27779_ (.B(net7495),
    .C(_14162_),
    .A(net7512),
    .Y(_14167_));
 sg13g2_a22oi_1 _27780_ (.Y(_14168_),
    .B1(_14166_),
    .B2(net6664),
    .A2(net7035),
    .A1(_00456_));
 sg13g2_o21ai_1 _27781_ (.B1(_14168_),
    .Y(_14169_),
    .A1(net6147),
    .A2(net6630));
 sg13g2_mux2_1 _27782_ (.A0(_14169_),
    .A1(_00366_),
    .S(net6515),
    .X(_14170_));
 sg13g2_mux2_1 _27783_ (.A0(_01932_),
    .A1(_01722_),
    .S(net6855),
    .X(_14171_));
 sg13g2_a22oi_1 _27784_ (.Y(_14172_),
    .B1(_14171_),
    .B2(net6663),
    .A2(net7035),
    .A1(_00455_));
 sg13g2_o21ai_1 _27785_ (.B1(_14172_),
    .Y(_14173_),
    .A1(net6145),
    .A2(net6630));
 sg13g2_mux2_1 _27786_ (.A0(_14173_),
    .A1(_00365_),
    .S(net6515),
    .X(_14174_));
 sg13g2_mux2_1 _27787_ (.A0(_01931_),
    .A1(_01721_),
    .S(net6855),
    .X(_14175_));
 sg13g2_a22oi_1 _27788_ (.Y(_14176_),
    .B1(_14175_),
    .B2(net6663),
    .A2(net7035),
    .A1(_00454_));
 sg13g2_o21ai_1 _27789_ (.B1(_14176_),
    .Y(_14177_),
    .A1(net6144),
    .A2(net6630));
 sg13g2_mux2_1 _27790_ (.A0(_14177_),
    .A1(_00364_),
    .S(net6515),
    .X(_14178_));
 sg13g2_mux2_1 _27791_ (.A0(_01930_),
    .A1(_01720_),
    .S(net6855),
    .X(_14179_));
 sg13g2_a22oi_1 _27792_ (.Y(_14180_),
    .B1(_14179_),
    .B2(net6664),
    .A2(net7035),
    .A1(_00453_));
 sg13g2_o21ai_1 _27793_ (.B1(_14180_),
    .Y(_14181_),
    .A1(net6143),
    .A2(net6630));
 sg13g2_mux2_1 _27794_ (.A0(_14181_),
    .A1(_00363_),
    .S(net6515),
    .X(_14182_));
 sg13g2_mux2_1 _27795_ (.A0(_01420_),
    .A1(_01455_),
    .S(net7892),
    .X(_14183_));
 sg13g2_mux2_1 _27796_ (.A0(_01929_),
    .A1(_01719_),
    .S(net6855),
    .X(_14184_));
 sg13g2_a22oi_1 _27797_ (.Y(_14185_),
    .B1(_14184_),
    .B2(net6663),
    .A2(net7035),
    .A1(_00452_));
 sg13g2_o21ai_1 _27798_ (.B1(_14185_),
    .Y(_14186_),
    .A1(_13506_),
    .A2(net6630));
 sg13g2_mux2_1 _27799_ (.A0(_14186_),
    .A1(_00362_),
    .S(net6515),
    .X(_14187_));
 sg13g2_nand3_1 _27800_ (.B(net7462),
    .C(_14183_),
    .A(net7496),
    .Y(_14188_));
 sg13g2_inv_1 _27801_ (.Y(_14189_),
    .A(_14190_));
 sg13g2_nand2_1 _27802_ (.Y(_14190_),
    .A(_13571_),
    .B(_13780_));
 sg13g2_mux2_1 _27803_ (.A0(_01928_),
    .A1(_01718_),
    .S(net6857),
    .X(_14191_));
 sg13g2_a21oi_1 _27804_ (.A1(_13570_),
    .A2(_14191_),
    .Y(_14192_),
    .B1(_14189_));
 sg13g2_nand2_1 _27805_ (.Y(_14193_),
    .A(net7983),
    .B(_00451_));
 sg13g2_o21ai_1 _27806_ (.B1(_14193_),
    .Y(_14194_),
    .A1(net7983),
    .A2(_13779_));
 sg13g2_a22oi_1 _27807_ (.Y(_14195_),
    .B1(_14194_),
    .B2(_09320_),
    .A2(_14100_),
    .A1(_13780_));
 sg13g2_o21ai_1 _27808_ (.B1(_14195_),
    .Y(_14196_),
    .A1(net6728),
    .A2(_14192_));
 sg13g2_mux2_1 _27809_ (.A0(_14196_),
    .A1(_00361_),
    .S(net6513),
    .X(_14197_));
 sg13g2_mux2_1 _27810_ (.A0(_01927_),
    .A1(_01717_),
    .S(net6854),
    .X(_14198_));
 sg13g2_mux2_1 _27811_ (.A0(_01350_),
    .A1(_01385_),
    .S(net7890),
    .X(_14199_));
 sg13g2_a22oi_1 _27812_ (.Y(_14200_),
    .B1(_14198_),
    .B2(net6666),
    .A2(net7034),
    .A1(_00450_));
 sg13g2_o21ai_1 _27813_ (.B1(_14200_),
    .Y(_14201_),
    .A1(_13511_),
    .A2(net6629));
 sg13g2_mux2_1 _27814_ (.A0(_14201_),
    .A1(_00360_),
    .S(net6514),
    .X(_14202_));
 sg13g2_nand2_1 _27815_ (.Y(_14203_),
    .A(_01716_),
    .B(net6854));
 sg13g2_nand3_1 _27816_ (.B(net7471),
    .C(_14199_),
    .A(net7496),
    .Y(_14204_));
 sg13g2_o21ai_1 _27817_ (.B1(_14203_),
    .Y(_14205_),
    .A1(_08227_),
    .A2(net6854));
 sg13g2_a22oi_1 _27818_ (.Y(_14206_),
    .B1(_14205_),
    .B2(net6666),
    .A2(net7034),
    .A1(_00449_));
 sg13g2_o21ai_1 _27819_ (.B1(_14206_),
    .Y(_14207_),
    .A1(net6140),
    .A2(net6629));
 sg13g2_mux2_1 _27820_ (.A0(_14207_),
    .A1(_00359_),
    .S(net6514),
    .X(_14208_));
 sg13g2_mux2_1 _27821_ (.A0(_01925_),
    .A1(_01715_),
    .S(net6853),
    .X(_14209_));
 sg13g2_a22oi_1 _27822_ (.Y(_14210_),
    .B1(_14209_),
    .B2(net6666),
    .A2(net7034),
    .A1(_00448_));
 sg13g2_o21ai_1 _27823_ (.B1(_14210_),
    .Y(_14211_),
    .A1(net6138),
    .A2(net6629));
 sg13g2_mux2_1 _27824_ (.A0(_14211_),
    .A1(_00358_),
    .S(net6514),
    .X(_14212_));
 sg13g2_mux2_1 _27825_ (.A0(_01924_),
    .A1(_01714_),
    .S(net6853),
    .X(_14213_));
 sg13g2_a22oi_1 _27826_ (.Y(_14214_),
    .B1(_14213_),
    .B2(net6660),
    .A2(net7038),
    .A1(_00447_));
 sg13g2_o21ai_1 _27827_ (.B1(_14214_),
    .Y(_14215_),
    .A1(_13527_),
    .A2(net6632));
 sg13g2_mux2_1 _27828_ (.A0(_14215_),
    .A1(_00357_),
    .S(net6517),
    .X(_14216_));
 sg13g2_mux2_1 _27829_ (.A0(_01923_),
    .A1(_01713_),
    .S(net6855),
    .X(_14217_));
 sg13g2_a22oi_1 _27830_ (.Y(_14218_),
    .B1(_14217_),
    .B2(net6659),
    .A2(_13895_),
    .A1(_00446_));
 sg13g2_o21ai_1 _27831_ (.B1(_14218_),
    .Y(_14219_),
    .A1(net6543),
    .A2(net6632));
 sg13g2_mux2_1 _27832_ (.A0(_14219_),
    .A1(_00356_),
    .S(net6513),
    .X(_14220_));
 sg13g2_mux2_1 _27833_ (.A0(_01922_),
    .A1(_01712_),
    .S(net6856),
    .X(_14221_));
 sg13g2_a22oi_1 _27834_ (.Y(_14222_),
    .B1(_14221_),
    .B2(_13572_),
    .A2(net7037),
    .A1(_00445_));
 sg13g2_o21ai_1 _27835_ (.B1(_14222_),
    .Y(_14223_),
    .A1(net6542),
    .A2(net6631));
 sg13g2_mux2_1 _27836_ (.A0(_14223_),
    .A1(_00355_),
    .S(net6516),
    .X(_14224_));
 sg13g2_mux2_1 _27837_ (.A0(_01921_),
    .A1(_01711_),
    .S(net6856),
    .X(_14225_));
 sg13g2_a22oi_1 _27838_ (.Y(_14226_),
    .B1(_14225_),
    .B2(net6669),
    .A2(net7037),
    .A1(_00444_));
 sg13g2_o21ai_1 _27839_ (.B1(_14226_),
    .Y(_14227_),
    .A1(net6136),
    .A2(net6631));
 sg13g2_nand4_1 _27840_ (.B(_14114_),
    .C(_14129_),
    .A(_14074_),
    .Y(_14228_),
    .D(_14188_));
 sg13g2_mux2_1 _27841_ (.A0(_14227_),
    .A1(_00354_),
    .S(net6516),
    .X(_14229_));
 sg13g2_mux2_1 _27842_ (.A0(_01920_),
    .A1(_01710_),
    .S(net6856),
    .X(_14230_));
 sg13g2_a22oi_1 _27843_ (.Y(_14231_),
    .B1(_14230_),
    .B2(net6669),
    .A2(net7037),
    .A1(_00443_));
 sg13g2_o21ai_1 _27844_ (.B1(_14231_),
    .Y(_14232_),
    .A1(_13547_),
    .A2(net6631));
 sg13g2_mux2_1 _27845_ (.A0(_14232_),
    .A1(_00353_),
    .S(net6516),
    .X(_14233_));
 sg13g2_mux2_1 _27846_ (.A0(_01919_),
    .A1(_01709_),
    .S(net6853),
    .X(_14234_));
 sg13g2_a22oi_1 _27847_ (.Y(_14235_),
    .B1(_14234_),
    .B2(net6660),
    .A2(net7038),
    .A1(_00442_));
 sg13g2_o21ai_1 _27848_ (.B1(_14235_),
    .Y(_14236_),
    .A1(net6134),
    .A2(net6632));
 sg13g2_mux2_1 _27849_ (.A0(_14236_),
    .A1(_00352_),
    .S(net6517),
    .X(_14237_));
 sg13g2_nand2_1 _27850_ (.Y(_14238_),
    .A(_01708_),
    .B(net6856));
 sg13g2_o21ai_1 _27851_ (.B1(_14238_),
    .Y(_14239_),
    .A1(_08414_),
    .A2(net6856));
 sg13g2_nand4_1 _27852_ (.B(_14151_),
    .C(_14167_),
    .A(_14091_),
    .Y(_14240_),
    .D(_14204_));
 sg13g2_a22oi_1 _27853_ (.Y(_14241_),
    .B1(_14239_),
    .B2(net6669),
    .A2(net7037),
    .A1(_00441_));
 sg13g2_o21ai_1 _27854_ (.B1(_14241_),
    .Y(_14242_),
    .A1(net6455),
    .A2(net6631));
 sg13g2_mux2_1 _27855_ (.A0(_14242_),
    .A1(_00351_),
    .S(net6516),
    .X(_14243_));
 sg13g2_a22oi_1 _27856_ (.Y(_14244_),
    .B1(_14075_),
    .B2(_00350_),
    .A2(net7036),
    .A1(_00440_));
 sg13g2_inv_1 _27857_ (.Y(_14245_),
    .A(_14244_));
 sg13g2_a221oi_1 _27858_ (.B2(net6592),
    .C1(net6668),
    .B1(_09565_),
    .A1(\cs_registers_i.nmi_mode_i ),
    .Y(_14246_),
    .A2(net7079));
 sg13g2_a22oi_1 _27859_ (.Y(_14247_),
    .B1(net7036),
    .B2(_00437_),
    .A2(_13568_),
    .A1(_07087_));
 sg13g2_o21ai_1 _27860_ (.B1(_14247_),
    .Y(_14248_),
    .A1(net6158),
    .A2(net6630));
 sg13g2_mux2_1 _27861_ (.A0(_14248_),
    .A1(_00349_),
    .S(net6512),
    .X(_14249_));
 sg13g2_nand2_1 _27862_ (.Y(_14250_),
    .A(_07735_),
    .B(net7075));
 sg13g2_a21oi_1 _27863_ (.A1(_14102_),
    .A2(_14250_),
    .Y(_14251_),
    .B1(net6728));
 sg13g2_nor4_1 _27864_ (.A(_13978_),
    .B(_14063_),
    .C(_14228_),
    .D(_14240_),
    .Y(_14252_));
 sg13g2_or4_1 _27865_ (.A(_13978_),
    .B(_14063_),
    .C(_14228_),
    .D(_14240_),
    .X(_14253_));
 sg13g2_nor2_1 _27866_ (.A(_02211_),
    .B(_00436_),
    .Y(_14254_));
 sg13g2_nor3_1 _27867_ (.A(net7078),
    .B(_14107_),
    .C(_14254_),
    .Y(_14255_));
 sg13g2_nor4_1 _27868_ (.A(_14101_),
    .B(net6512),
    .C(_14251_),
    .D(_14255_),
    .Y(_14256_));
 sg13g2_a21oi_1 _27869_ (.A1(_05827_),
    .A2(net6512),
    .Y(_14257_),
    .B1(_14256_));
 sg13g2_nand2_1 _27870_ (.Y(_14258_),
    .A(_07751_),
    .B(net7075));
 sg13g2_a21oi_1 _27871_ (.A1(_14113_),
    .A2(_14258_),
    .Y(_14259_),
    .B1(net6728));
 sg13g2_nor2_1 _27872_ (.A(_02211_),
    .B(_00435_),
    .Y(_14260_));
 sg13g2_nor3_1 _27873_ (.A(net7078),
    .B(_14119_),
    .C(_14260_),
    .Y(_14261_));
 sg13g2_nor4_1 _27874_ (.A(_14112_),
    .B(net6512),
    .C(_14259_),
    .D(_14261_),
    .Y(_14262_));
 sg13g2_a21oi_1 _27875_ (.A1(_05829_),
    .A2(net6512),
    .Y(_14263_),
    .B1(_14262_));
 sg13g2_nand2b_1 _27876_ (.Y(_14264_),
    .B(net7998),
    .A_N(_01637_));
 sg13g2_a21oi_1 _27877_ (.A1(net7982),
    .A2(_05552_),
    .Y(_14265_),
    .B1(_14139_));
 sg13g2_a21oi_1 _27878_ (.A1(_07763_),
    .A2(net7075),
    .Y(_14266_),
    .B1(_14136_));
 sg13g2_o21ai_1 _27879_ (.B1(_14264_),
    .Y(_14267_),
    .A1(_01660_),
    .A2(_09260_));
 sg13g2_a22oi_1 _27880_ (.Y(_14268_),
    .B1(_14265_),
    .B2(_09320_),
    .A2(_14100_),
    .A1(net6131));
 sg13g2_a21oi_1 _27881_ (.A1(_13566_),
    .A2(_14266_),
    .Y(_14269_),
    .B1(net6512));
 sg13g2_a22oi_1 _27882_ (.Y(_14270_),
    .B1(_14268_),
    .B2(_14269_),
    .A2(net6512),
    .A1(_05830_));
 sg13g2_inv_1 _27883_ (.Y(_14271_),
    .A(_14272_));
 sg13g2_o21ai_1 _27884_ (.B1(_14190_),
    .Y(_14272_),
    .A1(_07784_),
    .A2(_13571_));
 sg13g2_nand2_1 _27885_ (.Y(_14273_),
    .A(net7983),
    .B(_00433_));
 sg13g2_o21ai_1 _27886_ (.B1(_14273_),
    .Y(_14274_),
    .A1(net7983),
    .A2(net6454));
 sg13g2_a221oi_1 _27887_ (.B2(net8005),
    .C1(_14267_),
    .B1(net7275),
    .A1(_09275_),
    .Y(_14275_),
    .A2(net7074));
 sg13g2_a22oi_1 _27888_ (.Y(_14276_),
    .B1(_14274_),
    .B2(_09320_),
    .A2(_14100_),
    .A1(_13780_));
 sg13g2_o21ai_1 _27889_ (.B1(_14276_),
    .Y(_14277_),
    .A1(net6728),
    .A2(_14271_));
 sg13g2_mux2_1 _27890_ (.A0(_14277_),
    .A1(_00345_),
    .S(net6512),
    .X(_14278_));
 sg13g2_a22oi_1 _27891_ (.Y(_14279_),
    .B1(net7036),
    .B2(_00432_),
    .A2(net6662),
    .A1(_07837_));
 sg13g2_o21ai_1 _27892_ (.B1(_14279_),
    .Y(_14280_),
    .A1(_13874_),
    .A2(_14076_));
 sg13g2_mux2_1 _27893_ (.A0(_14280_),
    .A1(_00344_),
    .S(_14246_),
    .X(_14281_));
 sg13g2_nand2_1 _27894_ (.Y(_14282_),
    .A(net6692),
    .B(_13420_));
 sg13g2_nand2_1 _27895_ (.Y(_14283_),
    .A(_00343_),
    .B(net6508));
 sg13g2_o21ai_1 _27896_ (.B1(_14283_),
    .Y(_14284_),
    .A1(_13431_),
    .A2(net6508));
 sg13g2_nand2_1 _27897_ (.Y(_14285_),
    .A(_00342_),
    .B(net6511));
 sg13g2_o21ai_1 _27898_ (.B1(_14285_),
    .Y(_14286_),
    .A1(net6159),
    .A2(net6509));
 sg13g2_nand2_1 _27899_ (.Y(_14287_),
    .A(_00341_),
    .B(net6507));
 sg13g2_nor2_1 _27900_ (.A(net7364),
    .B(_14275_),
    .Y(_14288_));
 sg13g2_o21ai_1 _27901_ (.B1(_14287_),
    .Y(_14289_),
    .A1(net6132),
    .A2(net6507));
 sg13g2_nand2_1 _27902_ (.Y(_14290_),
    .A(_00340_),
    .B(net6506));
 sg13g2_a21oi_1 _27903_ (.A1(net6917),
    .A2(_13838_),
    .Y(_14291_),
    .B1(_14288_));
 sg13g2_o21ai_1 _27904_ (.B1(_14290_),
    .Y(_14292_),
    .A1(_13621_),
    .A2(net6506));
 sg13g2_nand2_1 _27905_ (.Y(_14293_),
    .A(_00339_),
    .B(_14282_));
 sg13g2_o21ai_1 _27906_ (.B1(_14293_),
    .Y(_14294_),
    .A1(net6533),
    .A2(_14282_));
 sg13g2_nand2_1 _27907_ (.Y(_14295_),
    .A(_00338_),
    .B(net6505));
 sg13g2_o21ai_1 _27908_ (.B1(_14295_),
    .Y(_14296_),
    .A1(_13645_),
    .A2(net6505));
 sg13g2_nand2_1 _27909_ (.Y(_14297_),
    .A(_00337_),
    .B(net6505));
 sg13g2_o21ai_1 _27910_ (.B1(_14297_),
    .Y(_14298_),
    .A1(_13656_),
    .A2(net6505));
 sg13g2_nand2_1 _27911_ (.Y(_14299_),
    .A(_00336_),
    .B(net6508));
 sg13g2_o21ai_1 _27912_ (.B1(_14291_),
    .Y(_14300_),
    .A1(_08228_),
    .A2(_13838_));
 sg13g2_o21ai_1 _27913_ (.B1(_14299_),
    .Y(_14301_),
    .A1(net6158),
    .A2(net6508));
 sg13g2_nand2_1 _27914_ (.Y(_14302_),
    .A(_00335_),
    .B(net6508));
 sg13g2_o21ai_1 _27915_ (.B1(_14302_),
    .Y(_14303_),
    .A1(net6156),
    .A2(net6508));
 sg13g2_nand2_1 _27916_ (.Y(_14304_),
    .A(_00334_),
    .B(net6507));
 sg13g2_o21ai_1 _27917_ (.B1(_14304_),
    .Y(_14305_),
    .A1(_13704_),
    .A2(net6507));
 sg13g2_nand2_1 _27918_ (.Y(_14306_),
    .A(_00333_),
    .B(net6510));
 sg13g2_o21ai_1 _27919_ (.B1(_14306_),
    .Y(_14307_),
    .A1(net6155),
    .A2(net6510));
 sg13g2_nand2_1 _27920_ (.Y(_14308_),
    .A(_00332_),
    .B(net6510));
 sg13g2_o21ai_1 _27921_ (.B1(_14308_),
    .Y(_14309_),
    .A1(net6458),
    .A2(net6510));
 sg13g2_nand2_1 _27922_ (.Y(_14310_),
    .A(_00331_),
    .B(net6504));
 sg13g2_o21ai_1 _27923_ (.B1(_14310_),
    .Y(_14311_),
    .A1(net6152),
    .A2(net6504));
 sg13g2_nand2_1 _27924_ (.Y(_14312_),
    .A(_00330_),
    .B(net6503));
 sg13g2_o21ai_1 _27925_ (.B1(_14312_),
    .Y(_14313_),
    .A1(net6151),
    .A2(net6503));
 sg13g2_nand2_1 _27926_ (.Y(_14314_),
    .A(_00329_),
    .B(net6511));
 sg13g2_o21ai_1 _27927_ (.B1(_14314_),
    .Y(_14315_),
    .A1(net6149),
    .A2(net6511));
 sg13g2_nand2_1 _27928_ (.Y(_14316_),
    .A(_00328_),
    .B(net6502));
 sg13g2_o21ai_1 _27929_ (.B1(_14316_),
    .Y(_14317_),
    .A1(net6148),
    .A2(net6502));
 sg13g2_nand2_1 _27930_ (.Y(_14318_),
    .A(_00327_),
    .B(net6502));
 sg13g2_o21ai_1 _27931_ (.B1(_14318_),
    .Y(_14319_),
    .A1(net6146),
    .A2(net6502));
 sg13g2_nand2_1 _27932_ (.Y(_14320_),
    .A(_00326_),
    .B(net6502));
 sg13g2_o21ai_1 _27933_ (.B1(_14320_),
    .Y(_14321_),
    .A1(_13495_),
    .A2(net6504));
 sg13g2_nand2_1 _27934_ (.Y(_14322_),
    .A(_00325_),
    .B(net6502));
 sg13g2_o21ai_1 _27935_ (.B1(_14322_),
    .Y(_14323_),
    .A1(net6143),
    .A2(net6502));
 sg13g2_nand2_1 _27936_ (.Y(_14324_),
    .A(_00324_),
    .B(net6503));
 sg13g2_o21ai_1 _27937_ (.B1(_14324_),
    .Y(_14325_),
    .A1(_13506_),
    .A2(net6503));
 sg13g2_nand2_1 _27938_ (.Y(_14326_),
    .A(_00323_),
    .B(net6506));
 sg13g2_o21ai_1 _27939_ (.B1(_14326_),
    .Y(_14327_),
    .A1(net6454),
    .A2(net6506));
 sg13g2_nand2_1 _27940_ (.Y(_14328_),
    .A(_00322_),
    .B(net6503));
 sg13g2_o21ai_1 _27941_ (.B1(_14328_),
    .Y(_14329_),
    .A1(net6141),
    .A2(net6503));
 sg13g2_nand2_1 _27942_ (.Y(_14330_),
    .A(_00321_),
    .B(net6510));
 sg13g2_o21ai_1 _27943_ (.B1(_14330_),
    .Y(_14331_),
    .A1(net6139),
    .A2(net6510));
 sg13g2_nand2_1 _27944_ (.Y(_14332_),
    .A(_00320_),
    .B(net6510));
 sg13g2_mux4_1 _27945_ (.S0(net7787),
    .A0(_00794_),
    .A1(_00826_),
    .A2(_00858_),
    .A3(_00893_),
    .S1(net7727),
    .X(_14333_));
 sg13g2_o21ai_1 _27946_ (.B1(_14332_),
    .Y(_14334_),
    .A1(net6138),
    .A2(net6510));
 sg13g2_nand2_1 _27947_ (.Y(_14335_),
    .A(_00319_),
    .B(net6503));
 sg13g2_o21ai_1 _27948_ (.B1(_14335_),
    .Y(_14336_),
    .A1(net6137),
    .A2(net6503));
 sg13g2_nor2_1 _27949_ (.A(net7713),
    .B(_14333_),
    .Y(_14337_));
 sg13g2_nand2_1 _27950_ (.Y(_14338_),
    .A(_00318_),
    .B(net6505));
 sg13g2_o21ai_1 _27951_ (.B1(_14338_),
    .Y(_14339_),
    .A1(_13532_),
    .A2(net6505));
 sg13g2_nand2_1 _27952_ (.Y(_14340_),
    .A(_00317_),
    .B(net6504));
 sg13g2_o21ai_1 _27953_ (.B1(_14340_),
    .Y(_14341_),
    .A1(net6542),
    .A2(net6504));
 sg13g2_nand2_1 _27954_ (.Y(_14342_),
    .A(_00316_),
    .B(net6508));
 sg13g2_o21ai_1 _27955_ (.B1(_14342_),
    .Y(_14343_),
    .A1(net6135),
    .A2(net6508));
 sg13g2_nand2_1 _27956_ (.Y(_14344_),
    .A(_00315_),
    .B(net6507));
 sg13g2_o21ai_1 _27957_ (.B1(_14344_),
    .Y(_14345_),
    .A1(net6457),
    .A2(net6507));
 sg13g2_nand2_1 _27958_ (.Y(_14346_),
    .A(_00314_),
    .B(net6509));
 sg13g2_o21ai_1 _27959_ (.B1(_14346_),
    .Y(_14347_),
    .A1(net6133),
    .A2(net6509));
 sg13g2_nand2_1 _27960_ (.Y(_14348_),
    .A(_00313_),
    .B(net6509));
 sg13g2_o21ai_1 _27961_ (.B1(_14348_),
    .Y(_14349_),
    .A1(net6455),
    .A2(net6509));
 sg13g2_nand2_1 _27962_ (.Y(_14350_),
    .A(_00312_),
    .B(net6505));
 sg13g2_mux2_1 _27963_ (.A0(_00999_),
    .A1(_01034_),
    .S(net7784),
    .X(_14351_));
 sg13g2_o21ai_1 _27964_ (.B1(_14350_),
    .Y(_14352_),
    .A1(_13874_),
    .A2(net6505));
 sg13g2_nand2_1 _27965_ (.Y(_14353_),
    .A(net6695),
    .B(_13420_));
 sg13g2_nand2_1 _27966_ (.Y(_14354_),
    .A(_00311_),
    .B(net6496));
 sg13g2_o21ai_1 _27967_ (.B1(_14354_),
    .Y(_14355_),
    .A1(_13431_),
    .A2(net6496));
 sg13g2_nand2_1 _27968_ (.Y(_14356_),
    .A(_00310_),
    .B(_14353_));
 sg13g2_o21ai_1 _27969_ (.B1(_14356_),
    .Y(_14357_),
    .A1(net6159),
    .A2(_14353_));
 sg13g2_nand2_1 _27970_ (.Y(_14358_),
    .A(_00309_),
    .B(net6499));
 sg13g2_nor2_1 _27971_ (.A(_08522_),
    .B(_14351_),
    .Y(_14359_));
 sg13g2_o21ai_1 _27972_ (.B1(_14358_),
    .Y(_14360_),
    .A1(net6132),
    .A2(net6500));
 sg13g2_nand2_1 _27973_ (.Y(_14361_),
    .A(_00308_),
    .B(net6494));
 sg13g2_o21ai_1 _27974_ (.B1(_14361_),
    .Y(_14362_),
    .A1(_13621_),
    .A2(net6494));
 sg13g2_nand2_1 _27975_ (.Y(_14363_),
    .A(_00307_),
    .B(_14353_));
 sg13g2_o21ai_1 _27976_ (.B1(_14363_),
    .Y(_14364_),
    .A1(net6533),
    .A2(_14353_));
 sg13g2_nand2_1 _27977_ (.Y(_14365_),
    .A(_00306_),
    .B(net6493));
 sg13g2_o21ai_1 _27978_ (.B1(_14365_),
    .Y(_14366_),
    .A1(_13645_),
    .A2(net6493));
 sg13g2_nand2_1 _27979_ (.Y(_14367_),
    .A(_00305_),
    .B(net6493));
 sg13g2_o21ai_1 _27980_ (.B1(_14367_),
    .Y(_14368_),
    .A1(_13656_),
    .A2(net6493));
 sg13g2_nand2_1 _27981_ (.Y(_14369_),
    .A(_00304_),
    .B(net6496));
 sg13g2_o21ai_1 _27982_ (.B1(_14369_),
    .Y(_14370_),
    .A1(net6158),
    .A2(net6496));
 sg13g2_nand2_1 _27983_ (.Y(_14371_),
    .A(_00303_),
    .B(net6496));
 sg13g2_o21ai_1 _27984_ (.B1(_14371_),
    .Y(_14372_),
    .A1(net6156),
    .A2(net6496));
 sg13g2_nand2_1 _27985_ (.Y(_14373_),
    .A(_00302_),
    .B(net6494));
 sg13g2_mux2_1 _27986_ (.A0(_00929_),
    .A1(_00964_),
    .S(net7784),
    .X(_14374_));
 sg13g2_o21ai_1 _27987_ (.B1(_14373_),
    .Y(_14375_),
    .A1(_13704_),
    .A2(net6494));
 sg13g2_nand2_1 _27988_ (.Y(_14376_),
    .A(_00301_),
    .B(net6497));
 sg13g2_o21ai_1 _27989_ (.B1(_14376_),
    .Y(_14377_),
    .A1(net6155),
    .A2(net6497));
 sg13g2_nand2_1 _27990_ (.Y(_14378_),
    .A(_00300_),
    .B(net6497));
 sg13g2_o21ai_1 _27991_ (.B1(_14378_),
    .Y(_14379_),
    .A1(net6458),
    .A2(net6497));
 sg13g2_nand2_1 _27992_ (.Y(_14380_),
    .A(_00299_),
    .B(net6499));
 sg13g2_o21ai_1 _27993_ (.B1(_14380_),
    .Y(_14381_),
    .A1(net6152),
    .A2(net6499));
 sg13g2_nand2_1 _27994_ (.Y(_14382_),
    .A(_00298_),
    .B(net6498));
 sg13g2_o21ai_1 _27995_ (.B1(_14382_),
    .Y(_14383_),
    .A1(net6151),
    .A2(net6498));
 sg13g2_nand2_1 _27996_ (.Y(_14384_),
    .A(_00297_),
    .B(net6499));
 sg13g2_o21ai_1 _27997_ (.B1(_14384_),
    .Y(_14385_),
    .A1(net6149),
    .A2(net6499));
 sg13g2_nand2_1 _27998_ (.Y(_14386_),
    .A(_00296_),
    .B(net6501));
 sg13g2_o21ai_1 _27999_ (.B1(net7695),
    .Y(_14387_),
    .A1(net7561),
    .A2(_14374_));
 sg13g2_o21ai_1 _28000_ (.B1(_14386_),
    .Y(_14388_),
    .A1(net6148),
    .A2(net6501));
 sg13g2_nand2_1 _28001_ (.Y(_14389_),
    .A(_00295_),
    .B(net6501));
 sg13g2_o21ai_1 _28002_ (.B1(_14389_),
    .Y(_14390_),
    .A1(net6146),
    .A2(net6501));
 sg13g2_nand2_1 _28003_ (.Y(_14391_),
    .A(_00294_),
    .B(net6501));
 sg13g2_o21ai_1 _28004_ (.B1(_14391_),
    .Y(_14392_),
    .A1(_13495_),
    .A2(net6501));
 sg13g2_nand2_1 _28005_ (.Y(_14393_),
    .A(_00293_),
    .B(net6501));
 sg13g2_o21ai_1 _28006_ (.B1(_14393_),
    .Y(_14394_),
    .A1(net6143),
    .A2(net6501));
 sg13g2_nand2_1 _28007_ (.Y(_14395_),
    .A(_00292_),
    .B(net6498));
 sg13g2_or3_1 _28008_ (.A(_14337_),
    .B(_14359_),
    .C(_14387_),
    .X(_14396_));
 sg13g2_o21ai_1 _28009_ (.B1(_14395_),
    .Y(_14397_),
    .A1(_13506_),
    .A2(net6498));
 sg13g2_nand2_1 _28010_ (.Y(_14398_),
    .A(_00291_),
    .B(net6494));
 sg13g2_o21ai_1 _28011_ (.B1(_14398_),
    .Y(_14399_),
    .A1(net6454),
    .A2(net6494));
 sg13g2_nand2_1 _28012_ (.Y(_14400_),
    .A(_00290_),
    .B(net6498));
 sg13g2_o21ai_1 _28013_ (.B1(_14400_),
    .Y(_14401_),
    .A1(net6141),
    .A2(net6498));
 sg13g2_nand2_1 _28014_ (.Y(_14402_),
    .A(_00289_),
    .B(net6497));
 sg13g2_o21ai_1 _28015_ (.B1(_14402_),
    .Y(_14403_),
    .A1(net6139),
    .A2(net6497));
 sg13g2_nand2_1 _28016_ (.Y(_14404_),
    .A(_00288_),
    .B(net6500));
 sg13g2_mux2_1 _28017_ (.A0(_00634_),
    .A1(_00762_),
    .S(net7712),
    .X(_14405_));
 sg13g2_o21ai_1 _28018_ (.B1(_14404_),
    .Y(_14406_),
    .A1(net6138),
    .A2(net6500));
 sg13g2_nand2_1 _28019_ (.Y(_14407_),
    .A(_00287_),
    .B(net6498));
 sg13g2_o21ai_1 _28020_ (.B1(_14407_),
    .Y(_14408_),
    .A1(net6137),
    .A2(net6498));
 sg13g2_nand2_1 _28021_ (.Y(_14409_),
    .A(_00286_),
    .B(net6493));
 sg13g2_o21ai_1 _28022_ (.B1(_14409_),
    .Y(_14410_),
    .A1(_13532_),
    .A2(net6493));
 sg13g2_and2_1 _28023_ (.A(net7774),
    .B(_00928_),
    .X(_14411_));
 sg13g2_nand2_1 _28024_ (.Y(_14412_),
    .A(_00285_),
    .B(net6495));
 sg13g2_o21ai_1 _28025_ (.B1(_14412_),
    .Y(_14413_),
    .A1(net6542),
    .A2(net6495));
 sg13g2_nand2_1 _28026_ (.Y(_14414_),
    .A(_00284_),
    .B(net6496));
 sg13g2_o21ai_1 _28027_ (.B1(_14414_),
    .Y(_14415_),
    .A1(net6135),
    .A2(net6496));
 sg13g2_nand2_1 _28028_ (.Y(_14416_),
    .A(_00283_),
    .B(net6500));
 sg13g2_o21ai_1 _28029_ (.B1(_14416_),
    .Y(_14417_),
    .A1(net6457),
    .A2(net6495));
 sg13g2_nand2_1 _28030_ (.Y(_14418_),
    .A(_00282_),
    .B(net6495));
 sg13g2_nor2b_1 _28031_ (.A(net7774),
    .B_N(_01280_),
    .Y(_14419_));
 sg13g2_o21ai_1 _28032_ (.B1(_14418_),
    .Y(_14420_),
    .A1(net6133),
    .A2(net6495));
 sg13g2_nand2_1 _28033_ (.Y(_14421_),
    .A(_00281_),
    .B(net6495));
 sg13g2_o21ai_1 _28034_ (.B1(_14421_),
    .Y(_14422_),
    .A1(net6455),
    .A2(net6495));
 sg13g2_nand2_1 _28035_ (.Y(_14423_),
    .A(_00280_),
    .B(net6493));
 sg13g2_o21ai_1 _28036_ (.B1(_14423_),
    .Y(_14424_),
    .A1(_13874_),
    .A2(net6493));
 sg13g2_nor4_1 _28037_ (.A(_06923_),
    .B(_06935_),
    .C(_09553_),
    .D(_13422_),
    .Y(_14425_));
 sg13g2_nand2b_1 _28038_ (.Y(_14426_),
    .B(_13568_),
    .A_N(net6591));
 sg13g2_nand2b_1 _28039_ (.Y(_14427_),
    .B(net7276),
    .A_N(_14077_));
 sg13g2_o21ai_1 _28040_ (.B1(_14427_),
    .Y(_14428_),
    .A1(_00279_),
    .A2(net6491));
 sg13g2_a21oi_1 _28041_ (.A1(net6459),
    .A2(net6589),
    .Y(_14429_),
    .B1(_14428_));
 sg13g2_nand2b_1 _28042_ (.Y(_14430_),
    .B(net7276),
    .A_N(_14081_));
 sg13g2_o21ai_1 _28043_ (.B1(_14430_),
    .Y(_14431_),
    .A1(_00278_),
    .A2(net6492));
 sg13g2_a21oi_1 _28044_ (.A1(_13436_),
    .A2(net6590),
    .Y(_14432_),
    .B1(_14431_));
 sg13g2_nand2b_1 _28045_ (.Y(_14433_),
    .B(net7277),
    .A_N(_14087_));
 sg13g2_o21ai_1 _28046_ (.B1(_14433_),
    .Y(_14434_),
    .A1(_00277_),
    .A2(net6491));
 sg13g2_a21oi_1 _28047_ (.A1(net6132),
    .A2(net6589),
    .Y(_14435_),
    .B1(_14434_));
 sg13g2_nand2b_1 _28048_ (.Y(_14436_),
    .B(net7277),
    .A_N(_14092_));
 sg13g2_o21ai_1 _28049_ (.B1(_14436_),
    .Y(_14437_),
    .A1(_00276_),
    .A2(_14426_));
 sg13g2_a21oi_1 _28050_ (.A1(_13621_),
    .A2(net6591),
    .Y(_14438_),
    .B1(_14437_));
 sg13g2_nand2b_1 _28051_ (.Y(_14439_),
    .B(net7277),
    .A_N(_14096_));
 sg13g2_o21ai_1 _28052_ (.B1(_14439_),
    .Y(_14440_),
    .A1(_00275_),
    .A2(net6491));
 sg13g2_a21oi_1 _28053_ (.A1(net6533),
    .A2(net6591),
    .Y(_14441_),
    .B1(_14440_));
 sg13g2_nand2b_1 _28054_ (.Y(_14442_),
    .B(net7280),
    .A_N(_14103_));
 sg13g2_o21ai_1 _28055_ (.B1(_14442_),
    .Y(_14443_),
    .A1(_00274_),
    .A2(_14426_));
 sg13g2_a21oi_1 _28056_ (.A1(_13645_),
    .A2(net6591),
    .Y(_14444_),
    .B1(_14443_));
 sg13g2_mux2_1 _28057_ (.A0(_00666_),
    .A1(_00698_),
    .S(net7774),
    .X(_14445_));
 sg13g2_nand2b_1 _28058_ (.Y(_14446_),
    .B(net7280),
    .A_N(_14116_));
 sg13g2_o21ai_1 _28059_ (.B1(_14446_),
    .Y(_14447_),
    .A1(_00273_),
    .A2(_14426_));
 sg13g2_a21oi_1 _28060_ (.A1(_13656_),
    .A2(net6591),
    .Y(_14448_),
    .B1(_14447_));
 sg13g2_nand2b_1 _28061_ (.Y(_14449_),
    .B(net7276),
    .A_N(_14125_));
 sg13g2_o21ai_1 _28062_ (.B1(_14449_),
    .Y(_14450_),
    .A1(_00272_),
    .A2(net6488));
 sg13g2_a21oi_1 _28063_ (.A1(net6158),
    .A2(net6589),
    .Y(_14451_),
    .B1(_14450_));
 sg13g2_nand2b_1 _28064_ (.Y(_14452_),
    .B(net7278),
    .A_N(_14130_));
 sg13g2_o21ai_1 _28065_ (.B1(_14452_),
    .Y(_14453_),
    .A1(_00271_),
    .A2(net6489));
 sg13g2_nor2b_1 _28066_ (.A(net7774),
    .B_N(_00730_),
    .Y(_14454_));
 sg13g2_a21oi_1 _28067_ (.A1(net6157),
    .A2(net6588),
    .Y(_14455_),
    .B1(_14453_));
 sg13g2_nand2_1 _28068_ (.Y(_14456_),
    .A(net7280),
    .B(_14134_));
 sg13g2_o21ai_1 _28069_ (.B1(_14456_),
    .Y(_14457_),
    .A1(_00270_),
    .A2(_14426_));
 sg13g2_a21oi_1 _28070_ (.A1(_13704_),
    .A2(net6591),
    .Y(_14458_),
    .B1(_14457_));
 sg13g2_nand2b_1 _28071_ (.Y(_14459_),
    .B(net7278),
    .A_N(_14143_));
 sg13g2_o21ai_1 _28072_ (.B1(_14459_),
    .Y(_14460_),
    .A1(_00269_),
    .A2(net6489));
 sg13g2_a21oi_1 _28073_ (.A1(net6154),
    .A2(net6588),
    .Y(_14461_),
    .B1(_14460_));
 sg13g2_nand2b_1 _28074_ (.Y(_14462_),
    .B(net7278),
    .A_N(_14148_));
 sg13g2_o21ai_1 _28075_ (.B1(_14462_),
    .Y(_14463_),
    .A1(_00268_),
    .A2(net6489));
 sg13g2_a21oi_1 _28076_ (.A1(net6458),
    .A2(net6588),
    .Y(_14464_),
    .B1(_14463_));
 sg13g2_nand2b_1 _28077_ (.Y(_14465_),
    .B(net7279),
    .A_N(_14153_));
 sg13g2_o21ai_1 _28078_ (.B1(_14465_),
    .Y(_14466_),
    .A1(_00267_),
    .A2(net6490));
 sg13g2_a21oi_1 _28079_ (.A1(net6153),
    .A2(net6587),
    .Y(_14467_),
    .B1(_14466_));
 sg13g2_nand2b_1 _28080_ (.Y(_14468_),
    .B(net7278),
    .A_N(_14157_));
 sg13g2_o21ai_1 _28081_ (.B1(_14468_),
    .Y(_14469_),
    .A1(_00266_),
    .A2(net6489));
 sg13g2_a21oi_1 _28082_ (.A1(net6150),
    .A2(net6588),
    .Y(_14470_),
    .B1(_14469_));
 sg13g2_nand2b_1 _28083_ (.Y(_14471_),
    .B(net7279),
    .A_N(_14161_));
 sg13g2_o21ai_1 _28084_ (.B1(_14471_),
    .Y(_14472_),
    .A1(_00265_),
    .A2(net6490));
 sg13g2_a21oi_1 _28085_ (.A1(net6149),
    .A2(net6587),
    .Y(_14473_),
    .B1(_14472_));
 sg13g2_nand2b_1 _28086_ (.Y(_14474_),
    .B(net7279),
    .A_N(_14166_));
 sg13g2_o21ai_1 _28087_ (.B1(_14474_),
    .Y(_14475_),
    .A1(_00264_),
    .A2(net6490));
 sg13g2_nor2b_1 _28088_ (.A(_01901_),
    .B_N(net7706),
    .Y(_14476_));
 sg13g2_a21oi_1 _28089_ (.A1(net6147),
    .A2(net6587),
    .Y(_14477_),
    .B1(_14475_));
 sg13g2_nand2b_1 _28090_ (.Y(_14478_),
    .B(net7279),
    .A_N(_14171_));
 sg13g2_o21ai_1 _28091_ (.B1(_14478_),
    .Y(_14479_),
    .A1(_00263_),
    .A2(net6488));
 sg13g2_a21oi_1 _28092_ (.A1(net6145),
    .A2(net6587),
    .Y(_14480_),
    .B1(_14479_));
 sg13g2_nand2b_1 _28093_ (.Y(_14481_),
    .B(net7279),
    .A_N(_14175_));
 sg13g2_o21ai_1 _28094_ (.B1(_14481_),
    .Y(_14482_),
    .A1(_00262_),
    .A2(net6488));
 sg13g2_a21oi_1 _28095_ (.A1(net6144),
    .A2(net6587),
    .Y(_14483_),
    .B1(_14482_));
 sg13g2_nand2b_1 _28096_ (.Y(_14484_),
    .B(net7277),
    .A_N(_14179_));
 sg13g2_o21ai_1 _28097_ (.B1(_14484_),
    .Y(_14485_),
    .A1(_00261_),
    .A2(net6488));
 sg13g2_a21oi_1 _28098_ (.A1(net6143),
    .A2(net6589),
    .Y(_14486_),
    .B1(_14485_));
 sg13g2_nand2b_1 _28099_ (.Y(_14487_),
    .B(net7277),
    .A_N(_14184_));
 sg13g2_o21ai_1 _28100_ (.B1(_14487_),
    .Y(_14488_),
    .A1(_00260_),
    .A2(net6491));
 sg13g2_a21oi_1 _28101_ (.A1(_13506_),
    .A2(net6589),
    .Y(_14489_),
    .B1(_14488_));
 sg13g2_nand2b_1 _28102_ (.Y(_14490_),
    .B(net7276),
    .A_N(_14191_));
 sg13g2_o21ai_1 _28103_ (.B1(_14490_),
    .Y(_14491_),
    .A1(_00259_),
    .A2(_14426_));
 sg13g2_a21oi_1 _28104_ (.A1(_13779_),
    .A2(net6590),
    .Y(_14492_),
    .B1(_14491_));
 sg13g2_nand2b_1 _28105_ (.Y(_14493_),
    .B(net7278),
    .A_N(_14198_));
 sg13g2_o21ai_1 _28106_ (.B1(_14493_),
    .Y(_14494_),
    .A1(_00258_),
    .A2(net6489));
 sg13g2_a21oi_1 _28107_ (.A1(net6141),
    .A2(net6588),
    .Y(_14495_),
    .B1(_14494_));
 sg13g2_nand2b_1 _28108_ (.Y(_14496_),
    .B(net7278),
    .A_N(_14205_));
 sg13g2_o21ai_1 _28109_ (.B1(_14496_),
    .Y(_14497_),
    .A1(_00257_),
    .A2(net6489));
 sg13g2_a21oi_1 _28110_ (.A1(net6140),
    .A2(net6588),
    .Y(_14498_),
    .B1(_14497_));
 sg13g2_nand2b_1 _28111_ (.Y(_14499_),
    .B(net7278),
    .A_N(_14209_));
 sg13g2_o21ai_1 _28112_ (.B1(_14499_),
    .Y(_14500_),
    .A1(_00256_),
    .A2(net6489));
 sg13g2_a21oi_1 _28113_ (.A1(net6138),
    .A2(net6588),
    .Y(_14501_),
    .B1(_14500_));
 sg13g2_nand2b_1 _28114_ (.Y(_14502_),
    .B(net7277),
    .A_N(_14213_));
 sg13g2_o21ai_1 _28115_ (.B1(_14502_),
    .Y(_14503_),
    .A1(_00255_),
    .A2(net6488));
 sg13g2_a21oi_1 _28116_ (.A1(_13527_),
    .A2(net6587),
    .Y(_14504_),
    .B1(_14503_));
 sg13g2_mux4_1 _28117_ (.S0(net7744),
    .A0(_14411_),
    .A1(_14419_),
    .A2(_14445_),
    .A3(_14454_),
    .S1(net7712),
    .X(_14505_));
 sg13g2_nand2b_1 _28118_ (.Y(_14506_),
    .B(net7277),
    .A_N(_14217_));
 sg13g2_o21ai_1 _28119_ (.B1(_14506_),
    .Y(_14507_),
    .A1(_00254_),
    .A2(net6491));
 sg13g2_a21oi_1 _28120_ (.A1(net6543),
    .A2(net6589),
    .Y(_14508_),
    .B1(_14507_));
 sg13g2_nand2b_1 _28121_ (.Y(_14509_),
    .B(net7276),
    .A_N(_14221_));
 sg13g2_o21ai_1 _28122_ (.B1(_14509_),
    .Y(_14510_),
    .A1(_00253_),
    .A2(net6492));
 sg13g2_a221oi_1 _28123_ (.B2(net7533),
    .C1(net7690),
    .B1(_14505_),
    .A1(net7435),
    .Y(_14511_),
    .A2(_14405_));
 sg13g2_a21oi_1 _28124_ (.A1(net6542),
    .A2(net6590),
    .Y(_14512_),
    .B1(_14510_));
 sg13g2_nand2b_1 _28125_ (.Y(_14513_),
    .B(net7276),
    .A_N(_14225_));
 sg13g2_o21ai_1 _28126_ (.B1(_14513_),
    .Y(_14514_),
    .A1(_00252_),
    .A2(net6492));
 sg13g2_a21oi_1 _28127_ (.A1(net6136),
    .A2(net6590),
    .Y(_14515_),
    .B1(_14514_));
 sg13g2_nand2b_1 _28128_ (.Y(_14516_),
    .B(net7276),
    .A_N(_14230_));
 sg13g2_o21ai_1 _28129_ (.B1(_14516_),
    .Y(_14517_),
    .A1(_00251_),
    .A2(net6492));
 sg13g2_a21oi_1 _28130_ (.A1(net6456),
    .A2(net6590),
    .Y(_14518_),
    .B1(_14517_));
 sg13g2_nand2b_1 _28131_ (.Y(_14519_),
    .B(net7277),
    .A_N(_14234_));
 sg13g2_o21ai_1 _28132_ (.B1(_14519_),
    .Y(_14520_),
    .A1(_00250_),
    .A2(net6488));
 sg13g2_a21oi_1 _28133_ (.A1(net6134),
    .A2(net6587),
    .Y(_14521_),
    .B1(_14520_));
 sg13g2_nand2b_1 _28134_ (.Y(_14522_),
    .B(net7276),
    .A_N(_14239_));
 sg13g2_o21ai_1 _28135_ (.B1(_14522_),
    .Y(_14523_),
    .A1(_00249_),
    .A2(net6492));
 sg13g2_a21oi_1 _28136_ (.A1(net6455),
    .A2(net6590),
    .Y(_14524_),
    .B1(_14523_));
 sg13g2_nand2_1 _28137_ (.Y(_14525_),
    .A(_01600_),
    .B(\cs_registers_i.debug_single_step_o ));
 sg13g2_o21ai_1 _28138_ (.B1(_14525_),
    .Y(_14526_),
    .A1(_06135_),
    .A2(net7279));
 sg13g2_nand2_1 _28139_ (.Y(_14527_),
    .A(_00247_),
    .B(_13568_));
 sg13g2_nand2_1 _28140_ (.Y(_14528_),
    .A(net349),
    .B(_01600_));
 sg13g2_o21ai_1 _28141_ (.B1(_14527_),
    .Y(_14529_),
    .A1(\cs_registers_i.debug_single_step_o ),
    .A2(_14528_));
 sg13g2_a22oi_1 _28142_ (.Y(_14530_),
    .B1(_13568_),
    .B2(_06140_),
    .A2(\cs_registers_i.debug_single_step_o ),
    .A1(_01600_));
 sg13g2_nand2_1 _28143_ (.Y(_14531_),
    .A(net6673),
    .B(net6592));
 sg13g2_nand2_1 _28144_ (.Y(_14532_),
    .A(\cs_registers_i.debug_single_step_o ),
    .B(net6487));
 sg13g2_o21ai_1 _28145_ (.B1(_14532_),
    .Y(_14533_),
    .A1(_13704_),
    .A2(net6487));
 sg13g2_a21oi_1 _28146_ (.A1(_09661_),
    .A2(net6592),
    .Y(_14534_),
    .B1(net7279));
 sg13g2_a22oi_1 _28147_ (.Y(_14535_),
    .B1(_14534_),
    .B2(_00001_),
    .A2(net7280),
    .A1(_00243_));
 sg13g2_nand2_1 _28148_ (.Y(_14536_),
    .A(net6454),
    .B(_13874_));
 sg13g2_o21ai_1 _28149_ (.B1(_14535_),
    .Y(_14537_),
    .A1(net6487),
    .A2(_14536_));
 sg13g2_nand2_1 _28150_ (.Y(_14538_),
    .A(\cs_registers_i.debug_ebreakm_o ),
    .B(net6487));
 sg13g2_o21ai_1 _28151_ (.B1(_14538_),
    .Y(_14539_),
    .A1(_13532_),
    .A2(net6487));
 sg13g2_mux2_1 _28152_ (.A0(_01421_),
    .A1(_01457_),
    .S(net7768),
    .X(_14540_));
 sg13g2_nand2_1 _28153_ (.Y(_14541_),
    .A(_00245_),
    .B(_14531_));
 sg13g2_o21ai_1 _28154_ (.B1(_14541_),
    .Y(_14542_),
    .A1(net6135),
    .A2(_14531_));
 sg13g2_nor3_1 _28155_ (.A(net7577),
    .B(net7569),
    .C(_14540_),
    .Y(_14543_));
 sg13g2_nand2_1 _28156_ (.Y(_14544_),
    .A(\cs_registers_i.debug_ebreaku_o ),
    .B(net6487));
 sg13g2_o21ai_1 _28157_ (.B1(_14544_),
    .Y(_14545_),
    .A1(net6457),
    .A2(net6487));
 sg13g2_nand2_1 _28158_ (.Y(_14546_),
    .A(_00244_),
    .B(_14531_));
 sg13g2_o21ai_1 _28159_ (.B1(_14546_),
    .Y(_14547_),
    .A1(net6133),
    .A2(_14531_));
 sg13g2_a22oi_1 _28160_ (.Y(_14548_),
    .B1(_14534_),
    .B2(_00000_),
    .A2(net7280),
    .A1(_00242_));
 sg13g2_o21ai_1 _28161_ (.B1(_14548_),
    .Y(_14549_),
    .A1(net6487),
    .A2(_14536_));
 sg13g2_a22oi_1 _28162_ (.Y(_14550_),
    .B1(net7313),
    .B2(_00474_),
    .A2(net7105),
    .A1(_06145_));
 sg13g2_nor2_1 _28163_ (.A(_07692_),
    .B(_14550_),
    .Y(_14551_));
 sg13g2_a21oi_1 _28164_ (.A1(_06965_),
    .A2(_07691_),
    .Y(_14552_),
    .B1(_00243_));
 sg13g2_nor3_1 _28165_ (.A(_13566_),
    .B(_14551_),
    .C(_14552_),
    .Y(_14553_));
 sg13g2_a22oi_1 _28166_ (.Y(_14554_),
    .B1(net7313),
    .B2(_00473_),
    .A2(net7105),
    .A1(_06149_));
 sg13g2_nor2_1 _28167_ (.A(_07692_),
    .B(_14554_),
    .Y(_14555_));
 sg13g2_a21oi_1 _28168_ (.A1(_06965_),
    .A2(_07691_),
    .Y(_14556_),
    .B1(_00242_));
 sg13g2_nor3_1 _28169_ (.A(_13566_),
    .B(_14555_),
    .C(_14556_),
    .Y(_14557_));
 sg13g2_nand2_1 _28170_ (.Y(_14558_),
    .A(net6950),
    .B(net6930));
 sg13g2_nand2_1 _28171_ (.Y(_14559_),
    .A(net6592),
    .B(_14558_));
 sg13g2_nand3_1 _28172_ (.B(_03638_),
    .C(_06626_),
    .A(net7607),
    .Y(_14560_));
 sg13g2_nor3_1 _28173_ (.A(\id_stage_i.controller_i.instr_fetch_err_i ),
    .B(_00113_),
    .C(_06963_),
    .Y(_14561_));
 sg13g2_and4_1 _28174_ (.A(_06767_),
    .B(_06911_),
    .C(_14560_),
    .D(_14561_),
    .X(_14562_));
 sg13g2_mux2_1 _28175_ (.A0(_01492_),
    .A1(_01527_),
    .S(net7787),
    .X(_14563_));
 sg13g2_nand3_1 _28176_ (.B(_09330_),
    .C(_14562_),
    .A(_07041_),
    .Y(_14564_));
 sg13g2_nand2_1 _28177_ (.Y(_14565_),
    .A(_13423_),
    .B(_14558_));
 sg13g2_nand4_1 _28178_ (.B(_06957_),
    .C(_13426_),
    .A(_06894_),
    .Y(_14566_),
    .D(_14558_));
 sg13g2_nor2_1 _28179_ (.A(net6794),
    .B(_14566_),
    .Y(_14567_));
 sg13g2_nor3_1 _28180_ (.A(net7577),
    .B(net7561),
    .C(_14563_),
    .Y(_14568_));
 sg13g2_nand2_1 _28181_ (.Y(_14569_),
    .A(net6709),
    .B(_14567_));
 sg13g2_nor3_2 _28182_ (.A(_06921_),
    .B(net6794),
    .C(_14565_),
    .Y(_14570_));
 sg13g2_or3_1 _28183_ (.A(_06921_),
    .B(net6794),
    .C(_14565_),
    .X(_14571_));
 sg13g2_a22oi_1 _28184_ (.Y(_14572_),
    .B1(_14570_),
    .B2(_06920_),
    .A2(_14569_),
    .A1(net5881));
 sg13g2_and3_1 _28185_ (.X(_14573_),
    .A(_00200_),
    .B(_00189_),
    .C(_00178_));
 sg13g2_and2_1 _28186_ (.A(_00211_),
    .B(_14573_),
    .X(_14574_));
 sg13g2_nand2_1 _28187_ (.Y(_14575_),
    .A(_00222_),
    .B(_14574_));
 sg13g2_and3_1 _28188_ (.X(_14576_),
    .A(_00233_),
    .B(_00222_),
    .C(_14574_));
 sg13g2_nand2_1 _28189_ (.Y(_14577_),
    .A(_00238_),
    .B(_14576_));
 sg13g2_and3_1 _28190_ (.X(_14578_),
    .A(_00239_),
    .B(_00238_),
    .C(_14576_));
 sg13g2_and2_1 _28191_ (.A(_00240_),
    .B(_14578_),
    .X(_14579_));
 sg13g2_nand2_1 _28192_ (.Y(_14580_),
    .A(_00240_),
    .B(_14578_));
 sg13g2_nor3_1 _28193_ (.A(_06866_),
    .B(net6794),
    .C(_14559_),
    .Y(_14581_));
 sg13g2_and2_1 _28194_ (.A(_06941_),
    .B(_14567_),
    .X(_14582_));
 sg13g2_o21ai_1 _28195_ (.B1(net5826),
    .Y(_14583_),
    .A1(net6443),
    .A2(_14579_));
 sg13g2_nand2_1 _28196_ (.Y(_14584_),
    .A(_00241_),
    .B(_14579_));
 sg13g2_nand2_1 _28197_ (.Y(_14585_),
    .A(_13431_),
    .B(net6444));
 sg13g2_o21ai_1 _28198_ (.B1(_14585_),
    .Y(_14586_),
    .A1(net6443),
    .A2(_14584_));
 sg13g2_a22oi_1 _28199_ (.Y(_14587_),
    .B1(_14586_),
    .B2(net5826),
    .A2(_14583_),
    .A1(_06168_));
 sg13g2_nand2_1 _28200_ (.Y(_14588_),
    .A(net6159),
    .B(net6441));
 sg13g2_o21ai_1 _28201_ (.B1(_14588_),
    .Y(_14589_),
    .A1(_14580_),
    .A2(_14581_));
 sg13g2_o21ai_1 _28202_ (.B1(net5823),
    .Y(_14590_),
    .A1(net6441),
    .A2(_14578_));
 sg13g2_a22oi_1 _28203_ (.Y(_14591_),
    .B1(_14590_),
    .B2(_06174_),
    .A2(_14589_),
    .A1(net5823));
 sg13g2_nand2_1 _28204_ (.Y(_14592_),
    .A(net6438),
    .B(_14578_));
 sg13g2_nand2_1 _28205_ (.Y(_14593_),
    .A(_13610_),
    .B(net6441));
 sg13g2_mux2_1 _28206_ (.A0(_01351_),
    .A1(_01386_),
    .S(net7768),
    .X(_14594_));
 sg13g2_nand2_1 _28207_ (.Y(_14595_),
    .A(_14592_),
    .B(_14593_));
 sg13g2_nand2_1 _28208_ (.Y(_14596_),
    .A(net6439),
    .B(_14577_));
 sg13g2_a21oi_1 _28209_ (.A1(net5823),
    .A2(_14596_),
    .Y(_14597_),
    .B1(_00239_));
 sg13g2_a21oi_1 _28210_ (.A1(net5823),
    .A2(_14595_),
    .Y(_14598_),
    .B1(_14597_));
 sg13g2_o21ai_1 _28211_ (.B1(net6930),
    .Y(_14599_),
    .A1(net6950),
    .A2(_06893_));
 sg13g2_nor3_1 _28212_ (.A(net7577),
    .B(_08503_),
    .C(_14594_),
    .Y(_14600_));
 sg13g2_and3_1 _28213_ (.X(_14601_),
    .A(_06941_),
    .B(_13426_),
    .C(_14599_));
 sg13g2_nor2b_1 _28214_ (.A(net6794),
    .B_N(_14601_),
    .Y(_14602_));
 sg13g2_nand2_1 _28215_ (.Y(_14603_),
    .A(_13621_),
    .B(net6441));
 sg13g2_o21ai_1 _28216_ (.B1(_14603_),
    .Y(_14604_),
    .A1(_14577_),
    .A2(_14602_));
 sg13g2_o21ai_1 _28217_ (.B1(net5823),
    .Y(_14605_),
    .A1(net6441),
    .A2(_14576_));
 sg13g2_a22oi_1 _28218_ (.Y(_14606_),
    .B1(_14605_),
    .B2(_06185_),
    .A2(_14604_),
    .A1(net5823));
 sg13g2_or2_1 _28219_ (.X(_14607_),
    .B(_14582_),
    .A(net5881));
 sg13g2_nand2_1 _28220_ (.Y(_14608_),
    .A(net6707),
    .B(_14567_));
 sg13g2_nand2_1 _28221_ (.Y(_14609_),
    .A(_14607_),
    .B(_14608_));
 sg13g2_and4_1 _28222_ (.A(_00192_),
    .B(_00191_),
    .C(_00190_),
    .D(_00188_),
    .X(_14610_));
 sg13g2_nand4_1 _28223_ (.B(_00194_),
    .C(_00193_),
    .A(_00195_),
    .Y(_14611_),
    .D(_14610_));
 sg13g2_nand2_1 _28224_ (.Y(_14612_),
    .A(_00204_),
    .B(_00203_));
 sg13g2_mux2_1 _28225_ (.A0(_01562_),
    .A1(_01597_),
    .S(net7768),
    .X(_14613_));
 sg13g2_and3_1 _28226_ (.X(_14614_),
    .A(_00205_),
    .B(_00204_),
    .C(_00203_));
 sg13g2_nand3_1 _28227_ (.B(_00204_),
    .C(_00203_),
    .A(_00205_),
    .Y(_14615_));
 sg13g2_nand3_1 _28228_ (.B(_00206_),
    .C(_14614_),
    .A(_00207_),
    .Y(_14616_));
 sg13g2_or2_1 _28229_ (.X(_14617_),
    .B(_14616_),
    .A(_06266_));
 sg13g2_nor2_1 _28230_ (.A(net7556),
    .B(_14613_),
    .Y(_14618_));
 sg13g2_and2_1 _28231_ (.A(_00201_),
    .B(_00199_),
    .X(_14619_));
 sg13g2_nand4_1 _28232_ (.B(_00198_),
    .C(_00197_),
    .A(_00202_),
    .Y(_14620_),
    .D(_14619_));
 sg13g2_nand3_1 _28233_ (.B(_00215_),
    .C(_00214_),
    .A(_00216_),
    .Y(_14621_));
 sg13g2_or4_1 _28234_ (.A(_14543_),
    .B(_14568_),
    .C(_14600_),
    .D(_14618_),
    .X(_14622_));
 sg13g2_nand4_1 _28235_ (.B(_00181_),
    .C(_00180_),
    .A(_00182_),
    .Y(_14623_),
    .D(_00179_));
 sg13g2_nor3_1 _28236_ (.A(_06168_),
    .B(_14580_),
    .C(_14623_),
    .Y(_14624_));
 sg13g2_and2_1 _28237_ (.A(_00183_),
    .B(_14624_),
    .X(_14625_));
 sg13g2_inv_1 _28238_ (.Y(_14626_),
    .A(_14625_));
 sg13g2_and2_1 _28239_ (.A(_00184_),
    .B(_14625_),
    .X(_14627_));
 sg13g2_nand2_1 _28240_ (.Y(_14628_),
    .A(_00184_),
    .B(_14625_));
 sg13g2_nand4_1 _28241_ (.B(_00187_),
    .C(_00186_),
    .A(_00196_),
    .Y(_14629_),
    .D(_00185_));
 sg13g2_inv_1 _28242_ (.Y(_14630_),
    .A(_14631_));
 sg13g2_or3_1 _28243_ (.A(_14611_),
    .B(_14628_),
    .C(_14629_),
    .X(_14631_));
 sg13g2_nand3_1 _28244_ (.B(_00210_),
    .C(_00209_),
    .A(_00212_),
    .Y(_14632_));
 sg13g2_nor4_1 _28245_ (.A(_14617_),
    .B(_14620_),
    .C(_14631_),
    .D(_14632_),
    .Y(_14633_));
 sg13g2_inv_1 _28246_ (.Y(_14634_),
    .A(_14633_));
 sg13g2_nand3_1 _28247_ (.B(_00217_),
    .C(_00213_),
    .A(_00218_),
    .Y(_14635_));
 sg13g2_nor3_1 _28248_ (.A(_14621_),
    .B(_14634_),
    .C(_14635_),
    .Y(_14636_));
 sg13g2_and2_1 _28249_ (.A(_00219_),
    .B(_14636_),
    .X(_14637_));
 sg13g2_nand2_1 _28250_ (.Y(_14638_),
    .A(_00219_),
    .B(_14636_));
 sg13g2_nor2_1 _28251_ (.A(_06240_),
    .B(_14638_),
    .Y(_14639_));
 sg13g2_nand2_1 _28252_ (.Y(_14640_),
    .A(_00220_),
    .B(_14637_));
 sg13g2_nor2_1 _28253_ (.A(_06239_),
    .B(_14640_),
    .Y(_14641_));
 sg13g2_nand2_1 _28254_ (.Y(_14642_),
    .A(_00221_),
    .B(_14639_));
 sg13g2_nor2_1 _28255_ (.A(_06235_),
    .B(_14642_),
    .Y(_14643_));
 sg13g2_nand2_1 _28256_ (.Y(_14644_),
    .A(_00223_),
    .B(_14641_));
 sg13g2_nor2_1 _28257_ (.A(_06231_),
    .B(_14644_),
    .Y(_14645_));
 sg13g2_nand2_1 _28258_ (.Y(_14646_),
    .A(_00224_),
    .B(_14643_));
 sg13g2_nor2_1 _28259_ (.A(_06227_),
    .B(_14646_),
    .Y(_14647_));
 sg13g2_nand2_1 _28260_ (.Y(_14648_),
    .A(_00225_),
    .B(_14645_));
 sg13g2_nand2_1 _28261_ (.Y(_14649_),
    .A(_00226_),
    .B(_14647_));
 sg13g2_and3_1 _28262_ (.X(_14650_),
    .A(_00227_),
    .B(_00226_),
    .C(_14647_));
 sg13g2_inv_1 _28263_ (.Y(_14651_),
    .A(_14650_));
 sg13g2_and4_1 _28264_ (.A(_00230_),
    .B(_00229_),
    .C(_00228_),
    .D(_14650_),
    .X(_14652_));
 sg13g2_and2_1 _28265_ (.A(_00231_),
    .B(_14652_),
    .X(_14653_));
 sg13g2_nand2_1 _28266_ (.Y(_14654_),
    .A(_00231_),
    .B(_14652_));
 sg13g2_nor2_1 _28267_ (.A(_06208_),
    .B(_14654_),
    .Y(_14655_));
 sg13g2_nand2_1 _28268_ (.Y(_14656_),
    .A(_00232_),
    .B(_14653_));
 sg13g2_mux2_1 _28269_ (.A0(_01140_),
    .A1(_01175_),
    .S(net7771),
    .X(_14657_));
 sg13g2_nor2_1 _28270_ (.A(_06199_),
    .B(_14656_),
    .Y(_14658_));
 sg13g2_nand2_1 _28271_ (.Y(_14659_),
    .A(_00234_),
    .B(_14655_));
 sg13g2_nand2_1 _28272_ (.Y(_14660_),
    .A(_00235_),
    .B(_14658_));
 sg13g2_nand3_1 _28273_ (.B(_00235_),
    .C(_14658_),
    .A(_00236_),
    .Y(_14661_));
 sg13g2_nand2_1 _28274_ (.Y(_14662_),
    .A(net6435),
    .B(_14661_));
 sg13g2_a21oi_1 _28275_ (.A1(net5770),
    .A2(_14662_),
    .Y(_14663_),
    .B1(_00237_));
 sg13g2_nor2_1 _28276_ (.A(net6453),
    .B(_14661_),
    .Y(_14664_));
 sg13g2_a22oi_1 _28277_ (.Y(_14665_),
    .B1(_14664_),
    .B2(_00237_),
    .A2(net6453),
    .A1(_13441_));
 sg13g2_inv_1 _28278_ (.Y(_14666_),
    .A(_14665_));
 sg13g2_a21oi_1 _28279_ (.A1(net5770),
    .A2(_14666_),
    .Y(_14667_),
    .B1(_14663_));
 sg13g2_nand2_1 _28280_ (.Y(_14668_),
    .A(net6435),
    .B(_14660_));
 sg13g2_a21oi_1 _28281_ (.A1(net5770),
    .A2(_14668_),
    .Y(_14669_),
    .B1(_00236_));
 sg13g2_nand2_1 _28282_ (.Y(_14670_),
    .A(_13446_),
    .B(net6447));
 sg13g2_o21ai_1 _28283_ (.B1(_14670_),
    .Y(_14671_),
    .A1(net6447),
    .A2(_14661_));
 sg13g2_a21oi_1 _28284_ (.A1(net5770),
    .A2(_14671_),
    .Y(_14672_),
    .B1(_14669_));
 sg13g2_o21ai_1 _28285_ (.B1(net5770),
    .Y(_14673_),
    .A1(net6434),
    .A2(_14658_));
 sg13g2_nand2_1 _28286_ (.Y(_14674_),
    .A(net6155),
    .B(net6447));
 sg13g2_o21ai_1 _28287_ (.B1(_14674_),
    .Y(_14675_),
    .A1(net6447),
    .A2(_14660_));
 sg13g2_a22oi_1 _28288_ (.Y(_14676_),
    .B1(_14675_),
    .B2(net5770),
    .A2(_14673_),
    .A1(_06195_));
 sg13g2_mux2_1 _28289_ (.A0(_01069_),
    .A1(_01105_),
    .S(net7771),
    .X(_14677_));
 sg13g2_o21ai_1 _28290_ (.B1(net5770),
    .Y(_14678_),
    .A1(net6434),
    .A2(_14655_));
 sg13g2_nand2_1 _28291_ (.Y(_14679_),
    .A(_13458_),
    .B(net6448));
 sg13g2_o21ai_1 _28292_ (.B1(_14679_),
    .Y(_14680_),
    .A1(net6448),
    .A2(_14659_));
 sg13g2_a22oi_1 _28293_ (.Y(_14681_),
    .B1(_14680_),
    .B2(net5770),
    .A2(_14678_),
    .A1(_06199_));
 sg13g2_mux2_1 _28294_ (.A0(_14576_),
    .A1(_13634_),
    .S(net6433),
    .X(_14682_));
 sg13g2_nand2_1 _28295_ (.Y(_14683_),
    .A(net6437),
    .B(_14575_));
 sg13g2_a21oi_1 _28296_ (.A1(net5827),
    .A2(_14683_),
    .Y(_14684_),
    .B1(_00233_));
 sg13g2_a21oi_1 _28297_ (.A1(net5823),
    .A2(_14682_),
    .Y(_14685_),
    .B1(_14684_));
 sg13g2_o21ai_1 _28298_ (.B1(net5769),
    .Y(_14686_),
    .A1(net6434),
    .A2(_14653_));
 sg13g2_nand2_1 _28299_ (.Y(_14687_),
    .A(net6152),
    .B(net6448));
 sg13g2_o21ai_1 _28300_ (.B1(_14687_),
    .Y(_14688_),
    .A1(net6448),
    .A2(_14656_));
 sg13g2_a22oi_1 _28301_ (.Y(_14689_),
    .B1(_14688_),
    .B2(net5769),
    .A2(_14686_),
    .A1(_06208_));
 sg13g2_mux2_1 _28302_ (.A0(_01281_),
    .A1(_01316_),
    .S(net7769),
    .X(_14690_));
 sg13g2_o21ai_1 _28303_ (.B1(net5769),
    .Y(_14691_),
    .A1(net6434),
    .A2(_14652_));
 sg13g2_nand2_1 _28304_ (.Y(_14692_),
    .A(_13471_),
    .B(net6450));
 sg13g2_o21ai_1 _28305_ (.B1(_14692_),
    .Y(_14693_),
    .A1(net6449),
    .A2(_14654_));
 sg13g2_a22oi_1 _28306_ (.Y(_14694_),
    .B1(_14693_),
    .B2(net5769),
    .A2(_14691_),
    .A1(_06210_));
 sg13g2_nand2_1 _28307_ (.Y(_14695_),
    .A(_00228_),
    .B(_14650_));
 sg13g2_nand3_1 _28308_ (.B(_00228_),
    .C(_14650_),
    .A(_00229_),
    .Y(_14696_));
 sg13g2_nand2_1 _28309_ (.Y(_14697_),
    .A(net6435),
    .B(_14696_));
 sg13g2_a21oi_1 _28310_ (.A1(net5768),
    .A2(_14697_),
    .Y(_14698_),
    .B1(_00230_));
 sg13g2_nand4_1 _28311_ (.B(_00229_),
    .C(_00228_),
    .A(_00230_),
    .Y(_14699_),
    .D(_14650_));
 sg13g2_nand2_1 _28312_ (.Y(_14700_),
    .A(_13477_),
    .B(net6451));
 sg13g2_o21ai_1 _28313_ (.B1(_14700_),
    .Y(_14701_),
    .A1(net6451),
    .A2(_14699_));
 sg13g2_a21oi_1 _28314_ (.A1(net5768),
    .A2(_14701_),
    .Y(_14702_),
    .B1(_14698_));
 sg13g2_nand2_1 _28315_ (.Y(_14703_),
    .A(net6435),
    .B(_14695_));
 sg13g2_a21oi_1 _28316_ (.A1(net5768),
    .A2(_14703_),
    .Y(_14704_),
    .B1(_00229_));
 sg13g2_nand2_1 _28317_ (.Y(_14705_),
    .A(_13484_),
    .B(net6451));
 sg13g2_o21ai_1 _28318_ (.B1(_14705_),
    .Y(_14706_),
    .A1(net6451),
    .A2(_14696_));
 sg13g2_a21oi_1 _28319_ (.A1(net5768),
    .A2(_14706_),
    .Y(_14707_),
    .B1(_14704_));
 sg13g2_mux2_1 _28320_ (.A0(_01210_),
    .A1(_01245_),
    .S(net7769),
    .X(_14708_));
 sg13g2_o21ai_1 _28321_ (.B1(net5767),
    .Y(_14709_),
    .A1(net6434),
    .A2(_14650_));
 sg13g2_nand2_1 _28322_ (.Y(_14710_),
    .A(net6146),
    .B(net6452));
 sg13g2_o21ai_1 _28323_ (.B1(_14710_),
    .Y(_14711_),
    .A1(net6452),
    .A2(_14695_));
 sg13g2_a22oi_1 _28324_ (.Y(_14712_),
    .B1(_14711_),
    .B2(net5768),
    .A2(_14709_),
    .A1(_06219_));
 sg13g2_nand2_1 _28325_ (.Y(_14713_),
    .A(net6436),
    .B(_14649_));
 sg13g2_mux4_1 _28326_ (.S0(net7518),
    .A0(_14657_),
    .A1(_14677_),
    .A2(_14690_),
    .A3(_14708_),
    .S1(net7713),
    .X(_14714_));
 sg13g2_a21oi_1 _28327_ (.A1(net5767),
    .A2(_14713_),
    .Y(_14715_),
    .B1(_00227_));
 sg13g2_inv_1 _28328_ (.Y(_14716_),
    .A(_14714_));
 sg13g2_nand2_1 _28329_ (.Y(_14717_),
    .A(_13495_),
    .B(net6449));
 sg13g2_o21ai_1 _28330_ (.B1(_14717_),
    .Y(_14718_),
    .A1(net6449),
    .A2(_14651_));
 sg13g2_a21oi_1 _28331_ (.A1(net5767),
    .A2(_14718_),
    .Y(_14719_),
    .B1(_14715_));
 sg13g2_a21o_1 _28332_ (.A2(_14716_),
    .A1(_08384_),
    .B1(_14622_),
    .X(_14720_));
 sg13g2_o21ai_1 _28333_ (.B1(net5767),
    .Y(_14721_),
    .A1(net6434),
    .A2(_14647_));
 sg13g2_a221oi_1 _28334_ (.B2(_08384_),
    .C1(_14622_),
    .B1(_14716_),
    .A1(_14396_),
    .Y(_14722_),
    .A2(_14511_));
 sg13g2_nand2_1 _28335_ (.Y(_14723_),
    .A(_13501_),
    .B(net6449));
 sg13g2_o21ai_1 _28336_ (.B1(_14723_),
    .Y(_14724_),
    .A1(net6449),
    .A2(_14649_));
 sg13g2_a21o_1 _28337_ (.A2(_14511_),
    .A1(_14396_),
    .B1(_14720_),
    .X(_14725_));
 sg13g2_a22oi_1 _28338_ (.Y(_14726_),
    .B1(_14724_),
    .B2(net5767),
    .A2(_14721_),
    .A1(_06224_));
 sg13g2_o21ai_1 _28339_ (.B1(net5767),
    .Y(_14727_),
    .A1(net6434),
    .A2(_14645_));
 sg13g2_nand2_1 _28340_ (.Y(_14728_),
    .A(net7683),
    .B(_13410_));
 sg13g2_nand2_1 _28341_ (.Y(_14729_),
    .A(net6142),
    .B(net6449));
 sg13g2_o21ai_1 _28342_ (.B1(_14729_),
    .Y(_14730_),
    .A1(net6449),
    .A2(_14648_));
 sg13g2_a22oi_1 _28343_ (.Y(_14731_),
    .B1(_14730_),
    .B2(net5767),
    .A2(_14727_),
    .A1(_06227_));
 sg13g2_o21ai_1 _28344_ (.B1(net5771),
    .Y(_14732_),
    .A1(net6432),
    .A2(_14643_));
 sg13g2_nand2_1 _28345_ (.Y(_14733_),
    .A(_13511_),
    .B(net6446));
 sg13g2_o21ai_1 _28346_ (.B1(_14733_),
    .Y(_14734_),
    .A1(net6446),
    .A2(_14646_));
 sg13g2_a22oi_1 _28347_ (.Y(_14735_),
    .B1(_14734_),
    .B2(net5767),
    .A2(_14732_),
    .A1(_06231_));
 sg13g2_o21ai_1 _28348_ (.B1(net5766),
    .Y(_14736_),
    .A1(net6432),
    .A2(_14641_));
 sg13g2_nand2_1 _28349_ (.Y(_14737_),
    .A(net6140),
    .B(net6446));
 sg13g2_o21ai_1 _28350_ (.B1(_14737_),
    .Y(_14738_),
    .A1(net6445),
    .A2(_14644_));
 sg13g2_a22oi_1 _28351_ (.Y(_14739_),
    .B1(_14738_),
    .B2(net5766),
    .A2(_14736_),
    .A1(_06235_));
 sg13g2_nand2_1 _28352_ (.Y(_14740_),
    .A(_13645_),
    .B(net6441));
 sg13g2_o21ai_1 _28353_ (.B1(_14740_),
    .Y(_14741_),
    .A1(_14575_),
    .A2(_14581_));
 sg13g2_o21ai_1 _28354_ (.B1(net5823),
    .Y(_14742_),
    .A1(net6441),
    .A2(_14574_));
 sg13g2_a22oi_1 _28355_ (.Y(_14743_),
    .B1(_14742_),
    .B2(_06236_),
    .A2(_14741_),
    .A1(net5821));
 sg13g2_o21ai_1 _28356_ (.B1(net5766),
    .Y(_14744_),
    .A1(net6432),
    .A2(_14639_));
 sg13g2_nand2_1 _28357_ (.Y(_14745_),
    .A(_13522_),
    .B(net6445));
 sg13g2_o21ai_1 _28358_ (.B1(_14745_),
    .Y(_14746_),
    .A1(net6445),
    .A2(_14642_));
 sg13g2_a22oi_1 _28359_ (.Y(_14747_),
    .B1(_14746_),
    .B2(net5766),
    .A2(_14744_),
    .A1(_06239_));
 sg13g2_o21ai_1 _28360_ (.B1(_14728_),
    .Y(_14748_),
    .A1(net7291),
    .A2(_14725_));
 sg13g2_o21ai_1 _28361_ (.B1(net5766),
    .Y(_14749_),
    .A1(net6432),
    .A2(_14637_));
 sg13g2_nand2_1 _28362_ (.Y(_14750_),
    .A(_13527_),
    .B(net6445));
 sg13g2_o21ai_1 _28363_ (.B1(_14750_),
    .Y(_14751_),
    .A1(net6445),
    .A2(_14640_));
 sg13g2_a22oi_1 _28364_ (.Y(_14752_),
    .B1(_14751_),
    .B2(net5766),
    .A2(_14749_),
    .A1(_06240_));
 sg13g2_o21ai_1 _28365_ (.B1(net5766),
    .Y(_14753_),
    .A1(net6432),
    .A2(_14636_));
 sg13g2_nand2_1 _28366_ (.Y(_14754_),
    .A(_13532_),
    .B(net6442));
 sg13g2_o21ai_1 _28367_ (.B1(_14754_),
    .Y(_14755_),
    .A1(net6442),
    .A2(_14638_));
 sg13g2_a22oi_1 _28368_ (.Y(_14756_),
    .B1(_14755_),
    .B2(net5766),
    .A2(_14753_),
    .A1(_06241_));
 sg13g2_and2_1 _28369_ (.A(_00213_),
    .B(_14633_),
    .X(_14757_));
 sg13g2_nand2_1 _28370_ (.Y(_14758_),
    .A(_00213_),
    .B(_14633_));
 sg13g2_nor2_1 _28371_ (.A(_14621_),
    .B(_14758_),
    .Y(_14759_));
 sg13g2_a21o_1 _28372_ (.A2(_14759_),
    .A1(_00217_),
    .B1(net6431),
    .X(_14760_));
 sg13g2_a21oi_1 _28373_ (.A1(net5762),
    .A2(_14760_),
    .Y(_14761_),
    .B1(_00218_));
 sg13g2_nand3_1 _28374_ (.B(_00217_),
    .C(_14759_),
    .A(_00218_),
    .Y(_14762_));
 sg13g2_nand2_1 _28375_ (.Y(_14763_),
    .A(_13537_),
    .B(net6442));
 sg13g2_o21ai_1 _28376_ (.B1(_14763_),
    .Y(_14764_),
    .A1(net6444),
    .A2(_14762_));
 sg13g2_a21oi_1 _28377_ (.A1(net5762),
    .A2(_14764_),
    .Y(_14765_),
    .B1(_14761_));
 sg13g2_nand2b_1 _28378_ (.Y(_14766_),
    .B(_14759_),
    .A_N(_14607_));
 sg13g2_a21oi_1 _28379_ (.A1(net6707),
    .A2(_14567_),
    .Y(_14767_),
    .B1(_00217_));
 sg13g2_mux2_1 _28380_ (.A0(_01280_),
    .A1(_00634_),
    .S(net7868),
    .X(_14768_));
 sg13g2_nand3_1 _28381_ (.B(net6136),
    .C(net6433),
    .A(net6707),
    .Y(_14769_));
 sg13g2_mux2_1 _28382_ (.A0(_00217_),
    .A1(_14767_),
    .S(_14766_),
    .X(_14770_));
 sg13g2_nor2b_1 _28383_ (.A(_14770_),
    .B_N(_14769_),
    .Y(_14771_));
 sg13g2_nand2_1 _28384_ (.Y(_14772_),
    .A(_00214_),
    .B(_14757_));
 sg13g2_and3_1 _28385_ (.X(_14773_),
    .A(_00215_),
    .B(_00214_),
    .C(_14757_));
 sg13g2_o21ai_1 _28386_ (.B1(net5763),
    .Y(_14774_),
    .A1(net6431),
    .A2(_14773_));
 sg13g2_nand3_1 _28387_ (.B(net6438),
    .C(_14773_),
    .A(_00216_),
    .Y(_14775_));
 sg13g2_nand2_1 _28388_ (.Y(_14776_),
    .A(_13547_),
    .B(net6444));
 sg13g2_nand2_1 _28389_ (.Y(_14777_),
    .A(_14775_),
    .B(_14776_));
 sg13g2_a22oi_1 _28390_ (.Y(_14778_),
    .B1(_14777_),
    .B2(net5763),
    .A2(_14774_),
    .A1(_06242_));
 sg13g2_nand2_1 _28391_ (.Y(_14779_),
    .A(net6438),
    .B(_14772_));
 sg13g2_a21oi_1 _28392_ (.A1(net5763),
    .A2(_14779_),
    .Y(_14780_),
    .B1(_00215_));
 sg13g2_nand2_1 _28393_ (.Y(_14781_),
    .A(_13553_),
    .B(net6443));
 sg13g2_mux2_1 _28394_ (.A0(_14773_),
    .A1(_13553_),
    .S(net6431),
    .X(_14782_));
 sg13g2_a21oi_1 _28395_ (.A1(net5763),
    .A2(_14782_),
    .Y(_14783_),
    .B1(_14780_));
 sg13g2_inv_1 _28396_ (.Y(_14784_),
    .A(_01731_));
 sg13g2_o21ai_1 _28397_ (.B1(net5763),
    .Y(_14785_),
    .A1(net6431),
    .A2(_14757_));
 sg13g2_nand2_1 _28398_ (.Y(_14786_),
    .A(_13559_),
    .B(net6444));
 sg13g2_o21ai_1 _28399_ (.B1(_14786_),
    .Y(_14787_),
    .A1(net6444),
    .A2(_14772_));
 sg13g2_a22oi_1 _28400_ (.Y(_14788_),
    .B1(_14787_),
    .B2(net5763),
    .A2(_14785_),
    .A1(_06247_));
 sg13g2_nand2b_1 _28401_ (.Y(_14789_),
    .B(_14634_),
    .A_N(net6431));
 sg13g2_a21oi_1 _28402_ (.A1(net5763),
    .A2(_14789_),
    .Y(_14790_),
    .B1(_00213_));
 sg13g2_a22oi_1 _28403_ (.Y(_14791_),
    .B1(_14768_),
    .B2(net7833),
    .A2(net7527),
    .A1(_00928_));
 sg13g2_o21ai_1 _28404_ (.B1(_14585_),
    .Y(_14792_),
    .A1(net6444),
    .A2(_14758_));
 sg13g2_a21oi_1 _28405_ (.A1(net5763),
    .A2(_14792_),
    .Y(_14793_),
    .B1(_14790_));
 sg13g2_nor2_1 _28406_ (.A(_14620_),
    .B(_14631_),
    .Y(_14794_));
 sg13g2_or2_1 _28407_ (.X(_14795_),
    .B(_14631_),
    .A(_14620_));
 sg13g2_nor2_1 _28408_ (.A(_14617_),
    .B(_14795_),
    .Y(_14796_));
 sg13g2_nor3_1 _28409_ (.A(_06263_),
    .B(_14617_),
    .C(_14795_),
    .Y(_14797_));
 sg13g2_nand2_1 _28410_ (.Y(_14798_),
    .A(_00209_),
    .B(_14796_));
 sg13g2_nand2_1 _28411_ (.Y(_14799_),
    .A(_00210_),
    .B(_14797_));
 sg13g2_nand2_1 _28412_ (.Y(_14800_),
    .A(net6439),
    .B(_14799_));
 sg13g2_a21oi_1 _28413_ (.A1(net5762),
    .A2(_14800_),
    .Y(_14801_),
    .B1(_00212_));
 sg13g2_nand3_1 _28414_ (.B(_00210_),
    .C(_14797_),
    .A(_00212_),
    .Y(_14802_));
 sg13g2_o21ai_1 _28415_ (.B1(_14588_),
    .Y(_14803_),
    .A1(net6442),
    .A2(_14802_));
 sg13g2_a21oi_1 _28416_ (.A1(net5762),
    .A2(_14803_),
    .Y(_14804_),
    .B1(_14801_));
 sg13g2_o21ai_1 _28417_ (.B1(net5822),
    .Y(_14805_),
    .A1(net6441),
    .A2(_14573_));
 sg13g2_nand2b_1 _28418_ (.Y(_14806_),
    .B(net7868),
    .A_N(_00698_));
 sg13g2_nand2_1 _28419_ (.Y(_14807_),
    .A(net6437),
    .B(_14574_));
 sg13g2_o21ai_1 _28420_ (.B1(_14807_),
    .Y(_14808_),
    .A1(_13657_),
    .A2(net6437));
 sg13g2_a22oi_1 _28421_ (.Y(_14809_),
    .B1(_14808_),
    .B2(net5820),
    .A2(_14805_),
    .A1(_06255_));
 sg13g2_nand2_1 _28422_ (.Y(_14810_),
    .A(net6439),
    .B(_14798_));
 sg13g2_a21oi_1 _28423_ (.A1(net5761),
    .A2(_14810_),
    .Y(_14811_),
    .B1(_00210_));
 sg13g2_o21ai_1 _28424_ (.B1(_14806_),
    .Y(_14812_),
    .A1(net7868),
    .A2(_00666_));
 sg13g2_o21ai_1 _28425_ (.B1(_14593_),
    .Y(_14813_),
    .A1(net6442),
    .A2(_14799_));
 sg13g2_inv_1 _28426_ (.Y(_14814_),
    .A(_01730_));
 sg13g2_a21oi_1 _28427_ (.A1(net5762),
    .A2(_14813_),
    .Y(_14815_),
    .B1(_14811_));
 sg13g2_o21ai_1 _28428_ (.B1(net5761),
    .Y(_14816_),
    .A1(net6431),
    .A2(_14796_));
 sg13g2_o21ai_1 _28429_ (.B1(_14603_),
    .Y(_14817_),
    .A1(net6442),
    .A2(_14798_));
 sg13g2_a22oi_1 _28430_ (.Y(_14818_),
    .B1(_14817_),
    .B2(net5761),
    .A2(_14816_),
    .A1(_06263_));
 sg13g2_o21ai_1 _28431_ (.B1(net6439),
    .Y(_14819_),
    .A1(_14616_),
    .A2(_14795_));
 sg13g2_nand2_1 _28432_ (.Y(_14820_),
    .A(net5765),
    .B(_14819_));
 sg13g2_nor4_1 _28433_ (.A(_06266_),
    .B(net6433),
    .C(_14616_),
    .D(_14795_),
    .Y(_14821_));
 sg13g2_a21o_1 _28434_ (.A2(net6433),
    .A1(_13634_),
    .B1(_14821_),
    .X(_14822_));
 sg13g2_a22oi_1 _28435_ (.Y(_14823_),
    .B1(_14822_),
    .B2(_14609_),
    .A2(_14820_),
    .A1(_06266_));
 sg13g2_mux2_1 _28436_ (.A0(_00730_),
    .A1(_00762_),
    .S(net7868),
    .X(_14824_));
 sg13g2_nand3_1 _28437_ (.B(_14614_),
    .C(_14794_),
    .A(_00206_),
    .Y(_14825_));
 sg13g2_nand2_1 _28438_ (.Y(_14826_),
    .A(net6439),
    .B(_14825_));
 sg13g2_a21oi_1 _28439_ (.A1(_14609_),
    .A2(_14826_),
    .Y(_14827_),
    .B1(_00207_));
 sg13g2_nand2_1 _28440_ (.Y(_14828_),
    .A(net6440),
    .B(_14794_));
 sg13g2_o21ai_1 _28441_ (.B1(_14740_),
    .Y(_14829_),
    .A1(_14616_),
    .A2(_14828_));
 sg13g2_a21oi_1 _28442_ (.A1(_14609_),
    .A2(_14829_),
    .Y(_14830_),
    .B1(_14827_));
 sg13g2_o21ai_1 _28443_ (.B1(net6440),
    .Y(_14831_),
    .A1(_14615_),
    .A2(_14795_));
 sg13g2_a21oi_1 _28444_ (.A1(_14609_),
    .A2(_14831_),
    .Y(_14832_),
    .B1(_00206_));
 sg13g2_nand4_1 _28445_ (.B(net6440),
    .C(_14614_),
    .A(_00206_),
    .Y(_14833_),
    .D(_14794_));
 sg13g2_o21ai_1 _28446_ (.B1(_14833_),
    .Y(_14834_),
    .A1(_13657_),
    .A2(net6440));
 sg13g2_a21oi_1 _28447_ (.A1(_14609_),
    .A2(_14834_),
    .Y(_14835_),
    .B1(_14832_));
 sg13g2_o21ai_1 _28448_ (.B1(net6440),
    .Y(_14836_),
    .A1(_14612_),
    .A2(_14795_));
 sg13g2_a21oi_1 _28449_ (.A1(net5765),
    .A2(_14836_),
    .Y(_14837_),
    .B1(_00205_));
 sg13g2_o21ai_1 _28450_ (.B1(net7530),
    .Y(_14838_),
    .A1(net7520),
    .A2(_14824_));
 sg13g2_nand2_1 _28451_ (.Y(_14839_),
    .A(_13704_),
    .B(net6446));
 sg13g2_o21ai_1 _28452_ (.B1(_14839_),
    .Y(_14840_),
    .A1(_14615_),
    .A2(_14828_));
 sg13g2_a221oi_1 _28453_ (.B2(net7515),
    .C1(_14838_),
    .B1(_14812_),
    .A1(net7484),
    .Y(_14841_),
    .A2(_14791_));
 sg13g2_a21oi_1 _28454_ (.A1(net5765),
    .A2(_14840_),
    .Y(_14842_),
    .B1(_14837_));
 sg13g2_a21o_1 _28455_ (.A2(_14794_),
    .A1(_00203_),
    .B1(net6433),
    .X(_14843_));
 sg13g2_a21oi_1 _28456_ (.A1(net5765),
    .A2(_14843_),
    .Y(_14844_),
    .B1(_00204_));
 sg13g2_nand2_1 _28457_ (.Y(_14845_),
    .A(net6454),
    .B(net6446));
 sg13g2_o21ai_1 _28458_ (.B1(_14845_),
    .Y(_14846_),
    .A1(_14612_),
    .A2(_14828_));
 sg13g2_a21oi_1 _28459_ (.A1(net5765),
    .A2(_14846_),
    .Y(_14847_),
    .B1(_14844_));
 sg13g2_o21ai_1 _28460_ (.B1(net5765),
    .Y(_14848_),
    .A1(net6433),
    .A2(_14794_));
 sg13g2_nand2_1 _28461_ (.Y(_14849_),
    .A(_13874_),
    .B(net6446));
 sg13g2_o21ai_1 _28462_ (.B1(_14849_),
    .Y(_14850_),
    .A1(_06280_),
    .A2(_14828_));
 sg13g2_a22oi_1 _28463_ (.Y(_14851_),
    .B1(_14850_),
    .B2(net5765),
    .A2(_14848_),
    .A1(_06280_));
 sg13g2_mux2_1 _28464_ (.A0(_01281_),
    .A1(_01316_),
    .S(net7864),
    .X(_14852_));
 sg13g2_and2_1 _28465_ (.A(_00197_),
    .B(_14630_),
    .X(_14853_));
 sg13g2_nand2_1 _28466_ (.Y(_14854_),
    .A(_00197_),
    .B(_14630_));
 sg13g2_and2_1 _28467_ (.A(_00198_),
    .B(_14853_),
    .X(_14855_));
 sg13g2_nand2_1 _28468_ (.Y(_14856_),
    .A(_00198_),
    .B(_14853_));
 sg13g2_nand2_1 _28469_ (.Y(_14857_),
    .A(_00199_),
    .B(_14855_));
 sg13g2_nand3_1 _28470_ (.B(_00199_),
    .C(_14855_),
    .A(_00201_),
    .Y(_14858_));
 sg13g2_nand2_1 _28471_ (.Y(_14859_),
    .A(net6435),
    .B(_14858_));
 sg13g2_inv_1 _28472_ (.Y(_14860_),
    .A(_01728_));
 sg13g2_nor2_1 _28473_ (.A(net7520),
    .B(_14852_),
    .Y(_14861_));
 sg13g2_a21oi_1 _28474_ (.A1(net5829),
    .A2(_14859_),
    .Y(_14862_),
    .B1(_00202_));
 sg13g2_nor2_1 _28475_ (.A(net6447),
    .B(_14858_),
    .Y(_14863_));
 sg13g2_a22oi_1 _28476_ (.Y(_14864_),
    .B1(_14863_),
    .B2(_00202_),
    .A2(net6447),
    .A1(_13441_));
 sg13g2_inv_1 _28477_ (.Y(_14865_),
    .A(_14864_));
 sg13g2_a21oi_1 _28478_ (.A1(net5828),
    .A2(_14865_),
    .Y(_14866_),
    .B1(_14862_));
 sg13g2_nand2_1 _28479_ (.Y(_14867_),
    .A(net6435),
    .B(_14857_));
 sg13g2_a21oi_1 _28480_ (.A1(net5829),
    .A2(_14867_),
    .Y(_14868_),
    .B1(_00201_));
 sg13g2_o21ai_1 _28481_ (.B1(_14670_),
    .Y(_14869_),
    .A1(net6447),
    .A2(_14858_));
 sg13g2_a21oi_1 _28482_ (.A1(net5828),
    .A2(_14869_),
    .Y(_14870_),
    .B1(_14868_));
 sg13g2_nand2_1 _28483_ (.Y(_14871_),
    .A(net6437),
    .B(_14573_));
 sg13g2_nand2_1 _28484_ (.Y(_14872_),
    .A(_14839_),
    .B(_14871_));
 sg13g2_o21ai_1 _28485_ (.B1(net6437),
    .Y(_14873_),
    .A1(_06328_),
    .A2(_06362_));
 sg13g2_a21oi_1 _28486_ (.A1(net5822),
    .A2(_14873_),
    .Y(_14874_),
    .B1(_00200_));
 sg13g2_a21oi_1 _28487_ (.A1(net5820),
    .A2(_14872_),
    .Y(_14875_),
    .B1(_14874_));
 sg13g2_nand2_1 _28488_ (.Y(_14876_),
    .A(net6435),
    .B(_14856_));
 sg13g2_mux2_1 _28489_ (.A0(_01069_),
    .A1(_01105_),
    .S(net7917),
    .X(_14877_));
 sg13g2_a21oi_1 _28490_ (.A1(net5829),
    .A2(_14876_),
    .Y(_14878_),
    .B1(_00199_));
 sg13g2_o21ai_1 _28491_ (.B1(_14674_),
    .Y(_14879_),
    .A1(net6448),
    .A2(_14857_));
 sg13g2_nor2_1 _28492_ (.A(_10182_),
    .B(_14877_),
    .Y(_14880_));
 sg13g2_a21oi_1 _28493_ (.A1(net5829),
    .A2(_14879_),
    .Y(_14881_),
    .B1(_14878_));
 sg13g2_nand2_1 _28494_ (.Y(_14882_),
    .A(_14571_),
    .B(_14854_));
 sg13g2_a21oi_1 _28495_ (.A1(net5829),
    .A2(_14882_),
    .Y(_14883_),
    .B1(_00198_));
 sg13g2_o21ai_1 _28496_ (.B1(_14679_),
    .Y(_14884_),
    .A1(net6448),
    .A2(_14856_));
 sg13g2_a21oi_1 _28497_ (.A1(net5829),
    .A2(_14884_),
    .Y(_14885_),
    .B1(_14883_));
 sg13g2_nand2_1 _28498_ (.Y(_14886_),
    .A(_14571_),
    .B(_14631_));
 sg13g2_a21oi_1 _28499_ (.A1(net5832),
    .A2(_14886_),
    .Y(_14887_),
    .B1(_00197_));
 sg13g2_o21ai_1 _28500_ (.B1(_14687_),
    .Y(_14888_),
    .A1(net6448),
    .A2(_14854_));
 sg13g2_a21oi_1 _28501_ (.A1(net5832),
    .A2(_14888_),
    .Y(_14889_),
    .B1(_14887_));
 sg13g2_nand2_1 _28502_ (.Y(_14890_),
    .A(_00185_),
    .B(_14627_));
 sg13g2_and3_1 _28503_ (.X(_14891_),
    .A(_00186_),
    .B(_00185_),
    .C(_14627_));
 sg13g2_inv_1 _28504_ (.Y(_14892_),
    .A(_14891_));
 sg13g2_and2_1 _28505_ (.A(_00187_),
    .B(_14891_),
    .X(_14893_));
 sg13g2_nand2_1 _28506_ (.Y(_14894_),
    .A(_00187_),
    .B(_14891_));
 sg13g2_nor2_1 _28507_ (.A(_14611_),
    .B(_14894_),
    .Y(_14895_));
 sg13g2_or2_1 _28508_ (.X(_14896_),
    .B(_14895_),
    .A(net6450));
 sg13g2_mux2_1 _28509_ (.A0(_01140_),
    .A1(_01175_),
    .S(net7917),
    .X(_14897_));
 sg13g2_a21oi_1 _28510_ (.A1(net5832),
    .A2(_14896_),
    .Y(_14898_),
    .B1(_00196_));
 sg13g2_nand2_1 _28511_ (.Y(_14899_),
    .A(_00196_),
    .B(_14895_));
 sg13g2_nor2_1 _28512_ (.A(net7460),
    .B(_14897_),
    .Y(_14900_));
 sg13g2_o21ai_1 _28513_ (.B1(_14692_),
    .Y(_14901_),
    .A1(net6450),
    .A2(_14899_));
 sg13g2_a21oi_1 _28514_ (.A1(net5829),
    .A2(_14901_),
    .Y(_14902_),
    .B1(_14898_));
 sg13g2_and2_1 _28515_ (.A(_00188_),
    .B(_14893_),
    .X(_14903_));
 sg13g2_nand2_1 _28516_ (.Y(_14904_),
    .A(_00188_),
    .B(_14893_));
 sg13g2_and2_1 _28517_ (.A(_00190_),
    .B(_14903_),
    .X(_14905_));
 sg13g2_nand2_1 _28518_ (.Y(_14906_),
    .A(_00190_),
    .B(_14903_));
 sg13g2_and2_1 _28519_ (.A(_00191_),
    .B(_14905_),
    .X(_14907_));
 sg13g2_nand2_1 _28520_ (.Y(_14908_),
    .A(_00191_),
    .B(_14905_));
 sg13g2_and2_1 _28521_ (.A(_00192_),
    .B(_14907_),
    .X(_14909_));
 sg13g2_nand2_1 _28522_ (.Y(_14910_),
    .A(_00192_),
    .B(_14907_));
 sg13g2_and2_1 _28523_ (.A(_00193_),
    .B(_14909_),
    .X(_14911_));
 sg13g2_nand2_1 _28524_ (.Y(_14912_),
    .A(_00193_),
    .B(_14909_));
 sg13g2_nand2_1 _28525_ (.Y(_14913_),
    .A(_00194_),
    .B(_14911_));
 sg13g2_nand2_1 _28526_ (.Y(_14914_),
    .A(net6436),
    .B(_14913_));
 sg13g2_a21oi_1 _28527_ (.A1(net5831),
    .A2(_14914_),
    .Y(_14915_),
    .B1(_00195_));
 sg13g2_nand3_1 _28528_ (.B(_00194_),
    .C(_14911_),
    .A(_00195_),
    .Y(_14916_));
 sg13g2_o21ai_1 _28529_ (.B1(_14700_),
    .Y(_14917_),
    .A1(net6451),
    .A2(_14916_));
 sg13g2_a21oi_1 _28530_ (.A1(net5831),
    .A2(_14917_),
    .Y(_14918_),
    .B1(_14915_));
 sg13g2_nand2_1 _28531_ (.Y(_14919_),
    .A(net6436),
    .B(_14912_));
 sg13g2_a21oi_1 _28532_ (.A1(net5831),
    .A2(_14919_),
    .Y(_14920_),
    .B1(_00194_));
 sg13g2_o21ai_1 _28533_ (.B1(_14705_),
    .Y(_14921_),
    .A1(net6451),
    .A2(_14913_));
 sg13g2_a21oi_1 _28534_ (.A1(net5831),
    .A2(_14921_),
    .Y(_14922_),
    .B1(_14920_));
 sg13g2_nand2_1 _28535_ (.Y(_14923_),
    .A(net6436),
    .B(_14910_));
 sg13g2_a21oi_1 _28536_ (.A1(net5831),
    .A2(_14923_),
    .Y(_14924_),
    .B1(_00193_));
 sg13g2_o21ai_1 _28537_ (.B1(_14710_),
    .Y(_14925_),
    .A1(net6452),
    .A2(_14912_));
 sg13g2_a21oi_1 _28538_ (.A1(net5831),
    .A2(_14925_),
    .Y(_14926_),
    .B1(_14924_));
 sg13g2_nand2_1 _28539_ (.Y(_14927_),
    .A(net6436),
    .B(_14908_));
 sg13g2_a21oi_1 _28540_ (.A1(net5830),
    .A2(_14927_),
    .Y(_14928_),
    .B1(_00192_));
 sg13g2_mux2_1 _28541_ (.A0(_01210_),
    .A1(_01245_),
    .S(net7864),
    .X(_14929_));
 sg13g2_o21ai_1 _28542_ (.B1(_14717_),
    .Y(_14930_),
    .A1(net6450),
    .A2(_14910_));
 sg13g2_a21oi_1 _28543_ (.A1(net5830),
    .A2(_14930_),
    .Y(_14931_),
    .B1(_14928_));
 sg13g2_nand2_1 _28544_ (.Y(_14932_),
    .A(net6436),
    .B(_14906_));
 sg13g2_a21oi_1 _28545_ (.A1(net5830),
    .A2(_14932_),
    .Y(_14933_),
    .B1(_00191_));
 sg13g2_o21ai_1 _28546_ (.B1(_14723_),
    .Y(_14934_),
    .A1(net6450),
    .A2(_14908_));
 sg13g2_o21ai_1 _28547_ (.B1(net7502),
    .Y(_14935_),
    .A1(net7504),
    .A2(_14929_));
 sg13g2_nor4_1 _28548_ (.A(_14861_),
    .B(_14880_),
    .C(_14900_),
    .D(_14935_),
    .Y(_14936_));
 sg13g2_a21oi_1 _28549_ (.A1(net5830),
    .A2(_14934_),
    .Y(_14937_),
    .B1(_14933_));
 sg13g2_nand2_1 _28550_ (.Y(_14938_),
    .A(net6436),
    .B(_14904_));
 sg13g2_a21oi_1 _28551_ (.A1(net5830),
    .A2(_14938_),
    .Y(_14939_),
    .B1(_00190_));
 sg13g2_o21ai_1 _28552_ (.B1(_14729_),
    .Y(_14940_),
    .A1(net6450),
    .A2(_14906_));
 sg13g2_a21oi_1 _28553_ (.A1(net5830),
    .A2(_14940_),
    .Y(_14941_),
    .B1(_14939_));
 sg13g2_nand3_1 _28554_ (.B(_00178_),
    .C(net6437),
    .A(_00189_),
    .Y(_14942_));
 sg13g2_o21ai_1 _28555_ (.B1(_14942_),
    .Y(_14943_),
    .A1(_13780_),
    .A2(net6437));
 sg13g2_o21ai_1 _28556_ (.B1(net5822),
    .Y(_14944_),
    .A1(_00178_),
    .A2(net6453));
 sg13g2_mux2_1 _28557_ (.A0(_01562_),
    .A1(_01597_),
    .S(net7876),
    .X(_14945_));
 sg13g2_a22oi_1 _28558_ (.Y(_14946_),
    .B1(_14944_),
    .B2(_06328_),
    .A2(_14943_),
    .A1(net5822));
 sg13g2_nand2_1 _28559_ (.Y(_14947_),
    .A(net6436),
    .B(_14894_));
 sg13g2_nand2_1 _28560_ (.Y(_14948_),
    .A(_10980_),
    .B(_14945_));
 sg13g2_a21oi_1 _28561_ (.A1(net5830),
    .A2(_14947_),
    .Y(_14949_),
    .B1(_00188_));
 sg13g2_o21ai_1 _28562_ (.B1(_14733_),
    .Y(_14950_),
    .A1(net6450),
    .A2(_14904_));
 sg13g2_a21oi_1 _28563_ (.A1(net5830),
    .A2(_14950_),
    .Y(_14951_),
    .B1(_14949_));
 sg13g2_nand2b_1 _28564_ (.Y(_14952_),
    .B(_14892_),
    .A_N(net6432));
 sg13g2_a21oi_1 _28565_ (.A1(net5824),
    .A2(_14952_),
    .Y(_14953_),
    .B1(_00187_));
 sg13g2_o21ai_1 _28566_ (.B1(_14737_),
    .Y(_14954_),
    .A1(net6445),
    .A2(_14894_));
 sg13g2_mux2_1 _28567_ (.A0(_01492_),
    .A1(_01527_),
    .S(net7870),
    .X(_14955_));
 sg13g2_a21oi_1 _28568_ (.A1(net5824),
    .A2(_14954_),
    .Y(_14956_),
    .B1(_14953_));
 sg13g2_nand2_1 _28569_ (.Y(_14957_),
    .A(net6439),
    .B(_14890_));
 sg13g2_nand3_1 _28570_ (.B(net7497),
    .C(_14955_),
    .A(net7513),
    .Y(_14958_));
 sg13g2_a21oi_1 _28571_ (.A1(net5824),
    .A2(_14957_),
    .Y(_14959_),
    .B1(_00186_));
 sg13g2_o21ai_1 _28572_ (.B1(_14745_),
    .Y(_14960_),
    .A1(net6445),
    .A2(_14892_));
 sg13g2_a21oi_1 _28573_ (.A1(net5824),
    .A2(_14960_),
    .Y(_14961_),
    .B1(_14959_));
 sg13g2_nand2_1 _28574_ (.Y(_14962_),
    .A(net6439),
    .B(_14628_));
 sg13g2_a21oi_1 _28575_ (.A1(net5824),
    .A2(_14962_),
    .Y(_14963_),
    .B1(_00185_));
 sg13g2_o21ai_1 _28576_ (.B1(_14750_),
    .Y(_14964_),
    .A1(net6445),
    .A2(_14890_));
 sg13g2_mux2_1 _28577_ (.A0(_01421_),
    .A1(_01457_),
    .S(net7876),
    .X(_14965_));
 sg13g2_a21oi_1 _28578_ (.A1(net5824),
    .A2(_14964_),
    .Y(_14966_),
    .B1(_14963_));
 sg13g2_nand2b_1 _28579_ (.Y(_14967_),
    .B(_14626_),
    .A_N(net6432));
 sg13g2_a21oi_1 _28580_ (.A1(net5824),
    .A2(_14967_),
    .Y(_14968_),
    .B1(_00184_));
 sg13g2_nand3_1 _28581_ (.B(net7463),
    .C(_14965_),
    .A(net7497),
    .Y(_14969_));
 sg13g2_o21ai_1 _28582_ (.B1(_14754_),
    .Y(_14970_),
    .A1(net6442),
    .A2(_14628_));
 sg13g2_a21oi_1 _28583_ (.A1(net5827),
    .A2(_14970_),
    .Y(_14971_),
    .B1(_14968_));
 sg13g2_or2_1 _28584_ (.X(_14972_),
    .B(_14624_),
    .A(net6432));
 sg13g2_a21oi_1 _28585_ (.A1(net5827),
    .A2(_14972_),
    .Y(_14973_),
    .B1(_00183_));
 sg13g2_o21ai_1 _28586_ (.B1(_14763_),
    .Y(_14974_),
    .A1(net6442),
    .A2(_14626_));
 sg13g2_mux2_1 _28587_ (.A0(_01351_),
    .A1(_01386_),
    .S(net7876),
    .X(_14975_));
 sg13g2_a21oi_1 _28588_ (.A1(net5827),
    .A2(_14974_),
    .Y(_14976_),
    .B1(_14973_));
 sg13g2_nand3_1 _28589_ (.B(_00179_),
    .C(_14579_),
    .A(_00241_),
    .Y(_14977_));
 sg13g2_nand4_1 _28590_ (.B(_00180_),
    .C(_00179_),
    .A(_00241_),
    .Y(_14978_),
    .D(_14579_));
 sg13g2_or2_1 _28591_ (.X(_14979_),
    .B(_14978_),
    .A(_06345_));
 sg13g2_nand3_1 _28592_ (.B(net7472),
    .C(_14975_),
    .A(net7497),
    .Y(_14980_));
 sg13g2_nand2_1 _28593_ (.Y(_14981_),
    .A(net6438),
    .B(_14979_));
 sg13g2_a21oi_1 _28594_ (.A1(net5825),
    .A2(_14981_),
    .Y(_14982_),
    .B1(_00182_));
 sg13g2_nor2_1 _28595_ (.A(net6443),
    .B(_14979_),
    .Y(_14983_));
 sg13g2_a22oi_1 _28596_ (.Y(_14984_),
    .B1(_14983_),
    .B2(_00182_),
    .A2(net6443),
    .A1(net6136));
 sg13g2_inv_1 _28597_ (.Y(_14985_),
    .A(_14984_));
 sg13g2_a21oi_1 _28598_ (.A1(net5825),
    .A2(_14985_),
    .Y(_14986_),
    .B1(_14982_));
 sg13g2_nand2_1 _28599_ (.Y(_14987_),
    .A(net6438),
    .B(_14978_));
 sg13g2_a21oi_1 _28600_ (.A1(net5825),
    .A2(_14987_),
    .Y(_14988_),
    .B1(_00181_));
 sg13g2_o21ai_1 _28601_ (.B1(_14776_),
    .Y(_14989_),
    .A1(net6443),
    .A2(_14979_));
 sg13g2_a21oi_1 _28602_ (.A1(net5825),
    .A2(_14989_),
    .Y(_14990_),
    .B1(_14988_));
 sg13g2_nand2_1 _28603_ (.Y(_14991_),
    .A(net6438),
    .B(_14977_));
 sg13g2_a21oi_1 _28604_ (.A1(net5825),
    .A2(_14991_),
    .Y(_14992_),
    .B1(_00180_));
 sg13g2_mux2_1 _28605_ (.A0(_00858_),
    .A1(_00893_),
    .S(net7870),
    .X(_14993_));
 sg13g2_o21ai_1 _28606_ (.B1(_14781_),
    .Y(_14994_),
    .A1(net6443),
    .A2(_14978_));
 sg13g2_nand3_1 _28607_ (.B(net7463),
    .C(_14993_),
    .A(net7544),
    .Y(_14995_));
 sg13g2_a21oi_1 _28608_ (.A1(net5825),
    .A2(_14994_),
    .Y(_14996_),
    .B1(_14992_));
 sg13g2_nand2_1 _28609_ (.Y(_14997_),
    .A(net6438),
    .B(_14584_));
 sg13g2_a21oi_1 _28610_ (.A1(net5825),
    .A2(_14997_),
    .Y(_14998_),
    .B1(_00179_));
 sg13g2_o21ai_1 _28611_ (.B1(_14786_),
    .Y(_14999_),
    .A1(net6443),
    .A2(_14977_));
 sg13g2_a21oi_1 _28612_ (.A1(net5825),
    .A2(_14999_),
    .Y(_15000_),
    .B1(_14998_));
 sg13g2_o21ai_1 _28613_ (.B1(net5822),
    .Y(_15001_),
    .A1(_13873_),
    .A2(net6437));
 sg13g2_a21oi_1 _28614_ (.A1(_13873_),
    .A2(_14581_),
    .Y(_15002_),
    .B1(_06362_));
 sg13g2_mux2_1 _28615_ (.A0(_00794_),
    .A1(_00826_),
    .S(net7870),
    .X(_15003_));
 sg13g2_nand3_1 _28616_ (.B(net7472),
    .C(_15003_),
    .A(net7544),
    .Y(_15004_));
 sg13g2_a22oi_1 _28617_ (.Y(_15005_),
    .B1(_15002_),
    .B2(net5822),
    .A2(_15001_),
    .A1(_06362_));
 sg13g2_nor2_1 _28618_ (.A(net6825),
    .B(_14565_),
    .Y(_15006_));
 sg13g2_nand2_1 _28619_ (.Y(_15007_),
    .A(net6711),
    .B(_15006_));
 sg13g2_nor2_1 _28620_ (.A(net6825),
    .B(_14566_),
    .Y(_15008_));
 sg13g2_and2_1 _28621_ (.A(_06920_),
    .B(_15006_),
    .X(_15009_));
 sg13g2_and2_1 _28622_ (.A(net6707),
    .B(_15008_),
    .X(_15010_));
 sg13g2_a21oi_1 _28623_ (.A1(_00112_),
    .A2(_15007_),
    .Y(_15011_),
    .B1(_15010_));
 sg13g2_a21o_1 _28624_ (.A2(_15007_),
    .A1(_00112_),
    .B1(_15010_),
    .X(_15012_));
 sg13g2_nor2_1 _28625_ (.A(_06569_),
    .B(_06615_),
    .Y(_15013_));
 sg13g2_and2_1 _28626_ (.A(_00136_),
    .B(_15013_),
    .X(_15014_));
 sg13g2_nand4_1 _28627_ (.B(_00158_),
    .C(_00147_),
    .A(_00169_),
    .Y(_15015_),
    .D(_15014_));
 sg13g2_nor2_1 _28628_ (.A(_06379_),
    .B(_15015_),
    .Y(_15016_));
 sg13g2_nand2_1 _28629_ (.Y(_15017_),
    .A(_00175_),
    .B(_15016_));
 sg13g2_and3_1 _28630_ (.X(_15018_),
    .A(_00176_),
    .B(_00175_),
    .C(_15016_));
 sg13g2_inv_1 _28631_ (.Y(_15019_),
    .A(_15018_));
 sg13g2_nor3_1 _28632_ (.A(net6825),
    .B(_06921_),
    .C(_14565_),
    .Y(_15020_));
 sg13g2_nand2b_1 _28633_ (.Y(_15021_),
    .B(_15006_),
    .A_N(_06921_));
 sg13g2_and2_1 _28634_ (.A(_06941_),
    .B(_15008_),
    .X(_15022_));
 sg13g2_mux2_1 _28635_ (.A0(_00929_),
    .A1(_00964_),
    .S(net7871),
    .X(_15023_));
 sg13g2_o21ai_1 _28636_ (.B1(net6061),
    .Y(_15024_),
    .A1(_15018_),
    .A2(net6427));
 sg13g2_nand2_1 _28637_ (.Y(_15025_),
    .A(_00177_),
    .B(_15018_));
 sg13g2_nand2_1 _28638_ (.Y(_15026_),
    .A(_13431_),
    .B(net6428));
 sg13g2_nand3_1 _28639_ (.B(net7513),
    .C(_15023_),
    .A(net7544),
    .Y(_15027_));
 sg13g2_o21ai_1 _28640_ (.B1(_15026_),
    .Y(_15028_),
    .A1(net6415),
    .A2(_15025_));
 sg13g2_a22oi_1 _28641_ (.Y(_15029_),
    .B1(_15028_),
    .B2(net6061),
    .A2(_15024_),
    .A1(_06369_));
 sg13g2_inv_1 _28642_ (.Y(_15030_),
    .A(_01722_));
 sg13g2_nand2_1 _28643_ (.Y(_15031_),
    .A(_15017_),
    .B(net6127));
 sg13g2_nand2_1 _28644_ (.Y(_15032_),
    .A(net6159),
    .B(net6428));
 sg13g2_o21ai_1 _28645_ (.B1(_15032_),
    .Y(_15033_),
    .A1(_15019_),
    .A2(net6415));
 sg13g2_a21oi_1 _28646_ (.A1(net6061),
    .A2(_15031_),
    .Y(_15034_),
    .B1(_00176_));
 sg13g2_a21oi_1 _28647_ (.A1(net6063),
    .A2(_15033_),
    .Y(_15035_),
    .B1(_15034_));
 sg13g2_mux2_1 _28648_ (.A0(_00999_),
    .A1(_01034_),
    .S(net7871),
    .X(_15036_));
 sg13g2_o21ai_1 _28649_ (.B1(net6063),
    .Y(_15037_),
    .A1(_15016_),
    .A2(net6429));
 sg13g2_nand2_1 _28650_ (.Y(_15038_),
    .A(_13610_),
    .B(net6415));
 sg13g2_nand3_1 _28651_ (.B(net7526),
    .C(_15036_),
    .A(net7544),
    .Y(_15039_));
 sg13g2_o21ai_1 _28652_ (.B1(_15038_),
    .Y(_15040_),
    .A1(_15017_),
    .A2(net6415));
 sg13g2_a22oi_1 _28653_ (.Y(_15041_),
    .B1(_15040_),
    .B2(net6063),
    .A2(_15037_),
    .A1(_06373_));
 sg13g2_a21o_1 _28654_ (.A2(net6128),
    .A1(_15015_),
    .B1(_15012_),
    .X(_15042_));
 sg13g2_nand2_1 _28655_ (.Y(_15043_),
    .A(_15016_),
    .B(net6128));
 sg13g2_nand2_1 _28656_ (.Y(_15044_),
    .A(_13621_),
    .B(net6430));
 sg13g2_a21oi_1 _28657_ (.A1(_15043_),
    .A2(_15044_),
    .Y(_15045_),
    .B1(_15012_));
 sg13g2_a21oi_1 _28658_ (.A1(_06379_),
    .A2(_15042_),
    .Y(_15046_),
    .B1(_15045_));
 sg13g2_a21oi_1 _28659_ (.A1(_06803_),
    .A2(_14601_),
    .Y(_15047_),
    .B1(_06628_));
 sg13g2_a21oi_1 _28660_ (.A1(net6711),
    .A2(_15008_),
    .Y(_15048_),
    .B1(_15047_));
 sg13g2_nand4_1 _28661_ (.B(_00117_),
    .C(_00116_),
    .A(_00176_),
    .Y(_15049_),
    .D(_00115_));
 sg13g2_or2_1 _28662_ (.X(_15050_),
    .B(_15049_),
    .A(_06369_));
 sg13g2_nand4_1 _28663_ (.B(_00127_),
    .C(_00126_),
    .A(_00128_),
    .Y(_15051_),
    .D(_00124_));
 sg13g2_nand4_1 _28664_ (.B(_00131_),
    .C(_00130_),
    .A(_00132_),
    .Y(_15052_),
    .D(_00129_));
 sg13g2_nor2_1 _28665_ (.A(_15051_),
    .B(_15052_),
    .Y(_15053_));
 sg13g2_nand4_1 _28666_ (.B(_14969_),
    .C(_14980_),
    .A(_14948_),
    .Y(_15054_),
    .D(_15027_));
 sg13g2_nand3_1 _28667_ (.B(_00135_),
    .C(_00134_),
    .A(_00137_),
    .Y(_15055_));
 sg13g2_nand4_1 _28668_ (.B(_00139_),
    .C(_00138_),
    .A(_00140_),
    .Y(_15056_),
    .D(_00133_));
 sg13g2_nor2_1 _28669_ (.A(_15055_),
    .B(_15056_),
    .Y(_15057_));
 sg13g2_nand2_1 _28670_ (.Y(_15058_),
    .A(_00145_),
    .B(_00144_));
 sg13g2_nand3_1 _28671_ (.B(_00145_),
    .C(_00144_),
    .A(_00146_),
    .Y(_15059_));
 sg13g2_nor2_1 _28672_ (.A(_06466_),
    .B(_15059_),
    .Y(_15060_));
 sg13g2_or2_1 _28673_ (.X(_15061_),
    .B(_15059_),
    .A(_06466_));
 sg13g2_and2_1 _28674_ (.A(_00149_),
    .B(_15060_),
    .X(_15062_));
 sg13g2_nand2_1 _28675_ (.Y(_15063_),
    .A(_00149_),
    .B(_15060_));
 sg13g2_nand3_1 _28676_ (.B(_00150_),
    .C(_15062_),
    .A(_00151_),
    .Y(_15064_));
 sg13g2_nor2_1 _28677_ (.A(_06458_),
    .B(_15064_),
    .Y(_15065_));
 sg13g2_or2_1 _28678_ (.X(_15066_),
    .B(_15064_),
    .A(_06458_));
 sg13g2_nand4_1 _28679_ (.B(_14995_),
    .C(_15004_),
    .A(_14958_),
    .Y(_15067_),
    .D(_15039_));
 sg13g2_nor3_1 _28680_ (.A(_06597_),
    .B(_15017_),
    .C(_15050_),
    .Y(_15068_));
 sg13g2_nand2_1 _28681_ (.Y(_15069_),
    .A(_00119_),
    .B(_15068_));
 sg13g2_and3_1 _28682_ (.X(_15070_),
    .A(_00120_),
    .B(_00119_),
    .C(_15068_));
 sg13g2_inv_1 _28683_ (.Y(_15071_),
    .A(_15070_));
 sg13g2_nor4_1 _28684_ (.A(_14841_),
    .B(_14936_),
    .C(_15054_),
    .D(_15067_),
    .Y(_15072_));
 sg13g2_and4_1 _28685_ (.A(_00123_),
    .B(_00122_),
    .C(_00121_),
    .D(_15070_),
    .X(_15073_));
 sg13g2_and2_1 _28686_ (.A(_15053_),
    .B(_15073_),
    .X(_15074_));
 sg13g2_or4_1 _28687_ (.A(_14841_),
    .B(_14936_),
    .C(_15054_),
    .D(_15067_),
    .X(_15075_));
 sg13g2_and4_1 _28688_ (.A(_00142_),
    .B(_00141_),
    .C(_15057_),
    .D(_15074_),
    .X(_15076_));
 sg13g2_inv_1 _28689_ (.Y(_15077_),
    .A(net6748));
 sg13g2_nand2_1 _28690_ (.Y(_15078_),
    .A(_00143_),
    .B(_15076_));
 sg13g2_nand3_1 _28691_ (.B(_00153_),
    .C(_15065_),
    .A(_00154_),
    .Y(_15079_));
 sg13g2_nor2_1 _28692_ (.A(net6748),
    .B(_15079_),
    .Y(_15080_));
 sg13g2_nor3_1 _28693_ (.A(_06454_),
    .B(_15078_),
    .C(_15079_),
    .Y(_15081_));
 sg13g2_nand2_1 _28694_ (.Y(_15082_),
    .A(_00155_),
    .B(_15080_));
 sg13g2_nor2_1 _28695_ (.A(_06449_),
    .B(_15082_),
    .Y(_15083_));
 sg13g2_nand2_1 _28696_ (.Y(_15084_),
    .A(_00156_),
    .B(_15081_));
 sg13g2_nor2_1 _28697_ (.A(_06444_),
    .B(_15084_),
    .Y(_15085_));
 sg13g2_inv_1 _28698_ (.Y(_15086_),
    .A(_15085_));
 sg13g2_nand3_1 _28699_ (.B(_00159_),
    .C(_15085_),
    .A(_00160_),
    .Y(_15087_));
 sg13g2_nor2_1 _28700_ (.A(_06421_),
    .B(_15087_),
    .Y(_15088_));
 sg13g2_or2_1 _28701_ (.X(_15089_),
    .B(_15087_),
    .A(_06421_));
 sg13g2_nor2_1 _28702_ (.A(_06413_),
    .B(_15089_),
    .Y(_15090_));
 sg13g2_inv_1 _28703_ (.Y(_15091_),
    .A(_15090_));
 sg13g2_and4_1 _28704_ (.A(_00165_),
    .B(_00164_),
    .C(_00163_),
    .D(_15090_),
    .X(_15092_));
 sg13g2_nand2_1 _28705_ (.Y(_15093_),
    .A(_00166_),
    .B(_15092_));
 sg13g2_and3_1 _28706_ (.X(_15094_),
    .A(_00167_),
    .B(_00166_),
    .C(_15092_));
 sg13g2_and2_1 _28707_ (.A(_00168_),
    .B(_15094_),
    .X(_15095_));
 sg13g2_inv_1 _28708_ (.Y(_15096_),
    .A(_15095_));
 sg13g2_nor2_1 _28709_ (.A(_06387_),
    .B(_15096_),
    .Y(_15097_));
 sg13g2_nand2_1 _28710_ (.Y(_15098_),
    .A(_00171_),
    .B(_15097_));
 sg13g2_and3_1 _28711_ (.X(_15099_),
    .A(_00172_),
    .B(_00171_),
    .C(_15097_));
 sg13g2_o21ai_1 _28712_ (.B1(_15048_),
    .Y(_15100_),
    .A1(_15022_),
    .A2(_15099_));
 sg13g2_nand2b_1 _28713_ (.Y(_15101_),
    .B(net7997),
    .A_N(_01639_));
 sg13g2_nand3_1 _28714_ (.B(_15021_),
    .C(_15099_),
    .A(_00173_),
    .Y(_15102_));
 sg13g2_nand2_1 _28715_ (.Y(_15103_),
    .A(_13441_),
    .B(net6419));
 sg13g2_nand2_1 _28716_ (.Y(_15104_),
    .A(_15102_),
    .B(_15103_));
 sg13g2_o21ai_1 _28717_ (.B1(_15101_),
    .Y(_15105_),
    .A1(_01669_),
    .A2(net7478));
 sg13g2_a22oi_1 _28718_ (.Y(_15106_),
    .B1(_15104_),
    .B2(_15048_),
    .A2(_15100_),
    .A1(_06384_));
 sg13g2_nand2_1 _28719_ (.Y(_15107_),
    .A(_15021_),
    .B(_15098_));
 sg13g2_inv_1 _28720_ (.Y(_15108_),
    .A(_01720_));
 sg13g2_a21oi_1 _28721_ (.A1(net8008),
    .A2(net7273),
    .Y(_15109_),
    .B1(_15105_));
 sg13g2_a21oi_1 _28722_ (.A1(_15048_),
    .A2(_15107_),
    .Y(_15110_),
    .B1(_00172_));
 sg13g2_mux2_1 _28723_ (.A0(_15099_),
    .A1(_13446_),
    .S(net6416),
    .X(_15111_));
 sg13g2_a21oi_1 _28724_ (.A1(_15048_),
    .A2(_15111_),
    .Y(_15112_),
    .B1(_15110_));
 sg13g2_o21ai_1 _28725_ (.B1(_15109_),
    .Y(_15113_),
    .A1(_09277_),
    .A2(net7274));
 sg13g2_o21ai_1 _28726_ (.B1(net6410),
    .Y(_15114_),
    .A1(_15022_),
    .A2(_15097_));
 sg13g2_nand2_1 _28727_ (.Y(_15115_),
    .A(_13451_),
    .B(net6419));
 sg13g2_o21ai_1 _28728_ (.B1(_15115_),
    .Y(_15116_),
    .A1(net6419),
    .A2(_15098_));
 sg13g2_a22oi_1 _28729_ (.Y(_15117_),
    .B1(_15116_),
    .B2(_15048_),
    .A2(_15114_),
    .A1(_06386_));
 sg13g2_o21ai_1 _28730_ (.B1(net6410),
    .Y(_15118_),
    .A1(_15022_),
    .A2(_15095_));
 sg13g2_nand2_1 _28731_ (.Y(_15119_),
    .A(_15021_),
    .B(_15097_));
 sg13g2_nand2_1 _28732_ (.Y(_15120_),
    .A(_13458_),
    .B(net6418));
 sg13g2_nand2_1 _28733_ (.Y(_15121_),
    .A(_15119_),
    .B(_15120_));
 sg13g2_a22oi_1 _28734_ (.Y(_15122_),
    .B1(_15121_),
    .B2(net6410),
    .A2(_15118_),
    .A1(_06387_));
 sg13g2_and2_1 _28735_ (.A(_00147_),
    .B(_15014_),
    .X(_15123_));
 sg13g2_and2_1 _28736_ (.A(_00158_),
    .B(_15123_),
    .X(_15124_));
 sg13g2_a22oi_1 _28737_ (.Y(_15125_),
    .B1(_15113_),
    .B2(net7377),
    .A2(_14748_),
    .A1(_08251_));
 sg13g2_o21ai_1 _28738_ (.B1(net6060),
    .Y(_15126_),
    .A1(net6430),
    .A2(_15124_));
 sg13g2_nand2_1 _28739_ (.Y(_15127_),
    .A(net6129),
    .B(_15123_));
 sg13g2_nand2_1 _28740_ (.Y(_15128_),
    .A(net6128),
    .B(_15124_));
 sg13g2_nand2_1 _28741_ (.Y(_15129_),
    .A(_13634_),
    .B(net6430));
 sg13g2_o21ai_1 _28742_ (.B1(_15129_),
    .Y(_15130_),
    .A1(_06388_),
    .A2(_15128_));
 sg13g2_a22oi_1 _28743_ (.Y(_15131_),
    .B1(_15130_),
    .B2(net6060),
    .A2(_15126_),
    .A1(_06388_));
 sg13g2_o21ai_1 _28744_ (.B1(_15125_),
    .Y(_15132_),
    .A1(net6980),
    .A2(_14748_));
 sg13g2_o21ai_1 _28745_ (.B1(net6410),
    .Y(_15133_),
    .A1(_15022_),
    .A2(_15094_));
 sg13g2_nand2_1 _28746_ (.Y(_15134_),
    .A(net6152),
    .B(net6418));
 sg13g2_o21ai_1 _28747_ (.B1(_15134_),
    .Y(_15135_),
    .A1(net6418),
    .A2(_15096_));
 sg13g2_a22oi_1 _28748_ (.Y(_15136_),
    .B1(_15135_),
    .B2(net6410),
    .A2(_15133_),
    .A1(_06391_));
 sg13g2_nand2_1 _28749_ (.Y(_15137_),
    .A(net6126),
    .B(_15093_));
 sg13g2_a21oi_1 _28750_ (.A1(net6414),
    .A2(_15137_),
    .Y(_15138_),
    .B1(_00167_));
 sg13g2_mux2_1 _28751_ (.A0(_15094_),
    .A1(_13471_),
    .S(_15022_),
    .X(_15139_));
 sg13g2_a21oi_1 _28752_ (.A1(net6410),
    .A2(_15139_),
    .Y(_15140_),
    .B1(_15138_));
 sg13g2_o21ai_1 _28753_ (.B1(net6414),
    .Y(_15141_),
    .A1(_15022_),
    .A2(_15092_));
 sg13g2_nand2_1 _28754_ (.Y(_15142_),
    .A(_13477_),
    .B(net6418));
 sg13g2_o21ai_1 _28755_ (.B1(_15142_),
    .Y(_15143_),
    .A1(net6418),
    .A2(_15093_));
 sg13g2_a22oi_1 _28756_ (.Y(_15144_),
    .B1(_15143_),
    .B2(net6414),
    .A2(_15141_),
    .A1(_06394_));
 sg13g2_nand2_1 _28757_ (.Y(_15145_),
    .A(_00163_),
    .B(_15090_));
 sg13g2_and3_1 _28758_ (.X(_15146_),
    .A(_00164_),
    .B(_00163_),
    .C(_15090_));
 sg13g2_o21ai_1 _28759_ (.B1(net6413),
    .Y(_15147_),
    .A1(net6417),
    .A2(_15146_));
 sg13g2_nand3_1 _28760_ (.B(net6126),
    .C(_15146_),
    .A(_00165_),
    .Y(_15148_));
 sg13g2_nand2_1 _28761_ (.Y(_15149_),
    .A(_13484_),
    .B(net6422));
 sg13g2_nand2_1 _28762_ (.Y(_15150_),
    .A(_15148_),
    .B(_15149_));
 sg13g2_a22oi_1 _28763_ (.Y(_15151_),
    .B1(_15150_),
    .B2(net6413),
    .A2(_15147_),
    .A1(_06399_));
 sg13g2_inv_1 _28764_ (.Y(_15152_),
    .A(_01718_));
 sg13g2_nand2_1 _28765_ (.Y(_15153_),
    .A(net6126),
    .B(_15145_));
 sg13g2_a21oi_1 _28766_ (.A1(net6413),
    .A2(_15153_),
    .Y(_15154_),
    .B1(_00164_));
 sg13g2_nand2_1 _28767_ (.Y(_15155_),
    .A(net6146),
    .B(net6422));
 sg13g2_mux2_1 _28768_ (.A0(_15146_),
    .A1(net6146),
    .S(net6417),
    .X(_15156_));
 sg13g2_a21oi_1 _28769_ (.A1(net6413),
    .A2(_15156_),
    .Y(_15157_),
    .B1(_15154_));
 sg13g2_o21ai_1 _28770_ (.B1(net6414),
    .Y(_15158_),
    .A1(net6417),
    .A2(_15090_));
 sg13g2_nand2_1 _28771_ (.Y(_15159_),
    .A(_13495_),
    .B(net6418));
 sg13g2_o21ai_1 _28772_ (.B1(_15159_),
    .Y(_15160_),
    .A1(net6423),
    .A2(_15145_));
 sg13g2_a22oi_1 _28773_ (.Y(_15161_),
    .B1(_15160_),
    .B2(net6414),
    .A2(_15158_),
    .A1(_06406_));
 sg13g2_mux4_1 _28774_ (.S0(net7795),
    .A0(_00795_),
    .A1(_00827_),
    .A2(_00859_),
    .A3(_00894_),
    .S1(net7738),
    .X(_15162_));
 sg13g2_nor2_1 _28775_ (.A(net7707),
    .B(_15162_),
    .Y(_15163_));
 sg13g2_o21ai_1 _28776_ (.B1(net6412),
    .Y(_15164_),
    .A1(net6417),
    .A2(_15088_));
 sg13g2_nand2_1 _28777_ (.Y(_15165_),
    .A(_13501_),
    .B(net6426));
 sg13g2_o21ai_1 _28778_ (.B1(_15165_),
    .Y(_15166_),
    .A1(net6426),
    .A2(_15091_));
 sg13g2_a22oi_1 _28779_ (.Y(_15167_),
    .B1(_15166_),
    .B2(net6412),
    .A2(_15164_),
    .A1(_06413_));
 sg13g2_nand2_1 _28780_ (.Y(_15168_),
    .A(net6125),
    .B(_15087_));
 sg13g2_a21oi_1 _28781_ (.A1(net6412),
    .A2(_15168_),
    .Y(_15169_),
    .B1(_00161_));
 sg13g2_nand2_1 _28782_ (.Y(_15170_),
    .A(net6142),
    .B(net6423));
 sg13g2_o21ai_1 _28783_ (.B1(_15170_),
    .Y(_15171_),
    .A1(net6426),
    .A2(_15089_));
 sg13g2_a21oi_1 _28784_ (.A1(net6412),
    .A2(_15171_),
    .Y(_15172_),
    .B1(_15169_));
 sg13g2_nand2_1 _28785_ (.Y(_15173_),
    .A(_00159_),
    .B(_15085_));
 sg13g2_nand2_1 _28786_ (.Y(_15174_),
    .A(net6125),
    .B(_15173_));
 sg13g2_a21oi_1 _28787_ (.A1(net6412),
    .A2(_15174_),
    .Y(_15175_),
    .B1(_00160_));
 sg13g2_nand4_1 _28788_ (.B(_00159_),
    .C(net6125),
    .A(_00160_),
    .Y(_15176_),
    .D(_15085_));
 sg13g2_nand2_1 _28789_ (.Y(_15177_),
    .A(_13511_),
    .B(net6426));
 sg13g2_nand2_1 _28790_ (.Y(_15178_),
    .A(_15176_),
    .B(_15177_));
 sg13g2_mux2_1 _28791_ (.A0(_01000_),
    .A1(_01035_),
    .S(net7794),
    .X(_15179_));
 sg13g2_a21oi_1 _28792_ (.A1(net6412),
    .A2(_15178_),
    .Y(_15180_),
    .B1(_15175_));
 sg13g2_o21ai_1 _28793_ (.B1(net6411),
    .Y(_15181_),
    .A1(net6417),
    .A2(_15085_));
 sg13g2_nand2_1 _28794_ (.Y(_15182_),
    .A(net6140),
    .B(net6426));
 sg13g2_o21ai_1 _28795_ (.B1(_15182_),
    .Y(_15183_),
    .A1(net6426),
    .A2(_15173_));
 sg13g2_a22oi_1 _28796_ (.Y(_15184_),
    .B1(_15183_),
    .B2(net6412),
    .A2(_15181_),
    .A1(_06433_));
 sg13g2_nor2_1 _28797_ (.A(_08522_),
    .B(_15179_),
    .Y(_15185_));
 sg13g2_o21ai_1 _28798_ (.B1(net6060),
    .Y(_15186_),
    .A1(net6430),
    .A2(_15123_));
 sg13g2_o21ai_1 _28799_ (.B1(_15128_),
    .Y(_15187_),
    .A1(_13646_),
    .A2(net6128));
 sg13g2_a22oi_1 _28800_ (.Y(_15188_),
    .B1(_15187_),
    .B2(net6060),
    .A2(_15186_),
    .A1(_06438_));
 sg13g2_o21ai_1 _28801_ (.B1(net6411),
    .Y(_15189_),
    .A1(net6417),
    .A2(_15083_));
 sg13g2_nand2_1 _28802_ (.Y(_15190_),
    .A(_13522_),
    .B(net6426));
 sg13g2_o21ai_1 _28803_ (.B1(_15190_),
    .Y(_15191_),
    .A1(net6425),
    .A2(_15086_));
 sg13g2_a22oi_1 _28804_ (.Y(_15192_),
    .B1(_15191_),
    .B2(net6411),
    .A2(_15189_),
    .A1(_06444_));
 sg13g2_o21ai_1 _28805_ (.B1(net6411),
    .Y(_15193_),
    .A1(net6417),
    .A2(_15081_));
 sg13g2_nand2_1 _28806_ (.Y(_15194_),
    .A(_13527_),
    .B(net6425));
 sg13g2_mux2_1 _28807_ (.A0(_00930_),
    .A1(_00965_),
    .S(net7794),
    .X(_15195_));
 sg13g2_o21ai_1 _28808_ (.B1(_15194_),
    .Y(_15196_),
    .A1(net6424),
    .A2(_15084_));
 sg13g2_a22oi_1 _28809_ (.Y(_15197_),
    .B1(_15196_),
    .B2(net6411),
    .A2(_15193_),
    .A1(_06449_));
 sg13g2_o21ai_1 _28810_ (.B1(net6411),
    .Y(_15198_),
    .A1(net6417),
    .A2(_15080_));
 sg13g2_nand2_1 _28811_ (.Y(_15199_),
    .A(_13532_),
    .B(net6424));
 sg13g2_o21ai_1 _28812_ (.B1(_15199_),
    .Y(_15200_),
    .A1(net6424),
    .A2(_15082_));
 sg13g2_a22oi_1 _28813_ (.Y(_15201_),
    .B1(_15200_),
    .B2(net6411),
    .A2(_15198_),
    .A1(_06454_));
 sg13g2_nand3_1 _28814_ (.B(_15065_),
    .C(_15077_),
    .A(_00153_),
    .Y(_15202_));
 sg13g2_nand2_1 _28815_ (.Y(_15203_),
    .A(net6127),
    .B(_15202_));
 sg13g2_a21oi_1 _28816_ (.A1(net6406),
    .A2(_15203_),
    .Y(_15204_),
    .B1(_00154_));
 sg13g2_nand2_1 _28817_ (.Y(_15205_),
    .A(_15021_),
    .B(_15077_));
 sg13g2_nand2_1 _28818_ (.Y(_15206_),
    .A(_13537_),
    .B(net6428));
 sg13g2_o21ai_1 _28819_ (.B1(net7694),
    .Y(_15207_),
    .A1(net7562),
    .A2(_15195_));
 sg13g2_o21ai_1 _28820_ (.B1(_15206_),
    .Y(_15208_),
    .A1(_15079_),
    .A2(_15205_));
 sg13g2_a21oi_1 _28821_ (.A1(net6406),
    .A2(_15208_),
    .Y(_15209_),
    .B1(_15204_));
 sg13g2_o21ai_1 _28822_ (.B1(net6127),
    .Y(_15210_),
    .A1(_15066_),
    .A2(net6748));
 sg13g2_a21oi_1 _28823_ (.A1(net6406),
    .A2(_15210_),
    .Y(_15211_),
    .B1(_00153_));
 sg13g2_nand3_1 _28824_ (.B(_15065_),
    .C(_15077_),
    .A(_00153_),
    .Y(_15212_));
 sg13g2_nand2_1 _28825_ (.Y(_15213_),
    .A(net6136),
    .B(net6427));
 sg13g2_o21ai_1 _28826_ (.B1(_15213_),
    .Y(_15214_),
    .A1(net6428),
    .A2(_15212_));
 sg13g2_a21oi_1 _28827_ (.A1(net6406),
    .A2(_15214_),
    .Y(_15215_),
    .B1(_15211_));
 sg13g2_or3_1 _28828_ (.A(_15163_),
    .B(_15185_),
    .C(_15207_),
    .X(_15216_));
 sg13g2_nor2_1 _28829_ (.A(_15064_),
    .B(net6748),
    .Y(_15217_));
 sg13g2_o21ai_1 _28830_ (.B1(net6406),
    .Y(_15218_),
    .A1(net6415),
    .A2(_15217_));
 sg13g2_nand2_1 _28831_ (.Y(_15219_),
    .A(_13547_),
    .B(net6429));
 sg13g2_o21ai_1 _28832_ (.B1(_15219_),
    .Y(_15220_),
    .A1(_15066_),
    .A2(_15205_));
 sg13g2_a22oi_1 _28833_ (.Y(_15221_),
    .B1(_15220_),
    .B2(net6406),
    .A2(_15218_),
    .A1(_06458_));
 sg13g2_mux2_1 _28834_ (.A0(_00635_),
    .A1(_00763_),
    .S(net7708),
    .X(_15222_));
 sg13g2_nand3_1 _28835_ (.B(_15062_),
    .C(_15077_),
    .A(_00150_),
    .Y(_15223_));
 sg13g2_nand2_1 _28836_ (.Y(_15224_),
    .A(net6127),
    .B(_15223_));
 sg13g2_a21oi_1 _28837_ (.A1(net6406),
    .A2(_15224_),
    .Y(_15225_),
    .B1(_00151_));
 sg13g2_nand2_1 _28838_ (.Y(_15226_),
    .A(_13553_),
    .B(net6427));
 sg13g2_o21ai_1 _28839_ (.B1(_15226_),
    .Y(_15227_),
    .A1(_15064_),
    .A2(_15205_));
 sg13g2_a21oi_1 _28840_ (.A1(net6406),
    .A2(_15227_),
    .Y(_15228_),
    .B1(_15225_));
 sg13g2_and2_1 _28841_ (.A(net7797),
    .B(_00939_),
    .X(_15229_));
 sg13g2_o21ai_1 _28842_ (.B1(net6128),
    .Y(_15230_),
    .A1(_15063_),
    .A2(net6748));
 sg13g2_a21oi_1 _28843_ (.A1(net6407),
    .A2(_15230_),
    .Y(_15231_),
    .B1(_00150_));
 sg13g2_nand3_1 _28844_ (.B(_15062_),
    .C(_15077_),
    .A(_00150_),
    .Y(_15232_));
 sg13g2_nand2_1 _28845_ (.Y(_15233_),
    .A(_13559_),
    .B(net6428));
 sg13g2_o21ai_1 _28846_ (.B1(_15233_),
    .Y(_15234_),
    .A1(net6428),
    .A2(_15232_));
 sg13g2_a21oi_1 _28847_ (.A1(net6407),
    .A2(_15234_),
    .Y(_15235_),
    .B1(_15231_));
 sg13g2_nor2b_1 _28848_ (.A(net7797),
    .B_N(_01291_),
    .Y(_15236_));
 sg13g2_o21ai_1 _28849_ (.B1(net6128),
    .Y(_15237_),
    .A1(_15061_),
    .A2(net6748));
 sg13g2_a21oi_1 _28850_ (.A1(net6407),
    .A2(_15237_),
    .Y(_15238_),
    .B1(_00149_));
 sg13g2_o21ai_1 _28851_ (.B1(_15026_),
    .Y(_15239_),
    .A1(_15063_),
    .A2(net6059));
 sg13g2_a21oi_1 _28852_ (.A1(net6407),
    .A2(_15239_),
    .Y(_15240_),
    .B1(_15238_));
 sg13g2_nor2_1 _28853_ (.A(_15059_),
    .B(net6748),
    .Y(_15241_));
 sg13g2_o21ai_1 _28854_ (.B1(net6407),
    .Y(_15242_),
    .A1(net6415),
    .A2(_15241_));
 sg13g2_o21ai_1 _28855_ (.B1(_15032_),
    .Y(_15243_),
    .A1(_15061_),
    .A2(net6059));
 sg13g2_a22oi_1 _28856_ (.Y(_15244_),
    .B1(_15243_),
    .B2(net6407),
    .A2(_15242_),
    .A1(_06466_));
 sg13g2_o21ai_1 _28857_ (.B1(net6060),
    .Y(_15245_),
    .A1(_15014_),
    .A2(net6430));
 sg13g2_nand2_1 _28858_ (.Y(_15246_),
    .A(_13656_),
    .B(_15020_));
 sg13g2_nand2_1 _28859_ (.Y(_15247_),
    .A(_15127_),
    .B(_15246_));
 sg13g2_a22oi_1 _28860_ (.Y(_15248_),
    .B1(_15247_),
    .B2(net6060),
    .A2(_15245_),
    .A1(_06472_));
 sg13g2_nor3_1 _28861_ (.A(_00112_),
    .B(_15058_),
    .C(net6059),
    .Y(_15249_));
 sg13g2_nor3_1 _28862_ (.A(_00146_),
    .B(_15010_),
    .C(_15249_),
    .Y(_15250_));
 sg13g2_mux2_1 _28863_ (.A0(_00667_),
    .A1(_00699_),
    .S(net7797),
    .X(_15251_));
 sg13g2_a221oi_1 _28864_ (.B2(_00146_),
    .C1(_15250_),
    .B1(_15249_),
    .A1(_13610_),
    .Y(_15252_),
    .A2(_15009_));
 sg13g2_o21ai_1 _28865_ (.B1(net6128),
    .Y(_15253_),
    .A1(_06489_),
    .A2(net6748));
 sg13g2_a21oi_1 _28866_ (.A1(net6408),
    .A2(_15253_),
    .Y(_15254_),
    .B1(_00145_));
 sg13g2_o21ai_1 _28867_ (.B1(_15044_),
    .Y(_15255_),
    .A1(_15058_),
    .A2(net6059));
 sg13g2_a21oi_1 _28868_ (.A1(net6408),
    .A2(_15255_),
    .Y(_15256_),
    .B1(_15254_));
 sg13g2_nor2b_1 _28869_ (.A(net7797),
    .B_N(_00731_),
    .Y(_15257_));
 sg13g2_o21ai_1 _28870_ (.B1(net6407),
    .Y(_15258_),
    .A1(net6415),
    .A2(_15077_));
 sg13g2_o21ai_1 _28871_ (.B1(_15129_),
    .Y(_15259_),
    .A1(_06489_),
    .A2(net6059));
 sg13g2_a22oi_1 _28872_ (.Y(_15260_),
    .B1(_15259_),
    .B2(net6408),
    .A2(_15258_),
    .A1(_06489_));
 sg13g2_o21ai_1 _28873_ (.B1(net6408),
    .Y(_15261_),
    .A1(net6416),
    .A2(_15076_));
 sg13g2_o21ai_1 _28874_ (.B1(net6059),
    .Y(_15262_),
    .A1(_13646_),
    .A2(net6129));
 sg13g2_a22oi_1 _28875_ (.Y(_15263_),
    .B1(_15262_),
    .B2(net6408),
    .A2(_15261_),
    .A1(_06495_));
 sg13g2_and2_1 _28876_ (.A(_15057_),
    .B(_15074_),
    .X(_15264_));
 sg13g2_and2_1 _28877_ (.A(_00141_),
    .B(_15264_),
    .X(_15265_));
 sg13g2_o21ai_1 _28878_ (.B1(net6409),
    .Y(_15266_),
    .A1(net6416),
    .A2(_15265_));
 sg13g2_nand2_1 _28879_ (.Y(_15267_),
    .A(net6130),
    .B(_15265_));
 sg13g2_o21ai_1 _28880_ (.B1(_15246_),
    .Y(_15268_),
    .A1(_06502_),
    .A2(_15267_));
 sg13g2_a22oi_1 _28881_ (.Y(_15269_),
    .B1(_15268_),
    .B2(net6409),
    .A2(_15266_),
    .A1(_06502_));
 sg13g2_o21ai_1 _28882_ (.B1(net6405),
    .Y(_15270_),
    .A1(net6416),
    .A2(_15264_));
 sg13g2_o21ai_1 _28883_ (.B1(_15267_),
    .Y(_15271_),
    .A1(_13703_),
    .A2(net6130));
 sg13g2_a22oi_1 _28884_ (.Y(_15272_),
    .B1(_15271_),
    .B2(net6409),
    .A2(_15270_),
    .A1(_06508_));
 sg13g2_and2_1 _28885_ (.A(_00133_),
    .B(_15074_),
    .X(_15273_));
 sg13g2_nand2_1 _28886_ (.Y(_15274_),
    .A(_00133_),
    .B(_15074_));
 sg13g2_nor2_1 _28887_ (.A(_15055_),
    .B(_15274_),
    .Y(_15275_));
 sg13g2_nand2_1 _28888_ (.Y(_15276_),
    .A(_00138_),
    .B(_15275_));
 sg13g2_and3_1 _28889_ (.X(_15277_),
    .A(_00139_),
    .B(_00138_),
    .C(_15275_));
 sg13g2_o21ai_1 _28890_ (.B1(net6405),
    .Y(_15278_),
    .A1(net6416),
    .A2(_15277_));
 sg13g2_nand2_1 _28891_ (.Y(_15279_),
    .A(net6130),
    .B(_15277_));
 sg13g2_nand2_1 _28892_ (.Y(_15280_),
    .A(net6454),
    .B(net6420));
 sg13g2_o21ai_1 _28893_ (.B1(_15280_),
    .Y(_15281_),
    .A1(_06512_),
    .A2(_15279_));
 sg13g2_a22oi_1 _28894_ (.Y(_15282_),
    .B1(_15281_),
    .B2(net6405),
    .A2(_15278_),
    .A1(_06512_));
 sg13g2_nand2_1 _28895_ (.Y(_15283_),
    .A(net6130),
    .B(_15276_));
 sg13g2_mux4_1 _28896_ (.S0(net7738),
    .A0(_15229_),
    .A1(_15236_),
    .A2(_15251_),
    .A3(_15257_),
    .S1(net7708),
    .X(_15284_));
 sg13g2_a21oi_1 _28897_ (.A1(net6405),
    .A2(_15283_),
    .Y(_15285_),
    .B1(_00139_));
 sg13g2_o21ai_1 _28898_ (.B1(_15279_),
    .Y(_15286_),
    .A1(_13873_),
    .A2(net6130));
 sg13g2_a21oi_1 _28899_ (.A1(net6405),
    .A2(_15286_),
    .Y(_15287_),
    .B1(_15285_));
 sg13g2_a221oi_1 _28900_ (.B2(net7531),
    .C1(net7690),
    .B1(_15284_),
    .A1(_08288_),
    .Y(_15288_),
    .A2(_15222_));
 sg13g2_o21ai_1 _28901_ (.B1(net6065),
    .Y(_15289_),
    .A1(net6420),
    .A2(_15275_));
 sg13g2_o21ai_1 _28902_ (.B1(_15103_),
    .Y(_15290_),
    .A1(net6420),
    .A2(_15276_));
 sg13g2_a22oi_1 _28903_ (.Y(_15291_),
    .B1(_15290_),
    .B2(net6065),
    .A2(_15289_),
    .A1(_06521_));
 sg13g2_nand2_1 _28904_ (.Y(_15292_),
    .A(_00134_),
    .B(_15273_));
 sg13g2_nand3_1 _28905_ (.B(_00134_),
    .C(_15273_),
    .A(_00135_),
    .Y(_15293_));
 sg13g2_nand2_1 _28906_ (.Y(_15294_),
    .A(_15021_),
    .B(_15293_));
 sg13g2_nor2_1 _28907_ (.A(net6419),
    .B(_15293_),
    .Y(_15295_));
 sg13g2_a22oi_1 _28908_ (.Y(_15296_),
    .B1(_15295_),
    .B2(_00137_),
    .A2(net6419),
    .A1(_13446_));
 sg13g2_inv_1 _28909_ (.Y(_15297_),
    .A(_15296_));
 sg13g2_a21oi_1 _28910_ (.A1(net6064),
    .A2(_15294_),
    .Y(_15298_),
    .B1(_00137_));
 sg13g2_a21oi_1 _28911_ (.A1(net6064),
    .A2(_15297_),
    .Y(_15299_),
    .B1(_15298_));
 sg13g2_o21ai_1 _28912_ (.B1(_15011_),
    .Y(_15300_),
    .A1(_15013_),
    .A2(net6430));
 sg13g2_nand2_1 _28913_ (.Y(_15301_),
    .A(_15014_),
    .B(net6129));
 sg13g2_o21ai_1 _28914_ (.B1(_15301_),
    .Y(_15302_),
    .A1(_13703_),
    .A2(net6129));
 sg13g2_a22oi_1 _28915_ (.Y(_15303_),
    .B1(_15302_),
    .B2(_15011_),
    .A2(_15300_),
    .A1(_06527_));
 sg13g2_nand2_1 _28916_ (.Y(_15304_),
    .A(_15021_),
    .B(_15292_));
 sg13g2_a21oi_1 _28917_ (.A1(net6064),
    .A2(_15304_),
    .Y(_15305_),
    .B1(_00135_));
 sg13g2_o21ai_1 _28918_ (.B1(_15115_),
    .Y(_15306_),
    .A1(net6419),
    .A2(_15293_));
 sg13g2_a21oi_1 _28919_ (.A1(net6064),
    .A2(_15306_),
    .Y(_15307_),
    .B1(_15305_));
 sg13g2_mux2_1 _28920_ (.A0(_01422_),
    .A1(_01458_),
    .S(net7795),
    .X(_15308_));
 sg13g2_o21ai_1 _28921_ (.B1(net6064),
    .Y(_15309_),
    .A1(net6418),
    .A2(_15273_));
 sg13g2_o21ai_1 _28922_ (.B1(_15120_),
    .Y(_15310_),
    .A1(net6418),
    .A2(_15292_));
 sg13g2_nor3_1 _28923_ (.A(net7573),
    .B(net7571),
    .C(_15308_),
    .Y(_15311_));
 sg13g2_a22oi_1 _28924_ (.Y(_15312_),
    .B1(_15310_),
    .B2(net6064),
    .A2(_15309_),
    .A1(_06532_));
 sg13g2_o21ai_1 _28925_ (.B1(net6064),
    .Y(_15313_),
    .A1(net6423),
    .A2(_15074_));
 sg13g2_o21ai_1 _28926_ (.B1(_15134_),
    .Y(_15314_),
    .A1(net6423),
    .A2(_15274_));
 sg13g2_a22oi_1 _28927_ (.Y(_15315_),
    .B1(_15314_),
    .B2(net6064),
    .A2(_15313_),
    .A1(_06535_));
 sg13g2_nand2_1 _28928_ (.Y(_15316_),
    .A(_00124_),
    .B(_15073_));
 sg13g2_and3_1 _28929_ (.X(_15317_),
    .A(_00126_),
    .B(_00124_),
    .C(_15073_));
 sg13g2_nand3_1 _28930_ (.B(_00124_),
    .C(_15073_),
    .A(_00126_),
    .Y(_15318_));
 sg13g2_nor2_1 _28931_ (.A(_06556_),
    .B(_15318_),
    .Y(_15319_));
 sg13g2_nand2_1 _28932_ (.Y(_15320_),
    .A(_00127_),
    .B(_15317_));
 sg13g2_nor2_1 _28933_ (.A(_06552_),
    .B(_15320_),
    .Y(_15321_));
 sg13g2_nand2_1 _28934_ (.Y(_15322_),
    .A(_00128_),
    .B(_15319_));
 sg13g2_nand2_1 _28935_ (.Y(_15323_),
    .A(_00129_),
    .B(_15321_));
 sg13g2_and3_1 _28936_ (.X(_15324_),
    .A(_00130_),
    .B(_00129_),
    .C(_15321_));
 sg13g2_nand2_1 _28937_ (.Y(_15325_),
    .A(_00131_),
    .B(_15324_));
 sg13g2_nand2_1 _28938_ (.Y(_15326_),
    .A(net6126),
    .B(_15325_));
 sg13g2_a21oi_1 _28939_ (.A1(net6067),
    .A2(_15326_),
    .Y(_15327_),
    .B1(_00132_));
 sg13g2_nor2_1 _28940_ (.A(net6422),
    .B(_15325_),
    .Y(_15328_));
 sg13g2_a22oi_1 _28941_ (.Y(_15329_),
    .B1(_15328_),
    .B2(_00132_),
    .A2(net6422),
    .A1(_13471_));
 sg13g2_inv_1 _28942_ (.Y(_15330_),
    .A(_15329_));
 sg13g2_mux2_1 _28943_ (.A0(_01493_),
    .A1(_01528_),
    .S(net7795),
    .X(_15331_));
 sg13g2_a21oi_1 _28944_ (.A1(net6067),
    .A2(_15330_),
    .Y(_15332_),
    .B1(_15327_));
 sg13g2_nor3_1 _28945_ (.A(net7573),
    .B(net7562),
    .C(_15331_),
    .Y(_15333_));
 sg13g2_o21ai_1 _28946_ (.B1(net6067),
    .Y(_15334_),
    .A1(net6422),
    .A2(_15324_));
 sg13g2_o21ai_1 _28947_ (.B1(_15142_),
    .Y(_15335_),
    .A1(net6422),
    .A2(_15325_));
 sg13g2_a22oi_1 _28948_ (.Y(_15336_),
    .B1(_15335_),
    .B2(net6067),
    .A2(_15334_),
    .A1(_06542_));
 sg13g2_nand2_1 _28949_ (.Y(_15337_),
    .A(net6126),
    .B(_15323_));
 sg13g2_a21oi_1 _28950_ (.A1(net6067),
    .A2(_15337_),
    .Y(_15338_),
    .B1(_00130_));
 sg13g2_nand2_1 _28951_ (.Y(_15339_),
    .A(net6126),
    .B(_15324_));
 sg13g2_a21oi_1 _28952_ (.A1(_15149_),
    .A2(_15339_),
    .Y(_15340_),
    .B1(_15012_));
 sg13g2_nor2_1 _28953_ (.A(_15338_),
    .B(_15340_),
    .Y(_15341_));
 sg13g2_o21ai_1 _28954_ (.B1(net6067),
    .Y(_15342_),
    .A1(net6421),
    .A2(_15321_));
 sg13g2_o21ai_1 _28955_ (.B1(_15155_),
    .Y(_15343_),
    .A1(net6421),
    .A2(_15323_));
 sg13g2_a22oi_1 _28956_ (.Y(_15344_),
    .B1(_15343_),
    .B2(net6067),
    .A2(_15342_),
    .A1(_06548_));
 sg13g2_o21ai_1 _28957_ (.B1(net6066),
    .Y(_15345_),
    .A1(net6421),
    .A2(_15319_));
 sg13g2_mux2_1 _28958_ (.A0(_01352_),
    .A1(_01387_),
    .S(net7793),
    .X(_15346_));
 sg13g2_o21ai_1 _28959_ (.B1(_15159_),
    .Y(_15347_),
    .A1(net6422),
    .A2(_15322_));
 sg13g2_nor3_1 _28960_ (.A(net7573),
    .B(net7558),
    .C(_15346_),
    .Y(_15348_));
 sg13g2_a22oi_1 _28961_ (.Y(_15349_),
    .B1(_15347_),
    .B2(net6066),
    .A2(_15345_),
    .A1(_06552_));
 sg13g2_o21ai_1 _28962_ (.B1(net6066),
    .Y(_15350_),
    .A1(net6421),
    .A2(_15317_));
 sg13g2_o21ai_1 _28963_ (.B1(_15165_),
    .Y(_15351_),
    .A1(net6421),
    .A2(_15320_));
 sg13g2_a22oi_1 _28964_ (.Y(_15352_),
    .B1(_15351_),
    .B2(net6066),
    .A2(_15350_),
    .A1(_06556_));
 sg13g2_nand2_1 _28965_ (.Y(_15353_),
    .A(net6125),
    .B(_15316_));
 sg13g2_a21oi_1 _28966_ (.A1(net6066),
    .A2(_15353_),
    .Y(_15354_),
    .B1(_00126_));
 sg13g2_o21ai_1 _28967_ (.B1(_15170_),
    .Y(_15355_),
    .A1(net6421),
    .A2(_15318_));
 sg13g2_a21oi_1 _28968_ (.A1(net6066),
    .A2(_15355_),
    .Y(_15356_),
    .B1(_15354_));
 sg13g2_o21ai_1 _28969_ (.B1(net6065),
    .Y(_15357_),
    .A1(_00114_),
    .A2(net6420));
 sg13g2_mux2_1 _28970_ (.A0(_15013_),
    .A1(net6454),
    .S(net6416),
    .X(_15358_));
 sg13g2_mux2_1 _28971_ (.A0(_01563_),
    .A1(_01598_),
    .S(net7793),
    .X(_15359_));
 sg13g2_a22oi_1 _28972_ (.Y(_15360_),
    .B1(_15358_),
    .B2(net6065),
    .A2(_15357_),
    .A1(_06569_));
 sg13g2_o21ai_1 _28973_ (.B1(net6066),
    .Y(_15361_),
    .A1(net6421),
    .A2(_15073_));
 sg13g2_nor2_1 _28974_ (.A(net7556),
    .B(_15359_),
    .Y(_15362_));
 sg13g2_o21ai_1 _28975_ (.B1(_15177_),
    .Y(_15363_),
    .A1(net6421),
    .A2(_15316_));
 sg13g2_a22oi_1 _28976_ (.Y(_15364_),
    .B1(_15363_),
    .B2(net6066),
    .A2(_15361_),
    .A1(_06574_));
 sg13g2_nand2_1 _28977_ (.Y(_15365_),
    .A(_00121_),
    .B(_15070_));
 sg13g2_nand3_1 _28978_ (.B(_00121_),
    .C(_15070_),
    .A(_00122_),
    .Y(_15366_));
 sg13g2_nand2_1 _28979_ (.Y(_15367_),
    .A(net6125),
    .B(_15366_));
 sg13g2_or4_1 _28980_ (.A(_15311_),
    .B(_15333_),
    .C(_15348_),
    .D(_15362_),
    .X(_15368_));
 sg13g2_a21oi_1 _28981_ (.A1(net6062),
    .A2(_15367_),
    .Y(_15369_),
    .B1(_00123_));
 sg13g2_nor2_1 _28982_ (.A(net6425),
    .B(_15366_),
    .Y(_15370_));
 sg13g2_a22oi_1 _28983_ (.Y(_15371_),
    .B1(_15370_),
    .B2(_00123_),
    .A2(net6425),
    .A1(net6140));
 sg13g2_inv_1 _28984_ (.Y(_15372_),
    .A(_15371_));
 sg13g2_a21oi_1 _28985_ (.A1(net6062),
    .A2(_15372_),
    .Y(_15373_),
    .B1(_15369_));
 sg13g2_nand2_1 _28986_ (.Y(_15374_),
    .A(net6125),
    .B(_15365_));
 sg13g2_a21oi_1 _28987_ (.A1(net6063),
    .A2(_15374_),
    .Y(_15375_),
    .B1(_00122_));
 sg13g2_o21ai_1 _28988_ (.B1(_15190_),
    .Y(_15376_),
    .A1(net6425),
    .A2(_15366_));
 sg13g2_a21oi_1 _28989_ (.A1(net6063),
    .A2(_15376_),
    .Y(_15377_),
    .B1(_15375_));
 sg13g2_o21ai_1 _28990_ (.B1(net6062),
    .Y(_15378_),
    .A1(net6425),
    .A2(_15070_));
 sg13g2_o21ai_1 _28991_ (.B1(_15194_),
    .Y(_15379_),
    .A1(net6425),
    .A2(_15365_));
 sg13g2_mux2_1 _28992_ (.A0(_01141_),
    .A1(_01176_),
    .S(net7791),
    .X(_15380_));
 sg13g2_a22oi_1 _28993_ (.Y(_15381_),
    .B1(_15379_),
    .B2(net6062),
    .A2(_15378_),
    .A1(_06585_));
 sg13g2_nand2_1 _28994_ (.Y(_15382_),
    .A(net6125),
    .B(_15069_));
 sg13g2_a21oi_1 _28995_ (.A1(net6062),
    .A2(_15382_),
    .Y(_15383_),
    .B1(_00120_));
 sg13g2_o21ai_1 _28996_ (.B1(_15199_),
    .Y(_15384_),
    .A1(net6424),
    .A2(_15071_));
 sg13g2_a21oi_1 _28997_ (.A1(net6062),
    .A2(_15384_),
    .Y(_15385_),
    .B1(_15383_));
 sg13g2_o21ai_1 _28998_ (.B1(net6062),
    .Y(_15386_),
    .A1(net6424),
    .A2(_15068_));
 sg13g2_o21ai_1 _28999_ (.B1(_15206_),
    .Y(_15387_),
    .A1(net6424),
    .A2(_15069_));
 sg13g2_a22oi_1 _29000_ (.Y(_15388_),
    .B1(_15387_),
    .B2(net6062),
    .A2(_15386_),
    .A1(_06592_));
 sg13g2_nor2_1 _29001_ (.A(_15017_),
    .B(_15050_),
    .Y(_15389_));
 sg13g2_o21ai_1 _29002_ (.B1(net6063),
    .Y(_15390_),
    .A1(net6427),
    .A2(_15389_));
 sg13g2_nand3_1 _29003_ (.B(net6127),
    .C(_15389_),
    .A(_00118_),
    .Y(_15391_));
 sg13g2_a21oi_1 _29004_ (.A1(_15213_),
    .A2(_15391_),
    .Y(_15392_),
    .B1(_15012_));
 sg13g2_mux2_1 _29005_ (.A0(_01070_),
    .A1(_01106_),
    .S(net7791),
    .X(_15393_));
 sg13g2_a21oi_1 _29006_ (.A1(_06597_),
    .A2(_15390_),
    .Y(_15394_),
    .B1(_15392_));
 sg13g2_and3_1 _29007_ (.X(_15395_),
    .A(_00177_),
    .B(_00115_),
    .C(_15018_));
 sg13g2_nand2_1 _29008_ (.Y(_15396_),
    .A(_00116_),
    .B(_15395_));
 sg13g2_nand2_1 _29009_ (.Y(_15397_),
    .A(net6127),
    .B(_15396_));
 sg13g2_a21oi_1 _29010_ (.A1(net6061),
    .A2(_15397_),
    .Y(_15398_),
    .B1(_00117_));
 sg13g2_nor2_1 _29011_ (.A(net6427),
    .B(_15396_),
    .Y(_15399_));
 sg13g2_a22oi_1 _29012_ (.Y(_15400_),
    .B1(_15399_),
    .B2(_00117_),
    .A2(net6427),
    .A1(_13547_));
 sg13g2_inv_1 _29013_ (.Y(_15401_),
    .A(_15400_));
 sg13g2_a21oi_1 _29014_ (.A1(net6061),
    .A2(_15401_),
    .Y(_15402_),
    .B1(_15398_));
 sg13g2_o21ai_1 _29015_ (.B1(net6061),
    .Y(_15403_),
    .A1(net6427),
    .A2(_15395_));
 sg13g2_o21ai_1 _29016_ (.B1(_15226_),
    .Y(_15404_),
    .A1(net6427),
    .A2(_15396_));
 sg13g2_a22oi_1 _29017_ (.Y(_15405_),
    .B1(_15404_),
    .B2(net6061),
    .A2(_15403_),
    .A1(_06607_));
 sg13g2_nand2_1 _29018_ (.Y(_15406_),
    .A(net6127),
    .B(_15025_));
 sg13g2_a21oi_1 _29019_ (.A1(net6061),
    .A2(_15406_),
    .Y(_15407_),
    .B1(_00115_));
 sg13g2_nand2_1 _29020_ (.Y(_15408_),
    .A(net6127),
    .B(_15395_));
 sg13g2_a21oi_1 _29021_ (.A1(_15233_),
    .A2(_15408_),
    .Y(_15409_),
    .B1(_15012_));
 sg13g2_nor2_1 _29022_ (.A(_15407_),
    .B(_15409_),
    .Y(_15410_));
 sg13g2_o21ai_1 _29023_ (.B1(net6065),
    .Y(_15411_),
    .A1(_13873_),
    .A2(net6130));
 sg13g2_a21oi_1 _29024_ (.A1(_13873_),
    .A2(net6420),
    .Y(_15412_),
    .B1(_06615_));
 sg13g2_mux2_1 _29025_ (.A0(_01282_),
    .A1(_01317_),
    .S(net7791),
    .X(_15413_));
 sg13g2_a22oi_1 _29026_ (.Y(_15414_),
    .B1(_15412_),
    .B2(net6065),
    .A2(_15411_),
    .A1(_06615_));
 sg13g2_nand2_1 _29027_ (.Y(_15415_),
    .A(_09555_),
    .B(_13423_));
 sg13g2_mux2_1 _29028_ (.A0(net6131),
    .A1(_00113_),
    .S(_15415_),
    .X(_15416_));
 sg13g2_nor2_1 _29029_ (.A(_13873_),
    .B(_15415_),
    .Y(_15417_));
 sg13g2_a21oi_1 _29030_ (.A1(_06628_),
    .A2(_15415_),
    .Y(_15418_),
    .B1(_15417_));
 sg13g2_or2_1 _29031_ (.X(_15419_),
    .B(core_busy_q),
    .A(net349));
 sg13g2_o21ai_1 _29032_ (.B1(fetch_enable_q),
    .Y(net439),
    .A1(_07002_),
    .A2(_15419_));
 sg13g2_nand2b_1 _29033_ (.Y(_15420_),
    .B(net439),
    .A_N(net438));
 sg13g2_nor2_1 _29034_ (.A(_01839_),
    .B(net7937),
    .Y(_15421_));
 sg13g2_and2_1 _29035_ (.A(_06910_),
    .B(_15421_),
    .X(_15422_));
 sg13g2_nand4_1 _29036_ (.B(_07668_),
    .C(_09355_),
    .A(_06959_),
    .Y(_15423_),
    .D(_15422_));
 sg13g2_nand2_1 _29037_ (.Y(_15424_),
    .A(\load_store_unit_i.handle_misaligned_q ),
    .B(_06684_));
 sg13g2_nor3_1 _29038_ (.A(_05957_),
    .B(_06657_),
    .C(_06659_),
    .Y(_15425_));
 sg13g2_a21oi_1 _29039_ (.A1(_06659_),
    .A2(_15424_),
    .Y(net470),
    .B1(_15425_));
 sg13g2_o21ai_1 _29040_ (.B1(_15424_),
    .Y(_15426_),
    .A1(net6747),
    .A2(_06684_));
 sg13g2_nand3_1 _29041_ (.B(net6726),
    .C(_06658_),
    .A(\load_store_unit_i.handle_misaligned_q ),
    .Y(_15427_));
 sg13g2_o21ai_1 _29042_ (.B1(_15427_),
    .Y(net471),
    .A1(net6726),
    .A2(_15426_));
 sg13g2_nand3_1 _29043_ (.B(net6747),
    .C(net6726),
    .A(\load_store_unit_i.handle_misaligned_q ),
    .Y(_15428_));
 sg13g2_o21ai_1 _29044_ (.B1(_15428_),
    .Y(_15429_),
    .A1(\load_store_unit_i.handle_misaligned_q ),
    .A2(net6726));
 sg13g2_nand2_1 _29045_ (.Y(_15430_),
    .A(_07026_),
    .B(net6727));
 sg13g2_nand2_1 _29046_ (.Y(_15431_),
    .A(_01889_),
    .B(net6747));
 sg13g2_o21ai_1 _29047_ (.B1(_15430_),
    .Y(_15432_),
    .A1(net6726),
    .A2(_15431_));
 sg13g2_mux2_1 _29048_ (.A0(_01211_),
    .A1(_01246_),
    .S(net7791),
    .X(_15433_));
 sg13g2_a22oi_1 _29049_ (.Y(_15434_),
    .B1(_15432_),
    .B2(_05957_),
    .A2(_15429_),
    .A1(_06658_));
 sg13g2_o21ai_1 _29050_ (.B1(_15434_),
    .Y(net472),
    .A1(_06684_),
    .A2(_15430_));
 sg13g2_a21oi_1 _29051_ (.A1(_01889_),
    .A2(net6726),
    .Y(_15435_),
    .B1(_06658_));
 sg13g2_nand3_1 _29052_ (.B(net6726),
    .C(_06683_),
    .A(net6746),
    .Y(_15436_));
 sg13g2_o21ai_1 _29053_ (.B1(_15436_),
    .Y(net473),
    .A1(\load_store_unit_i.handle_misaligned_q ),
    .A2(_15435_));
 sg13g2_a21oi_1 _29054_ (.A1(_08627_),
    .A2(_06644_),
    .Y(net474),
    .B1(net7657));
 sg13g2_mux2_1 _29055_ (.A0(_03122_),
    .A1(net7271),
    .S(net6718),
    .X(_15437_));
 sg13g2_and2_1 _29056_ (.A(net6744),
    .B(_15437_),
    .X(_15438_));
 sg13g2_nor2_1 _29057_ (.A(net7103),
    .B(net6718),
    .Y(_15439_));
 sg13g2_a21oi_1 _29058_ (.A1(_02584_),
    .A2(net6718),
    .Y(_15440_),
    .B1(_15439_));
 sg13g2_a21oi_1 _29059_ (.A1(net6732),
    .A2(_15440_),
    .Y(net475),
    .B1(_15438_));
 sg13g2_nor2_1 _29060_ (.A(_03192_),
    .B(net6721),
    .Y(_15441_));
 sg13g2_a21oi_1 _29061_ (.A1(net7270),
    .A2(net6721),
    .Y(_15442_),
    .B1(_15441_));
 sg13g2_and2_1 _29062_ (.A(net6745),
    .B(_15442_),
    .X(_15443_));
 sg13g2_nor2_1 _29063_ (.A(net7077),
    .B(net6720),
    .Y(_15444_));
 sg13g2_a21oi_1 _29064_ (.A1(net7345),
    .A2(net6720),
    .Y(_15445_),
    .B1(_15444_));
 sg13g2_a21oi_1 _29065_ (.A1(net6733),
    .A2(_15445_),
    .Y(net486),
    .B1(_15443_));
 sg13g2_mux4_1 _29066_ (.S0(net7516),
    .A0(_15380_),
    .A1(_15393_),
    .A2(_15413_),
    .A3(_15433_),
    .S1(net7709),
    .X(_15446_));
 sg13g2_inv_1 _29067_ (.Y(_15447_),
    .A(_15446_));
 sg13g2_mux4_1 _29068_ (.S0(net6727),
    .A0(_10750_),
    .A1(_02713_),
    .A2(_03256_),
    .A3(_02171_),
    .S1(net6746),
    .X(net497));
 sg13g2_mux2_1 _29069_ (.A0(_03327_),
    .A1(_02252_),
    .S(net6719),
    .X(_15448_));
 sg13g2_mux2_1 _29070_ (.A0(_11665_),
    .A1(_02778_),
    .S(net6719),
    .X(_15449_));
 sg13g2_mux2_1 _29071_ (.A0(_15448_),
    .A1(_15449_),
    .S(net6732),
    .X(net500));
 sg13g2_nor2_1 _29072_ (.A(net7260),
    .B(net6723),
    .Y(_15450_));
 sg13g2_a21oi_1 _29073_ (.A1(_02324_),
    .A2(net6723),
    .Y(_15451_),
    .B1(_15450_));
 sg13g2_and2_1 _29074_ (.A(net6742),
    .B(_15451_),
    .X(_15452_));
 sg13g2_nor2_1 _29075_ (.A(_12791_),
    .B(net6722),
    .Y(_15453_));
 sg13g2_a21oi_1 _29076_ (.A1(_02850_),
    .A2(net6722),
    .Y(_15454_),
    .B1(_15453_));
 sg13g2_a21o_1 _29077_ (.A2(_15447_),
    .A1(net7592),
    .B1(_15368_),
    .X(_15455_));
 sg13g2_a21oi_1 _29078_ (.A1(net6734),
    .A2(_15454_),
    .Y(net501),
    .B1(_15452_));
 sg13g2_nor2_1 _29079_ (.A(_03473_),
    .B(net6722),
    .Y(_15456_));
 sg13g2_a21oi_1 _29080_ (.A1(_02399_),
    .A2(net6723),
    .Y(_15457_),
    .B1(_15456_));
 sg13g2_a221oi_1 _29081_ (.B2(net7592),
    .C1(_15368_),
    .B1(_15447_),
    .A1(_15216_),
    .Y(_15458_),
    .A2(_15288_));
 sg13g2_and2_1 _29082_ (.A(net6742),
    .B(_15457_),
    .X(_15459_));
 sg13g2_nor2_1 _29083_ (.A(net7074),
    .B(net6722),
    .Y(_15460_));
 sg13g2_a21oi_1 _29084_ (.A1(_02918_),
    .A2(net6723),
    .Y(_15461_),
    .B1(_15460_));
 sg13g2_a21o_1 _29085_ (.A2(_15288_),
    .A1(_15216_),
    .B1(_15455_),
    .X(_15462_));
 sg13g2_a21oi_1 _29086_ (.A1(net6734),
    .A2(_15461_),
    .Y(net502),
    .B1(_15459_));
 sg13g2_nor2_1 _29087_ (.A(net7259),
    .B(net6721),
    .Y(_15463_));
 sg13g2_a21oi_1 _29088_ (.A1(_02475_),
    .A2(net6721),
    .Y(_15464_),
    .B1(_15463_));
 sg13g2_and2_1 _29089_ (.A(net6745),
    .B(_15464_),
    .X(_15465_));
 sg13g2_nor2_1 _29090_ (.A(net7291),
    .B(_15462_),
    .Y(_15466_));
 sg13g2_nor2_1 _29091_ (.A(_14725_),
    .B(net6721),
    .Y(_15467_));
 sg13g2_a21oi_1 _29092_ (.A1(net7339),
    .A2(net6721),
    .Y(_15468_),
    .B1(_15467_));
 sg13g2_a21oi_1 _29093_ (.A1(net6733),
    .A2(_15468_),
    .Y(net503),
    .B1(_15465_));
 sg13g2_mux2_1 _29094_ (.A0(_03608_),
    .A1(net7264),
    .S(net6724),
    .X(_15469_));
 sg13g2_and2_1 _29095_ (.A(net6743),
    .B(_15469_),
    .X(_15470_));
 sg13g2_nor2_1 _29096_ (.A(_15462_),
    .B(net6724),
    .Y(_15471_));
 sg13g2_a21oi_1 _29097_ (.A1(net7337),
    .A2(net6724),
    .Y(_15472_),
    .B1(_15471_));
 sg13g2_a21oi_1 _29098_ (.A1(net6735),
    .A2(_15472_),
    .Y(net504),
    .B1(_15470_));
 sg13g2_nor2_1 _29099_ (.A(net7271),
    .B(net6720),
    .Y(_15473_));
 sg13g2_a21oi_1 _29100_ (.A1(net7335),
    .A2(net6719),
    .Y(_15474_),
    .B1(_15473_));
 sg13g2_and2_1 _29101_ (.A(net6732),
    .B(_15474_),
    .X(_15475_));
 sg13g2_a21oi_1 _29102_ (.A1(net6744),
    .A2(_15440_),
    .Y(net505),
    .B1(_15475_));
 sg13g2_and2_1 _29103_ (.A(_03191_),
    .B(net6720),
    .X(_15476_));
 sg13g2_nor2_1 _29104_ (.A(_02104_),
    .B(net6717),
    .Y(_15477_));
 sg13g2_nor3_1 _29105_ (.A(net6747),
    .B(_15476_),
    .C(_15477_),
    .Y(_15478_));
 sg13g2_a21oi_1 _29106_ (.A1(net6745),
    .A2(_15445_),
    .Y(net506),
    .B1(_15478_));
 sg13g2_mux4_1 _29107_ (.S0(net6727),
    .A0(_02171_),
    .A1(_03256_),
    .A2(_10750_),
    .A3(_02713_),
    .S1(net6746),
    .X(net476));
 sg13g2_nor2_1 _29108_ (.A(net6732),
    .B(_15449_),
    .Y(_15479_));
 sg13g2_nor2_1 _29109_ (.A(net7269),
    .B(net6719),
    .Y(_15480_));
 sg13g2_a21oi_1 _29110_ (.A1(_03327_),
    .A2(net6719),
    .Y(_15481_),
    .B1(_15480_));
 sg13g2_a21oi_1 _29111_ (.A1(net6732),
    .A2(_15481_),
    .Y(net477),
    .B1(_15479_));
 sg13g2_and2_1 _29112_ (.A(net6742),
    .B(_15454_),
    .X(_15482_));
 sg13g2_nor2_1 _29113_ (.A(net7266),
    .B(net6723),
    .Y(_15483_));
 sg13g2_a21oi_1 _29114_ (.A1(_03403_),
    .A2(net6723),
    .Y(_15484_),
    .B1(_15483_));
 sg13g2_a21oi_1 _29115_ (.A1(net6734),
    .A2(_15484_),
    .Y(net478),
    .B1(_15482_));
 sg13g2_nor2_1 _29116_ (.A(net7265),
    .B(net6724),
    .Y(_15485_));
 sg13g2_a21oi_1 _29117_ (.A1(net7330),
    .A2(net6724),
    .Y(_15486_),
    .B1(_15485_));
 sg13g2_and2_1 _29118_ (.A(net6734),
    .B(_15486_),
    .X(_15487_));
 sg13g2_a21oi_1 _29119_ (.A1(net6742),
    .A2(_15461_),
    .Y(net479),
    .B1(_15487_));
 sg13g2_nor2_1 _29120_ (.A(_02476_),
    .B(net6725),
    .Y(_15488_));
 sg13g2_a21oi_1 _29121_ (.A1(_03537_),
    .A2(net6725),
    .Y(_15489_),
    .B1(_15488_));
 sg13g2_and2_1 _29122_ (.A(net6733),
    .B(_15489_),
    .X(_15490_));
 sg13g2_a21oi_1 _29123_ (.A1(net6745),
    .A2(_15468_),
    .Y(net480),
    .B1(_15490_));
 sg13g2_mux2_1 _29124_ (.A0(net7264),
    .A1(_03608_),
    .S(net6724),
    .X(_15491_));
 sg13g2_inv_1 _29125_ (.Y(_15492_),
    .A(_01704_));
 sg13g2_and2_1 _29126_ (.A(net6735),
    .B(_15491_),
    .X(_15493_));
 sg13g2_a21oi_1 _29127_ (.A1(net6742),
    .A2(_15472_),
    .Y(net481),
    .B1(_15493_));
 sg13g2_mux2_1 _29128_ (.A0(_02585_),
    .A1(net7103),
    .S(net6718),
    .X(_15494_));
 sg13g2_and2_1 _29129_ (.A(net6732),
    .B(_15494_),
    .X(_15495_));
 sg13g2_a21oi_1 _29130_ (.A1(net6744),
    .A2(_15474_),
    .Y(net482),
    .B1(_15495_));
 sg13g2_nor3_1 _29131_ (.A(_07026_),
    .B(_15476_),
    .C(_15477_),
    .Y(_15496_));
 sg13g2_mux2_1 _29132_ (.A0(_02652_),
    .A1(net7077),
    .S(net6720),
    .X(_15497_));
 sg13g2_a21oi_1 _29133_ (.A1(net6733),
    .A2(_15497_),
    .Y(net483),
    .B1(_15496_));
 sg13g2_mux4_1 _29134_ (.S0(net6746),
    .A0(_02713_),
    .A1(_02171_),
    .A2(_10750_),
    .A3(_03256_),
    .S1(net6727),
    .X(net484));
 sg13g2_nand2_1 _29135_ (.Y(_15498_),
    .A(_11665_),
    .B(net6719));
 sg13g2_o21ai_1 _29136_ (.B1(_15498_),
    .Y(_15499_),
    .A1(_02779_),
    .A2(net6719));
 sg13g2_nor2_1 _29137_ (.A(net6744),
    .B(_15499_),
    .Y(_15500_));
 sg13g2_a21oi_1 _29138_ (.A1(net6744),
    .A2(_15481_),
    .Y(net485),
    .B1(_15500_));
 sg13g2_and2_1 _29139_ (.A(net6742),
    .B(_15484_),
    .X(_15501_));
 sg13g2_nor2_1 _29140_ (.A(net7261),
    .B(net6722),
    .Y(_15502_));
 sg13g2_a21oi_1 _29141_ (.A1(net7281),
    .A2(net6722),
    .Y(_15503_),
    .B1(_15502_));
 sg13g2_a21oi_1 _29142_ (.A1(net6734),
    .A2(_15503_),
    .Y(net487),
    .B1(_15501_));
 sg13g2_mux2_1 _29143_ (.A0(_02919_),
    .A1(net7074),
    .S(\alu_adder_result_ex[1] ),
    .X(_15504_));
 sg13g2_and2_1 _29144_ (.A(_07026_),
    .B(_15504_),
    .X(_15505_));
 sg13g2_a21oi_1 _29145_ (.A1(net6743),
    .A2(_15486_),
    .Y(net488),
    .B1(_15505_));
 sg13g2_and2_1 _29146_ (.A(net6745),
    .B(_15489_),
    .X(_15506_));
 sg13g2_nor2_1 _29147_ (.A(_02986_),
    .B(net6721),
    .Y(_15507_));
 sg13g2_a21oi_1 _29148_ (.A1(net7274),
    .A2(net6721),
    .Y(_15508_),
    .B1(_15507_));
 sg13g2_a21oi_1 _29149_ (.A1(net6733),
    .A2(_15508_),
    .Y(net489),
    .B1(_15506_));
 sg13g2_and2_1 _29150_ (.A(net6743),
    .B(_15491_),
    .X(_15509_));
 sg13g2_nor2_1 _29151_ (.A(_03053_),
    .B(net6722),
    .Y(_15510_));
 sg13g2_a21oi_1 _29152_ (.A1(net7272),
    .A2(net6724),
    .Y(_15511_),
    .B1(_15510_));
 sg13g2_a21oi_1 _29153_ (.A1(net6735),
    .A2(_15511_),
    .Y(net490),
    .B1(_15509_));
 sg13g2_and2_1 _29154_ (.A(net6732),
    .B(_15437_),
    .X(_15512_));
 sg13g2_a21oi_1 _29155_ (.A1(net6744),
    .A2(_15494_),
    .Y(net491),
    .B1(_15512_));
 sg13g2_and2_1 _29156_ (.A(net6745),
    .B(_15497_),
    .X(_15513_));
 sg13g2_a21oi_1 _29157_ (.A1(net6733),
    .A2(_15442_),
    .Y(net492),
    .B1(_15513_));
 sg13g2_mux4_1 _29158_ (.S0(net6746),
    .A0(_03256_),
    .A1(_02713_),
    .A2(_02171_),
    .A3(_10750_),
    .S1(net6727),
    .X(net493));
 sg13g2_a21o_1 _29159_ (.A2(net7039),
    .A1(net7682),
    .B1(_15466_),
    .X(_15514_));
 sg13g2_mux2_1 _29160_ (.A0(_15448_),
    .A1(_15499_),
    .S(net6744),
    .X(net494));
 sg13g2_and2_1 _29161_ (.A(net6742),
    .B(_15503_),
    .X(_15515_));
 sg13g2_a21oi_1 _29162_ (.A1(net6734),
    .A2(_15451_),
    .Y(net495),
    .B1(_15515_));
 sg13g2_a21oi_1 _29163_ (.A1(net7682),
    .A2(net7039),
    .Y(_15516_),
    .B1(_15466_));
 sg13g2_and2_1 _29164_ (.A(net6742),
    .B(_15504_),
    .X(_15517_));
 sg13g2_a21oi_1 _29165_ (.A1(net6734),
    .A2(_15457_),
    .Y(net496),
    .B1(_15517_));
 sg13g2_and2_1 _29166_ (.A(net6733),
    .B(_15464_),
    .X(_15518_));
 sg13g2_a21oi_1 _29167_ (.A1(net6745),
    .A2(_15508_),
    .Y(net498),
    .B1(_15518_));
 sg13g2_and2_1 _29168_ (.A(net6734),
    .B(_15469_),
    .X(_15519_));
 sg13g2_a21oi_1 _29169_ (.A1(net6743),
    .A2(_15511_),
    .Y(net499),
    .B1(_15519_));
 sg13g2_nand2_1 _29170_ (.Y(_15520_),
    .A(net7883),
    .B(_01598_));
 sg13g2_nand2b_1 _29171_ (.Y(_15521_),
    .B(_01563_),
    .A_N(net7883));
 sg13g2_nand3_1 _29172_ (.B(_15520_),
    .C(_15521_),
    .A(net7450),
    .Y(_15522_));
 sg13g2_inv_1 _29173_ (.Y(_15523_),
    .A(_01702_));
 sg13g2_nand2_1 _29174_ (.Y(_15524_),
    .A(net7848),
    .B(_01528_));
 sg13g2_nand2b_1 _29175_ (.Y(_15525_),
    .B(_01493_),
    .A_N(net7848));
 sg13g2_nand4_1 _29176_ (.B(net7494),
    .C(_15524_),
    .A(net7512),
    .Y(_15526_),
    .D(_15525_));
 sg13g2_nand2_1 _29177_ (.Y(_15527_),
    .A(net7850),
    .B(_00827_));
 sg13g2_nand2b_1 _29178_ (.Y(_15528_),
    .B(_00795_),
    .A_N(net7849));
 sg13g2_inv_1 _29179_ (.Y(_15529_),
    .A(_01701_));
 sg13g2_nand4_1 _29180_ (.B(net7471),
    .C(_15527_),
    .A(net7548),
    .Y(_15530_),
    .D(_15528_));
 sg13g2_nand2_1 _29181_ (.Y(_15531_),
    .A(net7848),
    .B(_00894_));
 sg13g2_nand2b_1 _29182_ (.Y(_15532_),
    .B(_00859_),
    .A_N(net7848));
 sg13g2_nand4_1 _29183_ (.B(net7462),
    .C(_15531_),
    .A(net7548),
    .Y(_15533_),
    .D(_15532_));
 sg13g2_nand2_1 _29184_ (.Y(_15534_),
    .A(net7847),
    .B(_01035_));
 sg13g2_nand2b_1 _29185_ (.Y(_15535_),
    .B(_01000_),
    .A_N(net7847));
 sg13g2_inv_1 _29186_ (.Y(_15536_),
    .A(_01699_));
 sg13g2_nand4_1 _29187_ (.B(net7525),
    .C(_15534_),
    .A(net7548),
    .Y(_15537_),
    .D(_15535_));
 sg13g2_nand2_1 _29188_ (.Y(_15538_),
    .A(net7847),
    .B(_00965_));
 sg13g2_nand2b_1 _29189_ (.Y(_15539_),
    .B(_00930_),
    .A_N(net7847));
 sg13g2_nand4_1 _29190_ (.B(net7512),
    .C(_15538_),
    .A(net7548),
    .Y(_15540_),
    .D(_15539_));
 sg13g2_nand2_1 _29191_ (.Y(_15541_),
    .A(net7848),
    .B(_01387_));
 sg13g2_inv_1 _29192_ (.Y(_15542_),
    .A(_01698_));
 sg13g2_nand2b_1 _29193_ (.Y(_15543_),
    .B(_01352_),
    .A_N(net7848));
 sg13g2_nand4_1 _29194_ (.B(net7471),
    .C(_15541_),
    .A(net7494),
    .Y(_15544_),
    .D(_15543_));
 sg13g2_nand2_1 _29195_ (.Y(_15545_),
    .A(net7848),
    .B(_01458_));
 sg13g2_nand2b_1 _29196_ (.Y(_15546_),
    .B(_01422_),
    .A_N(net7848));
 sg13g2_nand4_1 _29197_ (.B(net7462),
    .C(_15545_),
    .A(net7494),
    .Y(_15547_),
    .D(_15546_));
 sg13g2_nand4_1 _29198_ (.B(_15537_),
    .C(_15544_),
    .A(_15530_),
    .Y(_15548_),
    .D(_15547_));
 sg13g2_nand4_1 _29199_ (.B(_15526_),
    .C(_15533_),
    .A(_15522_),
    .Y(_15549_),
    .D(_15540_));
 sg13g2_mux2_1 _29200_ (.A0(_01291_),
    .A1(_00635_),
    .S(net7851),
    .X(_15550_));
 sg13g2_and2_1 _29201_ (.A(net7851),
    .B(_00939_),
    .X(_15551_));
 sg13g2_mux2_1 _29202_ (.A0(_00667_),
    .A1(_00699_),
    .S(net7851),
    .X(_15552_));
 sg13g2_mux2_1 _29203_ (.A0(_00731_),
    .A1(_00763_),
    .S(net7851),
    .X(_15553_));
 sg13g2_mux4_1 _29204_ (.S0(net7811),
    .A0(_15551_),
    .A1(_15552_),
    .A2(_15550_),
    .A3(_15553_),
    .S1(net7826),
    .X(_15554_));
 sg13g2_nor2_1 _29205_ (.A(net7529),
    .B(_15554_),
    .Y(_15555_));
 sg13g2_inv_1 _29206_ (.Y(_15556_),
    .A(_01692_));
 sg13g2_mux4_1 _29207_ (.S0(net7892),
    .A0(_01070_),
    .A1(_01106_),
    .A2(_01141_),
    .A3(_01176_),
    .S1(net7825),
    .X(_15557_));
 sg13g2_mux4_1 _29208_ (.S0(net7892),
    .A0(_01211_),
    .A1(_01246_),
    .A2(_01282_),
    .A3(_01317_),
    .S1(net7825),
    .X(_15558_));
 sg13g2_or2_1 _29209_ (.X(_15559_),
    .B(_15558_),
    .A(net7443));
 sg13g2_inv_1 _29210_ (.Y(_15560_),
    .A(_01689_));
 sg13g2_o21ai_1 _29211_ (.B1(_15559_),
    .Y(_15561_),
    .A1(net7421),
    .A2(_15557_));
 sg13g2_nor4_1 _29212_ (.A(_15548_),
    .B(_15549_),
    .C(_15555_),
    .D(_15561_),
    .Y(_15562_));
 sg13g2_or4_1 _29213_ (.A(_15548_),
    .B(_15549_),
    .C(_15555_),
    .D(_15561_),
    .X(_15563_));
 sg13g2_nand2b_1 _29214_ (.Y(_15564_),
    .B(net7998),
    .A_N(_01640_));
 sg13g2_o21ai_1 _29215_ (.B1(_15564_),
    .Y(_15565_),
    .A1(_01670_),
    .A2(_09260_));
 sg13g2_a221oi_1 _29216_ (.B2(_00541_),
    .C1(_15565_),
    .B1(_15563_),
    .A1(_09275_),
    .Y(_15566_),
    .A2(_15462_));
 sg13g2_nor2_1 _29217_ (.A(net7366),
    .B(_15566_),
    .Y(_15567_));
 sg13g2_a21oi_1 _29218_ (.A1(net6917),
    .A2(_15514_),
    .Y(_15568_),
    .B1(_15567_));
 sg13g2_o21ai_1 _29219_ (.B1(_15568_),
    .Y(_15569_),
    .A1(_08228_),
    .A2(_15514_));
 sg13g2_mux4_1 _29220_ (.S0(net7777),
    .A0(_00796_),
    .A1(_00828_),
    .A2(_00860_),
    .A3(_00896_),
    .S1(net7726),
    .X(_15570_));
 sg13g2_and2_1 _29221_ (.A(net7605),
    .B(_15570_),
    .X(_15571_));
 sg13g2_nand2_1 _29222_ (.Y(_15572_),
    .A(net7714),
    .B(_00764_));
 sg13g2_nand2b_1 _29223_ (.Y(_15573_),
    .B(_00636_),
    .A_N(net7714));
 sg13g2_a21oi_1 _29224_ (.A1(_15572_),
    .A2(_15573_),
    .Y(_15574_),
    .B1(net7600));
 sg13g2_nand3b_1 _29225_ (.B(net7774),
    .C(_00950_),
    .Y(_15575_),
    .A_N(net7744));
 sg13g2_nand3b_1 _29226_ (.B(_01302_),
    .C(net7744),
    .Y(_15576_),
    .A_N(net7775));
 sg13g2_a21oi_1 _29227_ (.A1(_15575_),
    .A2(_15576_),
    .Y(_15577_),
    .B1(_08306_));
 sg13g2_nor4_1 _29228_ (.A(net7686),
    .B(_15571_),
    .C(_15574_),
    .D(_15577_),
    .Y(_15578_));
 sg13g2_mux4_1 _29229_ (.S0(net7777),
    .A0(_00931_),
    .A1(_00966_),
    .A2(_01001_),
    .A3(_01036_),
    .S1(net7728),
    .X(_15579_));
 sg13g2_mux2_1 _29230_ (.A0(_00668_),
    .A1(_00700_),
    .S(net7775),
    .X(_15580_));
 sg13g2_a221oi_1 _29231_ (.B2(net7518),
    .C1(net7695),
    .B1(_15580_),
    .A1(_00732_),
    .Y(_15581_),
    .A2(net7594));
 sg13g2_o21ai_1 _29232_ (.B1(net7714),
    .Y(_15582_),
    .A1(net7533),
    .A2(_15579_));
 \ALU_33_0_33_0_33_unused_CO_X_Y[0]_KOGGE_STONE  \alu_adder_result_ex\\ALU_33_0_33_0_33_unused_CO_X_Y[0]_HAN_CARLSON  (.A({_03632_,
    _03581_,
    _03511_,
    _03442_,
    _03373_,
    _03301_,
    _03230_,
    _03165_,
    _03091_,
    _03024_,
    _02957_,
    _02890_,
    _02824_,
    _02752_,
    _02687_,
    _02622_,
    _02555_,
    _02509_,
    _02445_,
    _02368_,
    _02289_,
    _02213_,
    _02146_,
    _02071_,
    _15569_,
    _15132_,
    _14300_,
    _13402_,
    _12286_,
    _11205_,
    _10414_,
    _09346_,
    _08254_}),
    .B({_03814_,
    _03808_,
    _03803_,
    _03798_,
    _03792_,
    _03787_,
    _03782_,
    _03777_,
    _03772_,
    _03767_,
    _03762_,
    _03757_,
    _03752_,
    _03747_,
    _03742_,
    _03737_,
    _03732_,
    _03727_,
    _03722_,
    _03717_,
    _03712_,
    _03707_,
    _03702_,
    _03697_,
    _03692_,
    _03687_,
    _03682_,
    _03677_,
    _03671_,
    _03665_,
    _03659_,
    _03652_,
    net_8}),
    .BI(net_6),
    .CI(net_7),
    .Y\[32:1\]({net462,
    net461,
    net459,
    net458,
    net457,
    net456,
    net455,
    net454,
    net453,
    net452,
    net451,
    net450,
    net449,
    net448,
    net447,
    net446,
    net445,
    net444,
    net443,
    net442,
    net441,
    net440,
    net469,
    net468,
    net467,
    net466,
    net465,
    net464,
    net463,
    net460,
    \alu_adder_result_ex[1] ,
    \alu_adder_result_ex[0] }));
 sg13g2_tielo \alu_adder_result_ex\\ALU_33_0_33_0_33_unused_CO_X_Y[0]_HAN_CARLSON_13  (.L_LO(net_6));
 sg13g2_tielo \alu_adder_result_ex\\ALU_33_0_33_0_33_unused_CO_X_Y[0]_HAN_CARLSON_14  (.L_LO(net_7));
 sg13g2_tiehi \alu_adder_result_ex\\ALU_33_0_33_0_33_unused_CO_X_Y[0]_HAN_CARLSON_15  (.L_HI(net_8));
 sg13g2_buf_16 clkbuf_0__06563_ (.X(clknet_0__06563_),
    .A(_06563_));
 sg13g2_buf_16 clkbuf_0_clk_i (.X(clknet_0_clk_i),
    .A(clk_i));
 sg13g2_buf_16 clkbuf_0_clk_i_regs (.X(clknet_0_clk_i_regs),
    .A(clk_i_regs));
 sg13g2_buf_16 clkbuf_1_0_0__06563_ (.X(clknet_1_0_0__06563_),
    .A(clknet_0__06563_));
 sg13g2_buf_16 clkbuf_1_0_0_clk_i_regs (.X(clknet_1_0_0_clk_i_regs),
    .A(clknet_0_clk_i_regs));
 sg13g2_buf_16 clkbuf_1_0__f_clk_i (.X(clknet_1_0__leaf_clk_i),
    .A(clknet_0_clk_i));
 sg13g2_buf_16 clkbuf_1_1_0__06563_ (.X(clknet_1_1_0__06563_),
    .A(clknet_0__06563_));
 sg13g2_buf_16 clkbuf_1_1_0_clk_i_regs (.X(clknet_1_1_0_clk_i_regs),
    .A(clknet_0_clk_i_regs));
 sg13g2_buf_16 clkbuf_2_0_0__06563_ (.X(clknet_2_0_0__06563_),
    .A(clknet_1_0_0__06563_));
 sg13g2_buf_16 clkbuf_2_0_0_clk_i_regs (.X(clknet_2_0_0_clk_i_regs),
    .A(clknet_1_0_0_clk_i_regs));
 sg13g2_buf_16 clkbuf_2_1_0__06563_ (.X(clknet_2_1_0__06563_),
    .A(clknet_1_0_0__06563_));
 sg13g2_buf_16 clkbuf_2_1_0_clk_i_regs (.X(clknet_2_1_0_clk_i_regs),
    .A(clknet_1_0_0_clk_i_regs));
 sg13g2_buf_16 clkbuf_2_2_0__06563_ (.X(clknet_2_2_0__06563_),
    .A(clknet_1_1_0__06563_));
 sg13g2_buf_16 clkbuf_2_2_0_clk_i_regs (.X(clknet_2_2_0_clk_i_regs),
    .A(clknet_1_1_0_clk_i_regs));
 sg13g2_buf_16 clkbuf_2_3_0__06563_ (.X(clknet_2_3_0__06563_),
    .A(clknet_1_1_0__06563_));
 sg13g2_buf_16 clkbuf_2_3_0_clk_i_regs (.X(clknet_2_3_0_clk_i_regs),
    .A(clknet_1_1_0_clk_i_regs));
 sg13g2_buf_16 clkbuf_3_0_0__06563_ (.X(clknet_3_0_0__06563_),
    .A(clknet_2_0_0__06563_));
 sg13g2_buf_16 clkbuf_3_0_0_clk_i_regs (.X(clknet_3_0_0_clk_i_regs),
    .A(clknet_2_0_0_clk_i_regs));
 sg13g2_buf_16 clkbuf_3_1_0__06563_ (.X(clknet_3_1_0__06563_),
    .A(clknet_2_0_0__06563_));
 sg13g2_buf_16 clkbuf_3_1_0_clk_i_regs (.X(clknet_3_1_0_clk_i_regs),
    .A(clknet_2_0_0_clk_i_regs));
 sg13g2_buf_16 clkbuf_3_2_0__06563_ (.X(clknet_3_2_0__06563_),
    .A(clknet_2_1_0__06563_));
 sg13g2_buf_16 clkbuf_3_2_0_clk_i_regs (.X(clknet_3_2_0_clk_i_regs),
    .A(clknet_2_1_0_clk_i_regs));
 sg13g2_buf_16 clkbuf_3_3_0__06563_ (.X(clknet_3_3_0__06563_),
    .A(clknet_2_1_0__06563_));
 sg13g2_buf_16 clkbuf_3_3_0_clk_i_regs (.X(clknet_3_3_0_clk_i_regs),
    .A(clknet_2_1_0_clk_i_regs));
 sg13g2_buf_16 clkbuf_3_4_0__06563_ (.X(clknet_3_4_0__06563_),
    .A(clknet_2_2_0__06563_));
 sg13g2_buf_16 clkbuf_3_4_0_clk_i_regs (.X(clknet_3_4_0_clk_i_regs),
    .A(clknet_2_2_0_clk_i_regs));
 sg13g2_buf_16 clkbuf_3_5_0__06563_ (.X(clknet_3_5_0__06563_),
    .A(clknet_2_2_0__06563_));
 sg13g2_buf_16 clkbuf_3_5_0_clk_i_regs (.X(clknet_3_5_0_clk_i_regs),
    .A(clknet_2_2_0_clk_i_regs));
 sg13g2_buf_16 clkbuf_3_6_0__06563_ (.X(clknet_3_6_0__06563_),
    .A(clknet_2_3_0__06563_));
 sg13g2_buf_16 clkbuf_3_6_0_clk_i_regs (.X(clknet_3_6_0_clk_i_regs),
    .A(clknet_2_3_0_clk_i_regs));
 sg13g2_buf_16 clkbuf_3_7_0__06563_ (.X(clknet_3_7_0__06563_),
    .A(clknet_2_3_0__06563_));
 sg13g2_buf_16 clkbuf_3_7_0_clk_i_regs (.X(clknet_3_7_0_clk_i_regs),
    .A(clknet_2_3_0_clk_i_regs));
 sg13g2_buf_16 clkbuf_leaf_0__06563_ (.X(clknet_leaf_0__06563_),
    .A(clknet_3_0_0__06563_));
 sg13g2_buf_16 clkbuf_leaf_0_clk_i_regs (.X(clknet_leaf_0_clk_i_regs),
    .A(clknet_3_0_0_clk_i_regs));
 sg13g2_buf_16 clkbuf_leaf_10__06563_ (.X(clknet_leaf_10__06563_),
    .A(clknet_3_6_0__06563_));
 sg13g2_buf_16 clkbuf_leaf_10_clk_i_regs (.X(clknet_leaf_10_clk_i_regs),
    .A(clknet_3_1_0_clk_i_regs));
 sg13g2_buf_16 clkbuf_leaf_11__06563_ (.X(clknet_leaf_11__06563_),
    .A(clknet_3_6_0__06563_));
 sg13g2_buf_16 clkbuf_leaf_11_clk_i_regs (.X(clknet_leaf_11_clk_i_regs),
    .A(clknet_3_4_0_clk_i_regs));
 sg13g2_buf_16 clkbuf_leaf_12__06563_ (.X(clknet_leaf_12__06563_),
    .A(clknet_3_7_0__06563_));
 sg13g2_buf_16 clkbuf_leaf_12_clk_i_regs (.X(clknet_leaf_12_clk_i_regs),
    .A(clknet_3_4_0_clk_i_regs));
 sg13g2_buf_16 clkbuf_leaf_13__06563_ (.X(clknet_leaf_13__06563_),
    .A(clknet_3_7_0__06563_));
 sg13g2_buf_16 clkbuf_leaf_13_clk_i_regs (.X(clknet_leaf_13_clk_i_regs),
    .A(clknet_3_4_0_clk_i_regs));
 sg13g2_buf_16 clkbuf_leaf_14__06563_ (.X(clknet_leaf_14__06563_),
    .A(clknet_3_7_0__06563_));
 sg13g2_buf_16 clkbuf_leaf_14_clk_i_regs (.X(clknet_leaf_14_clk_i_regs),
    .A(clknet_3_4_0_clk_i_regs));
 sg13g2_buf_16 clkbuf_leaf_15__06563_ (.X(clknet_leaf_15__06563_),
    .A(clknet_3_7_0__06563_));
 sg13g2_buf_16 clkbuf_leaf_15_clk_i_regs (.X(clknet_leaf_15_clk_i_regs),
    .A(clknet_3_5_0_clk_i_regs));
 sg13g2_buf_16 clkbuf_leaf_16__06563_ (.X(clknet_leaf_16__06563_),
    .A(clknet_3_7_0__06563_));
 sg13g2_buf_16 clkbuf_leaf_16_clk_i_regs (.X(clknet_leaf_16_clk_i_regs),
    .A(clknet_3_5_0_clk_i_regs));
 sg13g2_buf_16 clkbuf_leaf_17__06563_ (.X(clknet_leaf_17__06563_),
    .A(clknet_3_5_0__06563_));
 sg13g2_buf_16 clkbuf_leaf_17_clk_i_regs (.X(clknet_leaf_17_clk_i_regs),
    .A(clknet_3_5_0_clk_i_regs));
 sg13g2_buf_16 clkbuf_leaf_18__06563_ (.X(clknet_leaf_18__06563_),
    .A(clknet_3_7_0__06563_));
 sg13g2_buf_16 clkbuf_leaf_18_clk_i_regs (.X(clknet_leaf_18_clk_i_regs),
    .A(clknet_3_5_0_clk_i_regs));
 sg13g2_buf_16 clkbuf_leaf_19__06563_ (.X(clknet_leaf_19__06563_),
    .A(clknet_3_6_0__06563_));
 sg13g2_buf_16 clkbuf_leaf_19_clk_i_regs (.X(clknet_leaf_19_clk_i_regs),
    .A(clknet_3_5_0_clk_i_regs));
 sg13g2_buf_16 clkbuf_leaf_1__06563_ (.X(clknet_leaf_1__06563_),
    .A(clknet_3_2_0__06563_));
 sg13g2_buf_16 clkbuf_leaf_1_clk_i_regs (.X(clknet_leaf_1_clk_i_regs),
    .A(clknet_3_0_0_clk_i_regs));
 sg13g2_buf_16 clkbuf_leaf_20__06563_ (.X(clknet_leaf_20__06563_),
    .A(clknet_3_3_0__06563_));
 sg13g2_buf_16 clkbuf_leaf_20_clk_i_regs (.X(clknet_leaf_20_clk_i_regs),
    .A(clknet_3_4_0_clk_i_regs));
 sg13g2_buf_16 clkbuf_leaf_21__06563_ (.X(clknet_leaf_21__06563_),
    .A(clknet_3_3_0__06563_));
 sg13g2_buf_16 clkbuf_leaf_21_clk_i_regs (.X(clknet_leaf_21_clk_i_regs),
    .A(clknet_3_3_0_clk_i_regs));
 sg13g2_buf_16 clkbuf_leaf_22__06563_ (.X(clknet_leaf_22__06563_),
    .A(clknet_3_5_0__06563_));
 sg13g2_buf_16 clkbuf_leaf_22_clk_i_regs (.X(clknet_leaf_22_clk_i_regs),
    .A(clknet_3_6_0_clk_i_regs));
 sg13g2_buf_16 clkbuf_leaf_23__06563_ (.X(clknet_leaf_23__06563_),
    .A(clknet_3_5_0__06563_));
 sg13g2_buf_16 clkbuf_leaf_23_clk_i_regs (.X(clknet_leaf_23_clk_i_regs),
    .A(clknet_3_5_0_clk_i_regs));
 sg13g2_buf_16 clkbuf_leaf_24__06563_ (.X(clknet_leaf_24__06563_),
    .A(clknet_3_5_0__06563_));
 sg13g2_buf_16 clkbuf_leaf_24_clk_i_regs (.X(clknet_leaf_24_clk_i_regs),
    .A(clknet_3_7_0_clk_i_regs));
 sg13g2_buf_16 clkbuf_leaf_25__06563_ (.X(clknet_leaf_25__06563_),
    .A(clknet_3_5_0__06563_));
 sg13g2_buf_16 clkbuf_leaf_25_clk_i_regs (.X(clknet_leaf_25_clk_i_regs),
    .A(clknet_3_7_0_clk_i_regs));
 sg13g2_buf_16 clkbuf_leaf_26__06563_ (.X(clknet_leaf_26__06563_),
    .A(clknet_3_4_0__06563_));
 sg13g2_buf_16 clkbuf_leaf_26_clk_i_regs (.X(clknet_leaf_26_clk_i_regs),
    .A(clknet_3_7_0_clk_i_regs));
 sg13g2_buf_16 clkbuf_leaf_27__06563_ (.X(clknet_leaf_27__06563_),
    .A(clknet_3_4_0__06563_));
 sg13g2_buf_16 clkbuf_leaf_27_clk_i_regs (.X(clknet_leaf_27_clk_i_regs),
    .A(clknet_3_7_0_clk_i_regs));
 sg13g2_buf_16 clkbuf_leaf_28__06563_ (.X(clknet_leaf_28__06563_),
    .A(clknet_3_4_0__06563_));
 sg13g2_buf_16 clkbuf_leaf_28_clk_i_regs (.X(clknet_leaf_28_clk_i_regs),
    .A(clknet_3_7_0_clk_i_regs));
 sg13g2_buf_16 clkbuf_leaf_29__06563_ (.X(clknet_leaf_29__06563_),
    .A(clknet_3_5_0__06563_));
 sg13g2_buf_16 clkbuf_leaf_29_clk_i_regs (.X(clknet_leaf_29_clk_i_regs),
    .A(clknet_3_7_0_clk_i_regs));
 sg13g2_buf_16 clkbuf_leaf_2__06563_ (.X(clknet_leaf_2__06563_),
    .A(clknet_3_2_0__06563_));
 sg13g2_buf_16 clkbuf_leaf_2_clk_i_regs (.X(clknet_leaf_2_clk_i_regs),
    .A(clknet_3_1_0_clk_i_regs));
 sg13g2_buf_16 clkbuf_leaf_30__06563_ (.X(clknet_leaf_30__06563_),
    .A(clknet_3_4_0__06563_));
 sg13g2_buf_16 clkbuf_leaf_30_clk_i_regs (.X(clknet_leaf_30_clk_i_regs),
    .A(clknet_3_6_0_clk_i_regs));
 sg13g2_buf_16 clkbuf_leaf_31__06563_ (.X(clknet_leaf_31__06563_),
    .A(clknet_3_4_0__06563_));
 sg13g2_buf_16 clkbuf_leaf_31_clk_i_regs (.X(clknet_leaf_31_clk_i_regs),
    .A(clknet_3_6_0_clk_i_regs));
 sg13g2_buf_16 clkbuf_leaf_32__06563_ (.X(clknet_leaf_32__06563_),
    .A(clknet_3_4_0__06563_));
 sg13g2_buf_16 clkbuf_leaf_32_clk_i_regs (.X(clknet_leaf_32_clk_i_regs),
    .A(clknet_3_6_0_clk_i_regs));
 sg13g2_buf_16 clkbuf_leaf_33__06563_ (.X(clknet_leaf_33__06563_),
    .A(clknet_3_4_0__06563_));
 sg13g2_buf_16 clkbuf_leaf_33_clk_i_regs (.X(clknet_leaf_33_clk_i_regs),
    .A(clknet_3_6_0_clk_i_regs));
 sg13g2_buf_16 clkbuf_leaf_34__06563_ (.X(clknet_leaf_34__06563_),
    .A(clknet_3_1_0__06563_));
 sg13g2_buf_16 clkbuf_leaf_34_clk_i_regs (.X(clknet_leaf_34_clk_i_regs),
    .A(clknet_3_6_0_clk_i_regs));
 sg13g2_buf_16 clkbuf_leaf_35__06563_ (.X(clknet_leaf_35__06563_),
    .A(clknet_3_1_0__06563_));
 sg13g2_buf_16 clkbuf_leaf_35_clk_i_regs (.X(clknet_leaf_35_clk_i_regs),
    .A(clknet_3_3_0_clk_i_regs));
 sg13g2_buf_16 clkbuf_leaf_36__06563_ (.X(clknet_leaf_36__06563_),
    .A(clknet_3_1_0__06563_));
 sg13g2_buf_16 clkbuf_leaf_36_clk_i_regs (.X(clknet_leaf_36_clk_i_regs),
    .A(clknet_3_2_0_clk_i_regs));
 sg13g2_buf_16 clkbuf_leaf_37__06563_ (.X(clknet_leaf_37__06563_),
    .A(clknet_3_1_0__06563_));
 sg13g2_buf_16 clkbuf_leaf_37_clk_i_regs (.X(clknet_leaf_37_clk_i_regs),
    .A(clknet_3_2_0_clk_i_regs));
 sg13g2_buf_16 clkbuf_leaf_38__06563_ (.X(clknet_leaf_38__06563_),
    .A(clknet_3_1_0__06563_));
 sg13g2_buf_16 clkbuf_leaf_38_clk_i_regs (.X(clknet_leaf_38_clk_i_regs),
    .A(clknet_3_2_0_clk_i_regs));
 sg13g2_buf_16 clkbuf_leaf_39__06563_ (.X(clknet_leaf_39__06563_),
    .A(clknet_3_1_0__06563_));
 sg13g2_buf_16 clkbuf_leaf_39_clk_i_regs (.X(clknet_leaf_39_clk_i_regs),
    .A(clknet_3_2_0_clk_i_regs));
 sg13g2_buf_16 clkbuf_leaf_3__06563_ (.X(clknet_leaf_3__06563_),
    .A(clknet_3_2_0__06563_));
 sg13g2_buf_16 clkbuf_leaf_3_clk_i_regs (.X(clknet_leaf_3_clk_i_regs),
    .A(clknet_3_1_0_clk_i_regs));
 sg13g2_buf_16 clkbuf_leaf_40__06563_ (.X(clknet_leaf_40__06563_),
    .A(clknet_3_3_0__06563_));
 sg13g2_buf_16 clkbuf_leaf_40_clk_i_regs (.X(clknet_leaf_40_clk_i_regs),
    .A(clknet_3_2_0_clk_i_regs));
 sg13g2_buf_16 clkbuf_leaf_41__06563_ (.X(clknet_leaf_41__06563_),
    .A(clknet_3_3_0__06563_));
 sg13g2_buf_16 clkbuf_leaf_41_clk_i_regs (.X(clknet_leaf_41_clk_i_regs),
    .A(clknet_3_2_0_clk_i_regs));
 sg13g2_buf_16 clkbuf_leaf_42__06563_ (.X(clknet_leaf_42__06563_),
    .A(clknet_3_2_0__06563_));
 sg13g2_buf_16 clkbuf_leaf_42_clk_i_regs (.X(clknet_leaf_42_clk_i_regs),
    .A(clknet_3_3_0_clk_i_regs));
 sg13g2_buf_16 clkbuf_leaf_43__06563_ (.X(clknet_leaf_43__06563_),
    .A(clknet_3_2_0__06563_));
 sg13g2_buf_16 clkbuf_leaf_43_clk_i_regs (.X(clknet_leaf_43_clk_i_regs),
    .A(clknet_3_1_0_clk_i_regs));
 sg13g2_buf_16 clkbuf_leaf_44__06563_ (.X(clknet_leaf_44__06563_),
    .A(clknet_3_2_0__06563_));
 sg13g2_buf_16 clkbuf_leaf_44_clk_i_regs (.X(clknet_leaf_44_clk_i_regs),
    .A(clknet_3_0_0_clk_i_regs));
 sg13g2_buf_16 clkbuf_leaf_45__06563_ (.X(clknet_leaf_45__06563_),
    .A(clknet_3_3_0__06563_));
 sg13g2_buf_16 clkbuf_leaf_45_clk_i_regs (.X(clknet_leaf_45_clk_i_regs),
    .A(clknet_3_0_0_clk_i_regs));
 sg13g2_buf_16 clkbuf_leaf_46__06563_ (.X(clknet_leaf_46__06563_),
    .A(clknet_3_0_0__06563_));
 sg13g2_buf_16 clkbuf_leaf_46_clk_i_regs (.X(clknet_leaf_46_clk_i_regs),
    .A(clknet_3_0_0_clk_i_regs));
 sg13g2_buf_16 clkbuf_leaf_47__06563_ (.X(clknet_leaf_47__06563_),
    .A(clknet_3_0_0__06563_));
 sg13g2_buf_16 clkbuf_leaf_47_clk_i_regs (.X(clknet_leaf_47_clk_i_regs),
    .A(clknet_3_0_0_clk_i_regs));
 sg13g2_buf_16 clkbuf_leaf_48__06563_ (.X(clknet_leaf_48__06563_),
    .A(clknet_3_0_0__06563_));
 sg13g2_buf_16 clkbuf_leaf_48_clk_i_regs (.X(clknet_leaf_48_clk_i_regs),
    .A(clknet_3_0_0_clk_i_regs));
 sg13g2_buf_16 clkbuf_leaf_49__06563_ (.X(clknet_leaf_49__06563_),
    .A(clknet_3_0_0__06563_));
 sg13g2_buf_16 clkbuf_leaf_4__06563_ (.X(clknet_leaf_4__06563_),
    .A(clknet_3_2_0__06563_));
 sg13g2_buf_16 clkbuf_leaf_4_clk_i_regs (.X(clknet_leaf_4_clk_i_regs),
    .A(clknet_3_3_0_clk_i_regs));
 sg13g2_buf_16 clkbuf_leaf_50__06563_ (.X(clknet_leaf_50__06563_),
    .A(clknet_3_0_0__06563_));
 sg13g2_buf_16 clkbuf_leaf_51__06563_ (.X(clknet_leaf_51__06563_),
    .A(clknet_3_0_0__06563_));
 sg13g2_buf_16 clkbuf_leaf_5__06563_ (.X(clknet_leaf_5__06563_),
    .A(clknet_3_3_0__06563_));
 sg13g2_buf_16 clkbuf_leaf_5_clk_i_regs (.X(clknet_leaf_5_clk_i_regs),
    .A(clknet_3_1_0_clk_i_regs));
 sg13g2_buf_16 clkbuf_leaf_6__06563_ (.X(clknet_leaf_6__06563_),
    .A(clknet_3_6_0__06563_));
 sg13g2_buf_16 clkbuf_leaf_6_clk_i_regs (.X(clknet_leaf_6_clk_i_regs),
    .A(clknet_3_3_0_clk_i_regs));
 sg13g2_buf_16 clkbuf_leaf_7__06563_ (.X(clknet_leaf_7__06563_),
    .A(clknet_3_6_0__06563_));
 sg13g2_buf_16 clkbuf_leaf_7_clk_i_regs (.X(clknet_leaf_7_clk_i_regs),
    .A(clknet_3_3_0_clk_i_regs));
 sg13g2_buf_16 clkbuf_leaf_8__06563_ (.X(clknet_leaf_8__06563_),
    .A(clknet_3_6_0__06563_));
 sg13g2_buf_16 clkbuf_leaf_8_clk_i_regs (.X(clknet_leaf_8_clk_i_regs),
    .A(clknet_3_1_0_clk_i_regs));
 sg13g2_buf_16 clkbuf_leaf_9__06563_ (.X(clknet_leaf_9__06563_),
    .A(clknet_3_6_0__06563_));
 sg13g2_buf_16 clkbuf_leaf_9_clk_i_regs (.X(clknet_leaf_9_clk_i_regs),
    .A(clknet_3_4_0_clk_i_regs));
 sg13g2_buf_16 clkbuf_regs_0_core_clock (.X(clk_i_regs),
    .A(delaynet_2_core_clock));
 sg13g2_buf_16 clkload0 (.A(clknet_3_1_0_clk_i_regs));
 sg13g2_inv_4 clkload1 (.A(clknet_leaf_1_clk_i_regs));
 sg13g2_buf_8 clkload10 (.A(clknet_leaf_8_clk_i_regs));
 sg13g2_buf_8 clkload11 (.A(clknet_leaf_10_clk_i_regs));
 sg13g2_inv_8 clkload12 (.A(clknet_leaf_38_clk_i_regs));
 sg13g2_inv_1 clkload13 (.A(clknet_leaf_40_clk_i_regs));
 sg13g2_buf_8 clkload14 (.A(clknet_leaf_41_clk_i_regs));
 sg13g2_inv_1 clkload15 (.A(clknet_leaf_4_clk_i_regs));
 sg13g2_inv_1 clkload16 (.A(clknet_leaf_6_clk_i_regs));
 sg13g2_inv_2 clkload17 (.A(clknet_leaf_7_clk_i_regs));
 sg13g2_buf_8 clkload18 (.A(clknet_leaf_21_clk_i_regs));
 sg13g2_buf_8 clkload19 (.A(clknet_leaf_42_clk_i_regs));
 sg13g2_inv_2 clkload2 (.A(clknet_leaf_44_clk_i_regs));
 sg13g2_buf_16 clkload20 (.A(clknet_leaf_9_clk_i_regs));
 sg13g2_buf_16 clkload21 (.A(clknet_leaf_12_clk_i_regs));
 sg13g2_inv_4 clkload22 (.A(clknet_leaf_13_clk_i_regs));
 sg13g2_buf_16 clkload23 (.A(clknet_leaf_20_clk_i_regs));
 sg13g2_buf_8 clkload24 (.A(clknet_leaf_15_clk_i_regs));
 sg13g2_buf_16 clkload25 (.A(clknet_leaf_17_clk_i_regs));
 sg13g2_inv_4 clkload26 (.A(clknet_leaf_18_clk_i_regs));
 sg13g2_inv_4 clkload27 (.A(clknet_leaf_19_clk_i_regs));
 sg13g2_buf_16 clkload28 (.A(clknet_leaf_23_clk_i_regs));
 sg13g2_buf_8 clkload29 (.A(clknet_leaf_22_clk_i_regs));
 sg13g2_inv_2 clkload3 (.A(clknet_leaf_45_clk_i_regs));
 sg13g2_inv_4 clkload30 (.A(clknet_leaf_30_clk_i_regs));
 sg13g2_inv_2 clkload31 (.A(clknet_leaf_24_clk_i_regs));
 sg13g2_buf_8 clkload32 (.A(clknet_leaf_26_clk_i_regs));
 sg13g2_buf_8 clkload33 (.A(clknet_leaf_27_clk_i_regs));
 sg13g2_inv_2 clkload34 (.A(clknet_leaf_28_clk_i_regs));
 sg13g2_buf_16 clkload35 (.A(clknet_3_1_0__06563_));
 sg13g2_buf_16 clkload36 (.A(clknet_3_3_0__06563_));
 sg13g2_buf_16 clkload37 (.A(clknet_3_5_0__06563_));
 sg13g2_buf_16 clkload38 (.A(clknet_3_7_0__06563_));
 sg13g2_buf_16 clkload39 (.A(clknet_leaf_0__06563_));
 sg13g2_inv_4 clkload4 (.A(clknet_leaf_46_clk_i_regs));
 sg13g2_inv_2 clkload40 (.A(clknet_leaf_48__06563_));
 sg13g2_buf_8 clkload41 (.A(clknet_leaf_49__06563_));
 sg13g2_inv_1 clkload42 (.A(clknet_leaf_50__06563_));
 sg13g2_buf_8 clkload43 (.A(clknet_leaf_51__06563_));
 sg13g2_buf_8 clkload44 (.A(clknet_leaf_34__06563_));
 sg13g2_buf_8 clkload45 (.A(clknet_leaf_35__06563_));
 sg13g2_inv_8 clkload46 (.A(clknet_leaf_37__06563_));
 sg13g2_inv_1 clkload47 (.A(clknet_leaf_39__06563_));
 sg13g2_inv_8 clkload48 (.A(clknet_leaf_1__06563_));
 sg13g2_inv_4 clkload49 (.A(clknet_leaf_2__06563_));
 sg13g2_inv_2 clkload5 (.A(clknet_leaf_47_clk_i_regs));
 sg13g2_inv_8 clkload50 (.A(clknet_leaf_3__06563_));
 sg13g2_inv_16 clkload51 (.A(clknet_leaf_4__06563_));
 sg13g2_buf_8 clkload52 (.A(clknet_leaf_44__06563_));
 sg13g2_inv_8 clkload53 (.A(clknet_leaf_5__06563_));
 sg13g2_buf_8 clkload54 (.A(clknet_leaf_21__06563_));
 sg13g2_inv_8 clkload55 (.A(clknet_leaf_40__06563_));
 sg13g2_buf_16 clkload56 (.A(clknet_leaf_41__06563_));
 sg13g2_buf_16 clkload57 (.A(clknet_leaf_45__06563_));
 sg13g2_inv_2 clkload58 (.A(clknet_leaf_27__06563_));
 sg13g2_inv_2 clkload59 (.A(clknet_leaf_28__06563_));
 sg13g2_inv_16 clkload6 (.A(clknet_leaf_48_clk_i_regs));
 sg13g2_inv_1 clkload60 (.A(clknet_leaf_31__06563_));
 sg13g2_buf_16 clkload61 (.A(clknet_leaf_32__06563_));
 sg13g2_inv_1 clkload62 (.A(clknet_leaf_33__06563_));
 sg13g2_inv_4 clkload63 (.A(clknet_leaf_17__06563_));
 sg13g2_inv_1 clkload64 (.A(clknet_leaf_22__06563_));
 sg13g2_inv_4 clkload65 (.A(clknet_leaf_23__06563_));
 sg13g2_buf_8 clkload66 (.A(clknet_leaf_25__06563_));
 sg13g2_inv_1 clkload67 (.A(clknet_leaf_29__06563_));
 sg13g2_inv_8 clkload68 (.A(clknet_leaf_6__06563_));
 sg13g2_buf_16 clkload69 (.A(clknet_leaf_7__06563_));
 sg13g2_inv_1 clkload7 (.A(clknet_leaf_2_clk_i_regs));
 sg13g2_inv_4 clkload70 (.A(clknet_leaf_8__06563_));
 sg13g2_buf_16 clkload71 (.A(clknet_leaf_9__06563_));
 sg13g2_buf_16 clkload72 (.A(clknet_leaf_10__06563_));
 sg13g2_inv_8 clkload73 (.A(clknet_leaf_19__06563_));
 sg13g2_inv_4 clkload74 (.A(clknet_leaf_12__06563_));
 sg13g2_buf_16 clkload75 (.A(clknet_leaf_13__06563_));
 sg13g2_inv_2 clkload76 (.A(clknet_leaf_14__06563_));
 sg13g2_buf_8 clkload77 (.A(clknet_leaf_16__06563_));
 sg13g2_buf_8 clkload78 (.A(clknet_leaf_18__06563_));
 sg13g2_inv_8 clkload8 (.A(clknet_leaf_3_clk_i_regs));
 sg13g2_inv_4 clkload9 (.A(clknet_leaf_5_clk_i_regs));
 sg13g2_dfrbpq_1 \core_busy_q$_DFF_PN0_  (.RESET_B(net8242),
    .D(_15423_),
    .Q(core_busy_q),
    .CLK(clknet_leaf_38_clk_i_regs));
 sg13g2_dllrq_1 \core_clock_gate_i.en_latch$_DLATCH_N_  (.D(_15420_),
    .GATE_N(clknet_leaf_38_clk_i_regs),
    .RESET_B(net15),
    .Q(\core_clock_gate_i.en_latch ));
 sg13g2_tiehi \core_clock_gate_i.en_latch$_DLATCH_N__16  (.L_HI(net15));
 sg13g2_dfrbpq_1 \cs_registers_i.mcountinhibit_q[0]$_DFFE_PN0P_  (.RESET_B(net8174),
    .D(_15418_),
    .Q(_00112_),
    .CLK(clknet_leaf_22__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.mcountinhibit_q[2]$_DFFE_PN0P_  (.RESET_B(net8252),
    .D(_15416_),
    .Q(_00113_),
    .CLK(clknet_leaf_22__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.mcycle_counter_i.counter_val_o[0]$_DFFE_PN0P_  (.RESET_B(net8172),
    .D(_15414_),
    .Q(_00114_),
    .CLK(clknet_leaf_18__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.mcycle_counter_i.counter_val_o[10]$_DFFE_PN0P_  (.RESET_B(net8204),
    .D(_15410_),
    .Q(_00115_),
    .CLK(clknet_leaf_12__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.mcycle_counter_i.counter_val_o[11]$_DFFE_PN0P_  (.RESET_B(net8198),
    .D(_15405_),
    .Q(_00116_),
    .CLK(clknet_leaf_12__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.mcycle_counter_i.counter_val_o[12]$_DFFE_PN0P_  (.RESET_B(net8204),
    .D(_15402_),
    .Q(_00117_),
    .CLK(clknet_leaf_12__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.mcycle_counter_i.counter_val_o[13]$_DFFE_PN0P_  (.RESET_B(net8198),
    .D(_15394_),
    .Q(_00118_),
    .CLK(clknet_leaf_12__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.mcycle_counter_i.counter_val_o[14]$_DFFE_PN0P_  (.RESET_B(net8199),
    .D(_15388_),
    .Q(_00119_),
    .CLK(clknet_leaf_12__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.mcycle_counter_i.counter_val_o[15]$_DFFE_PN0P_  (.RESET_B(net8199),
    .D(_15385_),
    .Q(_00120_),
    .CLK(clknet_leaf_13__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.mcycle_counter_i.counter_val_o[16]$_DFFE_PN0P_  (.RESET_B(net8199),
    .D(_15381_),
    .Q(_00121_),
    .CLK(clknet_leaf_13__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.mcycle_counter_i.counter_val_o[17]$_DFFE_PN0P_  (.RESET_B(net8202),
    .D(_15377_),
    .Q(_00122_),
    .CLK(clknet_leaf_16__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.mcycle_counter_i.counter_val_o[18]$_DFFE_PN0P_  (.RESET_B(net8203),
    .D(_15373_),
    .Q(_00123_),
    .CLK(clknet_leaf_13__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.mcycle_counter_i.counter_val_o[19]$_DFFE_PN0P_  (.RESET_B(net8203),
    .D(_15364_),
    .Q(_00124_),
    .CLK(clknet_leaf_16__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.mcycle_counter_i.counter_val_o[1]$_DFFE_PN0P_  (.RESET_B(net8173),
    .D(_15360_),
    .Q(_00125_),
    .CLK(clknet_leaf_18__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.mcycle_counter_i.counter_val_o[20]$_DFFE_PN0P_  (.RESET_B(net8203),
    .D(_15356_),
    .Q(_00126_),
    .CLK(clknet_leaf_16__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.mcycle_counter_i.counter_val_o[21]$_DFFE_PN0P_  (.RESET_B(net8203),
    .D(_15352_),
    .Q(_00127_),
    .CLK(clknet_leaf_17__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.mcycle_counter_i.counter_val_o[22]$_DFFE_PN0P_  (.RESET_B(net8203),
    .D(_15349_),
    .Q(_00128_),
    .CLK(clknet_leaf_17__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.mcycle_counter_i.counter_val_o[23]$_DFFE_PN0P_  (.RESET_B(net8203),
    .D(_15344_),
    .Q(_00129_),
    .CLK(clknet_leaf_17__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.mcycle_counter_i.counter_val_o[24]$_DFFE_PN0P_  (.RESET_B(net8194),
    .D(_15341_),
    .Q(_00130_),
    .CLK(clknet_leaf_17__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.mcycle_counter_i.counter_val_o[25]$_DFFE_PN0P_  (.RESET_B(net8201),
    .D(_15336_),
    .Q(_00131_),
    .CLK(clknet_leaf_17__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.mcycle_counter_i.counter_val_o[26]$_DFFE_PN0P_  (.RESET_B(net8201),
    .D(_15332_),
    .Q(_00132_),
    .CLK(clknet_leaf_17__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.mcycle_counter_i.counter_val_o[27]$_DFFE_PN0P_  (.RESET_B(net8187),
    .D(_15315_),
    .Q(_00133_),
    .CLK(clknet_leaf_18__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.mcycle_counter_i.counter_val_o[28]$_DFFE_PN0P_  (.RESET_B(net8187),
    .D(_15312_),
    .Q(_00134_),
    .CLK(clknet_leaf_18__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.mcycle_counter_i.counter_val_o[29]$_DFFE_PN0P_  (.RESET_B(net8187),
    .D(_15307_),
    .Q(_00135_),
    .CLK(clknet_leaf_18__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.mcycle_counter_i.counter_val_o[2]$_DFFE_PN0P_  (.RESET_B(net8173),
    .D(_15303_),
    .Q(_00136_),
    .CLK(clknet_leaf_18__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.mcycle_counter_i.counter_val_o[30]$_DFFE_PN0P_  (.RESET_B(net8172),
    .D(_15299_),
    .Q(_00137_),
    .CLK(clknet_leaf_18__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.mcycle_counter_i.counter_val_o[31]$_DFFE_PN0P_  (.RESET_B(net8172),
    .D(_15291_),
    .Q(_00138_),
    .CLK(clknet_leaf_18__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.mcycle_counter_i.counter_val_o[32]$_DFFE_PN0P_  (.RESET_B(net8181),
    .D(_15287_),
    .Q(_00139_),
    .CLK(clknet_leaf_18__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.mcycle_counter_i.counter_val_o[33]$_DFFE_PN0P_  (.RESET_B(net8181),
    .D(_15282_),
    .Q(_00140_),
    .CLK(clknet_leaf_18__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.mcycle_counter_i.counter_val_o[34]$_DFFE_PN0P_  (.RESET_B(net8181),
    .D(_15272_),
    .Q(_00141_),
    .CLK(clknet_leaf_17__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.mcycle_counter_i.counter_val_o[35]$_DFFE_PN0P_  (.RESET_B(net8181),
    .D(_15269_),
    .Q(_00142_),
    .CLK(clknet_leaf_17__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.mcycle_counter_i.counter_val_o[36]$_DFFE_PN0P_  (.RESET_B(net8181),
    .D(_15263_),
    .Q(_00143_),
    .CLK(clknet_leaf_15__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.mcycle_counter_i.counter_val_o[37]$_DFFE_PN0P_  (.RESET_B(net8169),
    .D(_15260_),
    .Q(_00144_),
    .CLK(clknet_leaf_14__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.mcycle_counter_i.counter_val_o[38]$_DFFE_PN0P_  (.RESET_B(net8169),
    .D(_15256_),
    .Q(_00145_),
    .CLK(clknet_leaf_15__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.mcycle_counter_i.counter_val_o[39]$_DFFE_PN0P_  (.RESET_B(net8173),
    .D(_15252_),
    .Q(_00146_),
    .CLK(clknet_leaf_15__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.mcycle_counter_i.counter_val_o[3]$_DFFE_PN0P_  (.RESET_B(net8168),
    .D(_15248_),
    .Q(_00147_),
    .CLK(clknet_leaf_15__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.mcycle_counter_i.counter_val_o[40]$_DFFE_PN0P_  (.RESET_B(net8169),
    .D(_15244_),
    .Q(_00148_),
    .CLK(clknet_leaf_15__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.mcycle_counter_i.counter_val_o[41]$_DFFE_PN0P_  (.RESET_B(net8193),
    .D(_15240_),
    .Q(_00149_),
    .CLK(clknet_leaf_14__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.mcycle_counter_i.counter_val_o[42]$_DFFE_PN0P_  (.RESET_B(net8193),
    .D(_15235_),
    .Q(_00150_),
    .CLK(clknet_leaf_14__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.mcycle_counter_i.counter_val_o[43]$_DFFE_PN0P_  (.RESET_B(net8205),
    .D(_15228_),
    .Q(_00151_),
    .CLK(clknet_leaf_13__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.mcycle_counter_i.counter_val_o[44]$_DFFE_PN0P_  (.RESET_B(net8195),
    .D(_15221_),
    .Q(_00152_),
    .CLK(clknet_leaf_13__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.mcycle_counter_i.counter_val_o[45]$_DFFE_PN0P_  (.RESET_B(net8205),
    .D(_15215_),
    .Q(_00153_),
    .CLK(clknet_leaf_13__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.mcycle_counter_i.counter_val_o[46]$_DFFE_PN0P_  (.RESET_B(net8198),
    .D(_15209_),
    .Q(_00154_),
    .CLK(clknet_leaf_13__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.mcycle_counter_i.counter_val_o[47]$_DFFE_PN0P_  (.RESET_B(net8199),
    .D(_15201_),
    .Q(_00155_),
    .CLK(clknet_leaf_13__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.mcycle_counter_i.counter_val_o[48]$_DFFE_PN0P_  (.RESET_B(net8199),
    .D(_15197_),
    .Q(_00156_),
    .CLK(clknet_leaf_13__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.mcycle_counter_i.counter_val_o[49]$_DFFE_PN0P_  (.RESET_B(net8199),
    .D(_15192_),
    .Q(_00157_),
    .CLK(clknet_leaf_13__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.mcycle_counter_i.counter_val_o[4]$_DFFE_PN0P_  (.RESET_B(net8168),
    .D(_15188_),
    .Q(_00158_),
    .CLK(clknet_leaf_15__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.mcycle_counter_i.counter_val_o[50]$_DFFE_PN0P_  (.RESET_B(net8202),
    .D(_15184_),
    .Q(_00159_),
    .CLK(clknet_leaf_16__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.mcycle_counter_i.counter_val_o[51]$_DFFE_PN0P_  (.RESET_B(net8202),
    .D(_15180_),
    .Q(_00160_),
    .CLK(clknet_leaf_16__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.mcycle_counter_i.counter_val_o[52]$_DFFE_PN0P_  (.RESET_B(net8194),
    .D(_15172_),
    .Q(_00161_),
    .CLK(clknet_leaf_16__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.mcycle_counter_i.counter_val_o[53]$_DFFE_PN0P_  (.RESET_B(net8205),
    .D(_15167_),
    .Q(_00162_),
    .CLK(clknet_leaf_17__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.mcycle_counter_i.counter_val_o[54]$_DFFE_PN0P_  (.RESET_B(net8196),
    .D(_15161_),
    .Q(_00163_),
    .CLK(clknet_leaf_17__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.mcycle_counter_i.counter_val_o[55]$_DFFE_PN0P_  (.RESET_B(net8196),
    .D(_15157_),
    .Q(_00164_),
    .CLK(clknet_leaf_17__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.mcycle_counter_i.counter_val_o[56]$_DFFE_PN0P_  (.RESET_B(net8196),
    .D(_15151_),
    .Q(_00165_),
    .CLK(clknet_leaf_17__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.mcycle_counter_i.counter_val_o[57]$_DFFE_PN0P_  (.RESET_B(net8196),
    .D(_15144_),
    .Q(_00166_),
    .CLK(clknet_leaf_17__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.mcycle_counter_i.counter_val_o[58]$_DFFE_PN0P_  (.RESET_B(net8196),
    .D(_15140_),
    .Q(_00167_),
    .CLK(clknet_leaf_17__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.mcycle_counter_i.counter_val_o[59]$_DFFE_PN0P_  (.RESET_B(net8187),
    .D(_15136_),
    .Q(_00168_),
    .CLK(clknet_leaf_18__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.mcycle_counter_i.counter_val_o[5]$_DFFE_PN0P_  (.RESET_B(net8168),
    .D(_15131_),
    .Q(_00169_),
    .CLK(clknet_leaf_15__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.mcycle_counter_i.counter_val_o[60]$_DFFE_PN0P_  (.RESET_B(net8187),
    .D(_15122_),
    .Q(_00170_),
    .CLK(clknet_leaf_23__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.mcycle_counter_i.counter_val_o[61]$_DFFE_PN0P_  (.RESET_B(net8172),
    .D(_15117_),
    .Q(_00171_),
    .CLK(clknet_leaf_18__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.mcycle_counter_i.counter_val_o[62]$_DFFE_PN0P_  (.RESET_B(net8172),
    .D(_15112_),
    .Q(_00172_),
    .CLK(clknet_leaf_18__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.mcycle_counter_i.counter_val_o[63]$_DFFE_PN0P_  (.RESET_B(net8172),
    .D(_15106_),
    .Q(_00173_),
    .CLK(clknet_leaf_18__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.mcycle_counter_i.counter_val_o[6]$_DFFE_PN0P_  (.RESET_B(net8169),
    .D(_15046_),
    .Q(_00174_),
    .CLK(clknet_leaf_15__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.mcycle_counter_i.counter_val_o[7]$_DFFE_PN0P_  (.RESET_B(net8193),
    .D(_15041_),
    .Q(_00175_),
    .CLK(clknet_leaf_14__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.mcycle_counter_i.counter_val_o[8]$_DFFE_PN0P_  (.RESET_B(net8193),
    .D(_15035_),
    .Q(_00176_),
    .CLK(clknet_leaf_14__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.mcycle_counter_i.counter_val_o[9]$_DFFE_PN0P_  (.RESET_B(net8198),
    .D(_15029_),
    .Q(_00177_),
    .CLK(clknet_leaf_12__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.minstret_counter_i.counter_val_o[0]$_DFFE_PN0P_  (.RESET_B(net8173),
    .D(_15005_),
    .Q(_00178_),
    .CLK(clknet_leaf_18__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.minstret_counter_i.counter_val_o[10]$_DFFE_PN0P_  (.RESET_B(net8199),
    .D(_15000_),
    .Q(_00179_),
    .CLK(clknet_leaf_12__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.minstret_counter_i.counter_val_o[11]$_DFFE_PN0P_  (.RESET_B(net8204),
    .D(_14996_),
    .Q(_00180_),
    .CLK(clknet_leaf_12__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.minstret_counter_i.counter_val_o[12]$_DFFE_PN0P_  (.RESET_B(net8204),
    .D(_14990_),
    .Q(_00181_),
    .CLK(clknet_leaf_12__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.minstret_counter_i.counter_val_o[13]$_DFFE_PN0P_  (.RESET_B(net8204),
    .D(_14986_),
    .Q(_00182_),
    .CLK(clknet_leaf_12__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.minstret_counter_i.counter_val_o[14]$_DFFE_PN0P_  (.RESET_B(net8197),
    .D(_14976_),
    .Q(_00183_),
    .CLK(clknet_leaf_13__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.minstret_counter_i.counter_val_o[15]$_DFFE_PN0P_  (.RESET_B(net8197),
    .D(_14971_),
    .Q(_00184_),
    .CLK(clknet_leaf_16__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.minstret_counter_i.counter_val_o[16]$_DFFE_PN0P_  (.RESET_B(net8202),
    .D(_14966_),
    .Q(_00185_),
    .CLK(clknet_leaf_16__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.minstret_counter_i.counter_val_o[17]$_DFFE_PN0P_  (.RESET_B(net8202),
    .D(_14961_),
    .Q(_00186_),
    .CLK(clknet_leaf_16__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.minstret_counter_i.counter_val_o[18]$_DFFE_PN0P_  (.RESET_B(net8202),
    .D(_14956_),
    .Q(_00187_),
    .CLK(clknet_leaf_16__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.minstret_counter_i.counter_val_o[19]$_DFFE_PN0P_  (.RESET_B(net8201),
    .D(_14951_),
    .Q(_00188_),
    .CLK(clknet_leaf_17__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.minstret_counter_i.counter_val_o[1]$_DFFE_PN0P_  (.RESET_B(net8173),
    .D(_14946_),
    .Q(_00189_),
    .CLK(clknet_leaf_18__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.minstret_counter_i.counter_val_o[20]$_DFFE_PN0P_  (.RESET_B(net8201),
    .D(_14941_),
    .Q(_00190_),
    .CLK(clknet_leaf_17__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.minstret_counter_i.counter_val_o[21]$_DFFE_PN0P_  (.RESET_B(net8201),
    .D(_14937_),
    .Q(_00191_),
    .CLK(clknet_leaf_23__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.minstret_counter_i.counter_val_o[22]$_DFFE_PN0P_  (.RESET_B(net8201),
    .D(_14931_),
    .Q(_00192_),
    .CLK(clknet_leaf_23__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.minstret_counter_i.counter_val_o[23]$_DFFE_PN0P_  (.RESET_B(net8200),
    .D(_14926_),
    .Q(_00193_),
    .CLK(clknet_leaf_23__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.minstret_counter_i.counter_val_o[24]$_DFFE_PN0P_  (.RESET_B(net8200),
    .D(_14922_),
    .Q(_00194_),
    .CLK(clknet_leaf_23__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.minstret_counter_i.counter_val_o[25]$_DFFE_PN0P_  (.RESET_B(net8200),
    .D(_14918_),
    .Q(_00195_),
    .CLK(clknet_leaf_23__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.minstret_counter_i.counter_val_o[26]$_DFFE_PN0P_  (.RESET_B(net8201),
    .D(_14902_),
    .Q(_00196_),
    .CLK(clknet_leaf_23__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.minstret_counter_i.counter_val_o[27]$_DFFE_PN0P_  (.RESET_B(net8187),
    .D(_14889_),
    .Q(_00197_),
    .CLK(clknet_leaf_23__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.minstret_counter_i.counter_val_o[28]$_DFFE_PN0P_  (.RESET_B(net8182),
    .D(_14885_),
    .Q(_00198_),
    .CLK(clknet_leaf_23__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.minstret_counter_i.counter_val_o[29]$_DFFE_PN0P_  (.RESET_B(net8182),
    .D(_14881_),
    .Q(_00199_),
    .CLK(clknet_leaf_23__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.minstret_counter_i.counter_val_o[2]$_DFFE_PN0P_  (.RESET_B(net8173),
    .D(_14875_),
    .Q(_00200_),
    .CLK(clknet_leaf_18__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.minstret_counter_i.counter_val_o[30]$_DFFE_PN0P_  (.RESET_B(net8182),
    .D(_14870_),
    .Q(_00201_),
    .CLK(clknet_leaf_23__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.minstret_counter_i.counter_val_o[31]$_DFFE_PN0P_  (.RESET_B(net8182),
    .D(_14866_),
    .Q(_00202_),
    .CLK(clknet_leaf_24__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.minstret_counter_i.counter_val_o[32]$_DFFE_PN0P_  (.RESET_B(net8194),
    .D(_14851_),
    .Q(_00203_),
    .CLK(clknet_leaf_16__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.minstret_counter_i.counter_val_o[33]$_DFFE_PN0P_  (.RESET_B(net8194),
    .D(_14847_),
    .Q(_00204_),
    .CLK(clknet_leaf_17__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.minstret_counter_i.counter_val_o[34]$_DFFE_PN0P_  (.RESET_B(net8194),
    .D(_14842_),
    .Q(_00205_),
    .CLK(clknet_leaf_16__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.minstret_counter_i.counter_val_o[35]$_DFFE_PN0P_  (.RESET_B(net8181),
    .D(_14835_),
    .Q(_00206_),
    .CLK(clknet_leaf_15__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.minstret_counter_i.counter_val_o[36]$_DFFE_PN0P_  (.RESET_B(net8181),
    .D(_14830_),
    .Q(_00207_),
    .CLK(clknet_leaf_15__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.minstret_counter_i.counter_val_o[37]$_DFFE_PN0P_  (.RESET_B(net8194),
    .D(_14823_),
    .Q(_00208_),
    .CLK(clknet_leaf_15__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.minstret_counter_i.counter_val_o[38]$_DFFE_PN0P_  (.RESET_B(net8195),
    .D(_14818_),
    .Q(_00209_),
    .CLK(clknet_leaf_15__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.minstret_counter_i.counter_val_o[39]$_DFFE_PN0P_  (.RESET_B(net8195),
    .D(_14815_),
    .Q(_00210_),
    .CLK(clknet_leaf_15__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.minstret_counter_i.counter_val_o[3]$_DFFE_PN0P_  (.RESET_B(net8173),
    .D(_14809_),
    .Q(_00211_),
    .CLK(clknet_leaf_19__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.minstret_counter_i.counter_val_o[40]$_DFFE_PN0P_  (.RESET_B(net8195),
    .D(_14804_),
    .Q(_00212_),
    .CLK(clknet_leaf_15__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.minstret_counter_i.counter_val_o[41]$_DFFE_PN0P_  (.RESET_B(net8197),
    .D(_14793_),
    .Q(_00213_),
    .CLK(clknet_leaf_13__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.minstret_counter_i.counter_val_o[42]$_DFFE_PN0P_  (.RESET_B(net8197),
    .D(_14788_),
    .Q(_00214_),
    .CLK(clknet_leaf_13__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.minstret_counter_i.counter_val_o[43]$_DFFE_PN0P_  (.RESET_B(net8197),
    .D(_14783_),
    .Q(_00215_),
    .CLK(clknet_leaf_13__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.minstret_counter_i.counter_val_o[44]$_DFFE_PN0P_  (.RESET_B(net8198),
    .D(_14778_),
    .Q(_00216_),
    .CLK(clknet_leaf_12__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.minstret_counter_i.counter_val_o[45]$_DFFE_PN0P_  (.RESET_B(net8181),
    .D(_14771_),
    .Q(_00217_),
    .CLK(clknet_leaf_15__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.minstret_counter_i.counter_val_o[46]$_DFFE_PN0P_  (.RESET_B(net8195),
    .D(_14765_),
    .Q(_00218_),
    .CLK(clknet_leaf_13__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.minstret_counter_i.counter_val_o[47]$_DFFE_PN0P_  (.RESET_B(net8197),
    .D(_14756_),
    .Q(_00219_),
    .CLK(clknet_leaf_16__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.minstret_counter_i.counter_val_o[48]$_DFFE_PN0P_  (.RESET_B(net8197),
    .D(_14752_),
    .Q(_00220_),
    .CLK(clknet_leaf_16__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.minstret_counter_i.counter_val_o[49]$_DFFE_PN0P_  (.RESET_B(net8197),
    .D(_14747_),
    .Q(_00221_),
    .CLK(clknet_leaf_16__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.minstret_counter_i.counter_val_o[4]$_DFFE_PN0P_  (.RESET_B(net8168),
    .D(_14743_),
    .Q(_00222_),
    .CLK(clknet_leaf_19__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.minstret_counter_i.counter_val_o[50]$_DFFE_PN0P_  (.RESET_B(net8194),
    .D(_14739_),
    .Q(_00223_),
    .CLK(clknet_leaf_16__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.minstret_counter_i.counter_val_o[51]$_DFFE_PN0P_  (.RESET_B(net8194),
    .D(_14735_),
    .Q(_00224_),
    .CLK(clknet_leaf_16__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.minstret_counter_i.counter_val_o[52]$_DFFE_PN0P_  (.RESET_B(net8196),
    .D(_14731_),
    .Q(_00225_),
    .CLK(clknet_leaf_17__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.minstret_counter_i.counter_val_o[53]$_DFFE_PN0P_  (.RESET_B(net8196),
    .D(_14726_),
    .Q(_00226_),
    .CLK(clknet_leaf_23__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.minstret_counter_i.counter_val_o[54]$_DFFE_PN0P_  (.RESET_B(net8196),
    .D(_14719_),
    .Q(_00227_),
    .CLK(clknet_leaf_23__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.minstret_counter_i.counter_val_o[55]$_DFFE_PN0P_  (.RESET_B(net8201),
    .D(_14712_),
    .Q(_00228_),
    .CLK(clknet_leaf_23__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.minstret_counter_i.counter_val_o[56]$_DFFE_PN0P_  (.RESET_B(net8200),
    .D(_14707_),
    .Q(_00229_),
    .CLK(clknet_leaf_23__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.minstret_counter_i.counter_val_o[57]$_DFFE_PN0P_  (.RESET_B(net8182),
    .D(_14702_),
    .Q(_00230_),
    .CLK(clknet_leaf_24__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.minstret_counter_i.counter_val_o[58]$_DFFE_PN0P_  (.RESET_B(net8182),
    .D(_14694_),
    .Q(_00231_),
    .CLK(clknet_leaf_23__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.minstret_counter_i.counter_val_o[59]$_DFFE_PN0P_  (.RESET_B(net8182),
    .D(_14689_),
    .Q(_00232_),
    .CLK(clknet_leaf_24__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.minstret_counter_i.counter_val_o[5]$_DFFE_PN0P_  (.RESET_B(net8168),
    .D(_14685_),
    .Q(_00233_),
    .CLK(clknet_leaf_15__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.minstret_counter_i.counter_val_o[60]$_DFFE_PN0P_  (.RESET_B(net8182),
    .D(_14681_),
    .Q(_00234_),
    .CLK(clknet_leaf_24__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.minstret_counter_i.counter_val_o[61]$_DFFE_PN0P_  (.RESET_B(net8172),
    .D(_14676_),
    .Q(_00235_),
    .CLK(clknet_leaf_23__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.minstret_counter_i.counter_val_o[62]$_DFFE_PN0P_  (.RESET_B(net8176),
    .D(_14672_),
    .Q(_00236_),
    .CLK(clknet_leaf_22__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.minstret_counter_i.counter_val_o[63]$_DFFE_PN0P_  (.RESET_B(net8172),
    .D(_14667_),
    .Q(_00237_),
    .CLK(clknet_leaf_22__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.minstret_counter_i.counter_val_o[6]$_DFFE_PN0P_  (.RESET_B(net8169),
    .D(_14606_),
    .Q(_00238_),
    .CLK(clknet_leaf_15__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.minstret_counter_i.counter_val_o[7]$_DFFE_PN0P_  (.RESET_B(net8195),
    .D(_14598_),
    .Q(_00239_),
    .CLK(clknet_leaf_15__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.minstret_counter_i.counter_val_o[8]$_DFFE_PN0P_  (.RESET_B(net8195),
    .D(_14591_),
    .Q(_00240_),
    .CLK(clknet_leaf_15__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.minstret_counter_i.counter_val_o[9]$_DFFE_PN0P_  (.RESET_B(net8199),
    .D(_14587_),
    .Q(_00241_),
    .CLK(clknet_leaf_12__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.priv_mode_id_o[0]$_DFFE_PN1P_  (.RESET_B(net8245),
    .D(_14557_),
    .Q(_00242_),
    .CLK(clknet_leaf_21__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.priv_mode_id_o[1]$_DFFE_PN1P_  (.RESET_B(net8245),
    .D(_14553_),
    .Q(_00243_),
    .CLK(clknet_leaf_21__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dcsr_csr.rd_data_o[0]$_DFFE_PN1P_  (.RESET_B(net8248),
    .D(_14549_),
    .Q(_00000_),
    .CLK(clknet_leaf_21__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dcsr_csr.rd_data_o[11]$_DFFE_PN0P_  (.RESET_B(net8179),
    .D(_14547_),
    .Q(_00244_),
    .CLK(clknet_leaf_28__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dcsr_csr.rd_data_o[12]$_DFFE_PN0P_  (.RESET_B(net8178),
    .D(_14545_),
    .Q(\cs_registers_i.debug_ebreaku_o ),
    .CLK(clknet_leaf_28__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dcsr_csr.rd_data_o[13]$_DFFE_PN0P_  (.RESET_B(net8280),
    .D(_14542_),
    .Q(_00245_),
    .CLK(clknet_leaf_28__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dcsr_csr.rd_data_o[15]$_DFFE_PN0P_  (.RESET_B(net8249),
    .D(_14539_),
    .Q(\cs_registers_i.debug_ebreakm_o ),
    .CLK(clknet_leaf_21__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dcsr_csr.rd_data_o[1]$_DFFE_PN1P_  (.RESET_B(net8248),
    .D(_14537_),
    .Q(_00001_),
    .CLK(clknet_leaf_21__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dcsr_csr.rd_data_o[2]$_DFFE_PN0P_  (.RESET_B(net8249),
    .D(_14533_),
    .Q(\cs_registers_i.debug_single_step_o ),
    .CLK(clknet_leaf_26__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dcsr_csr.rd_data_o[6]$_DFFE_PN0P_  (.RESET_B(net8267),
    .D(_14530_),
    .Q(_00246_),
    .CLK(clknet_leaf_26__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dcsr_csr.rd_data_o[7]$_DFFE_PN0P_  (.RESET_B(net8267),
    .D(_14529_),
    .Q(_00247_),
    .CLK(clknet_leaf_27__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dcsr_csr.rd_data_o[8]$_DFFE_PN0P_  (.RESET_B(net8267),
    .D(_14526_),
    .Q(_00248_),
    .CLK(clknet_leaf_27__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_depc_csr.rd_data_o[10]$_DFFE_PN0P_  (.RESET_B(net8258),
    .D(_14524_),
    .Q(_00249_),
    .CLK(clknet_leaf_39__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_depc_csr.rd_data_o[11]$_DFFE_PN0P_  (.RESET_B(net8259),
    .D(_14521_),
    .Q(_00250_),
    .CLK(clknet_leaf_33__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_depc_csr.rd_data_o[12]$_DFFE_PN0P_  (.RESET_B(net8258),
    .D(_14518_),
    .Q(_00251_),
    .CLK(clknet_leaf_39__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_depc_csr.rd_data_o[13]$_DFFE_PN0P_  (.RESET_B(net8258),
    .D(_14515_),
    .Q(_00252_),
    .CLK(clknet_leaf_39__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_depc_csr.rd_data_o[14]$_DFFE_PN0P_  (.RESET_B(net8258),
    .D(_14512_),
    .Q(_00253_),
    .CLK(clknet_leaf_39__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_depc_csr.rd_data_o[15]$_DFFE_PN0P_  (.RESET_B(net8260),
    .D(_14508_),
    .Q(_00254_),
    .CLK(clknet_leaf_34__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_depc_csr.rd_data_o[16]$_DFFE_PN0P_  (.RESET_B(net8259),
    .D(_14504_),
    .Q(_00255_),
    .CLK(clknet_leaf_33__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_depc_csr.rd_data_o[17]$_DFFE_PN0P_  (.RESET_B(net8264),
    .D(_14501_),
    .Q(_00256_),
    .CLK(clknet_leaf_32__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_depc_csr.rd_data_o[18]$_DFFE_PN0P_  (.RESET_B(net8263),
    .D(_14498_),
    .Q(_00257_),
    .CLK(clknet_leaf_32__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_depc_csr.rd_data_o[19]$_DFFE_PN0P_  (.RESET_B(net8268),
    .D(_14495_),
    .Q(_00258_),
    .CLK(clknet_leaf_33__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_depc_csr.rd_data_o[1]$_DFFE_PN0P_  (.RESET_B(net8245),
    .D(_14492_),
    .Q(_00259_),
    .CLK(clknet_leaf_21__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_depc_csr.rd_data_o[20]$_DFFE_PN0P_  (.RESET_B(net8260),
    .D(_14489_),
    .Q(_00260_),
    .CLK(clknet_leaf_34__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_depc_csr.rd_data_o[21]$_DFFE_PN0P_  (.RESET_B(net8260),
    .D(_14486_),
    .Q(_00261_),
    .CLK(clknet_leaf_33__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_depc_csr.rd_data_o[22]$_DFFE_PN0P_  (.RESET_B(net8281),
    .D(_14483_),
    .Q(_00262_),
    .CLK(clknet_leaf_27__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_depc_csr.rd_data_o[23]$_DFFE_PN0P_  (.RESET_B(net8281),
    .D(_14480_),
    .Q(_00263_),
    .CLK(clknet_leaf_27__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_depc_csr.rd_data_o[24]$_DFFE_PN0P_  (.RESET_B(net8269),
    .D(_14477_),
    .Q(_00264_),
    .CLK(clknet_leaf_33__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_depc_csr.rd_data_o[25]$_DFFE_PN0P_  (.RESET_B(net8268),
    .D(_14473_),
    .Q(_00265_),
    .CLK(clknet_leaf_33__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_depc_csr.rd_data_o[26]$_DFFE_PN0P_  (.RESET_B(net8268),
    .D(_14470_),
    .Q(_00266_),
    .CLK(clknet_leaf_33__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_depc_csr.rd_data_o[27]$_DFFE_PN0P_  (.RESET_B(net8269),
    .D(_14467_),
    .Q(_00267_),
    .CLK(clknet_leaf_33__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_depc_csr.rd_data_o[28]$_DFFE_PN0P_  (.RESET_B(net8263),
    .D(_14464_),
    .Q(_00268_),
    .CLK(clknet_leaf_32__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_depc_csr.rd_data_o[29]$_DFFE_PN0P_  (.RESET_B(net8263),
    .D(_14461_),
    .Q(_00269_),
    .CLK(clknet_leaf_32__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_depc_csr.rd_data_o[2]$_DFFE_PN0P_  (.RESET_B(net8247),
    .D(_14458_),
    .Q(_00270_),
    .CLK(clknet_leaf_21__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_depc_csr.rd_data_o[30]$_DFFE_PN0P_  (.RESET_B(net8263),
    .D(_14455_),
    .Q(_00271_),
    .CLK(clknet_leaf_32__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_depc_csr.rd_data_o[31]$_DFFE_PN0P_  (.RESET_B(net8265),
    .D(_14451_),
    .Q(_00272_),
    .CLK(clknet_leaf_33__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_depc_csr.rd_data_o[3]$_DFFE_PN0P_  (.RESET_B(net8248),
    .D(_14448_),
    .Q(_00273_),
    .CLK(clknet_leaf_21__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_depc_csr.rd_data_o[4]$_DFFE_PN0P_  (.RESET_B(net8248),
    .D(_14444_),
    .Q(_00274_),
    .CLK(clknet_leaf_21__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_depc_csr.rd_data_o[5]$_DFFE_PN0P_  (.RESET_B(net8282),
    .D(_14441_),
    .Q(_00275_),
    .CLK(clknet_leaf_27__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_depc_csr.rd_data_o[6]$_DFFE_PN0P_  (.RESET_B(net8282),
    .D(_14438_),
    .Q(_00276_),
    .CLK(clknet_leaf_27__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_depc_csr.rd_data_o[7]$_DFFE_PN0P_  (.RESET_B(net8266),
    .D(_14435_),
    .Q(_00277_),
    .CLK(clknet_leaf_34__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_depc_csr.rd_data_o[8]$_DFFE_PN0P_  (.RESET_B(net8258),
    .D(_14432_),
    .Q(_00278_),
    .CLK(clknet_leaf_39__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_depc_csr.rd_data_o[9]$_DFFE_PN0P_  (.RESET_B(net8266),
    .D(_14429_),
    .Q(_00279_),
    .CLK(clknet_leaf_34__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dscratch0_csr.rd_data_o[0]$_DFFE_PN0P_  (.RESET_B(net8174),
    .D(_14424_),
    .Q(_00280_),
    .CLK(clknet_leaf_22__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dscratch0_csr.rd_data_o[10]$_DFFE_PN0P_  (.RESET_B(net8179),
    .D(_14422_),
    .Q(_00281_),
    .CLK(clknet_leaf_28__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dscratch0_csr.rd_data_o[11]$_DFFE_PN0P_  (.RESET_B(net8179),
    .D(_14420_),
    .Q(_00282_),
    .CLK(clknet_leaf_29__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dscratch0_csr.rd_data_o[12]$_DFFE_PN0P_  (.RESET_B(net8274),
    .D(_14417_),
    .Q(_00283_),
    .CLK(clknet_leaf_28__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dscratch0_csr.rd_data_o[13]$_DFFE_PN0P_  (.RESET_B(net8273),
    .D(_14415_),
    .Q(_00284_),
    .CLK(clknet_leaf_30__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dscratch0_csr.rd_data_o[14]$_DFFE_PN0P_  (.RESET_B(net8185),
    .D(_14413_),
    .Q(_00285_),
    .CLK(clknet_leaf_28__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dscratch0_csr.rd_data_o[15]$_DFFE_PN0P_  (.RESET_B(net8174),
    .D(_14410_),
    .Q(_00286_),
    .CLK(clknet_leaf_22__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dscratch0_csr.rd_data_o[16]$_DFFE_PN0P_  (.RESET_B(net8278),
    .D(_14408_),
    .Q(_00287_),
    .CLK(clknet_leaf_29__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dscratch0_csr.rd_data_o[17]$_DFFE_PN0P_  (.RESET_B(net8279),
    .D(_14406_),
    .Q(_00288_),
    .CLK(clknet_leaf_29__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dscratch0_csr.rd_data_o[18]$_DFFE_PN0P_  (.RESET_B(net8276),
    .D(_14403_),
    .Q(_00289_),
    .CLK(clknet_leaf_30__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dscratch0_csr.rd_data_o[19]$_DFFE_PN0P_  (.RESET_B(net8277),
    .D(_14401_),
    .Q(_00290_),
    .CLK(clknet_leaf_30__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dscratch0_csr.rd_data_o[1]$_DFFE_PN0P_  (.RESET_B(net8176),
    .D(_14399_),
    .Q(_00291_),
    .CLK(clknet_leaf_24__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dscratch0_csr.rd_data_o[20]$_DFFE_PN0P_  (.RESET_B(net8278),
    .D(_14397_),
    .Q(_00292_),
    .CLK(clknet_leaf_30__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dscratch0_csr.rd_data_o[21]$_DFFE_PN0P_  (.RESET_B(net8185),
    .D(_14394_),
    .Q(_00293_),
    .CLK(clknet_leaf_25__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dscratch0_csr.rd_data_o[22]$_DFFE_PN0P_  (.RESET_B(net8184),
    .D(_14392_),
    .Q(_00294_),
    .CLK(clknet_leaf_25__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dscratch0_csr.rd_data_o[23]$_DFFE_PN0P_  (.RESET_B(net8183),
    .D(_14390_),
    .Q(_00295_),
    .CLK(clknet_leaf_25__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dscratch0_csr.rd_data_o[24]$_DFFE_PN0P_  (.RESET_B(net8183),
    .D(_14388_),
    .Q(_00296_),
    .CLK(clknet_leaf_25__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dscratch0_csr.rd_data_o[25]$_DFFE_PN0P_  (.RESET_B(net8277),
    .D(_14385_),
    .Q(_00297_),
    .CLK(clknet_leaf_29__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dscratch0_csr.rd_data_o[26]$_DFFE_PN0P_  (.RESET_B(net8278),
    .D(_14383_),
    .Q(_00298_),
    .CLK(clknet_leaf_29__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dscratch0_csr.rd_data_o[27]$_DFFE_PN0P_  (.RESET_B(net8179),
    .D(_14381_),
    .Q(_00299_),
    .CLK(clknet_leaf_29__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dscratch0_csr.rd_data_o[28]$_DFFE_PN0P_  (.RESET_B(net8276),
    .D(_14379_),
    .Q(_00300_),
    .CLK(clknet_leaf_30__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dscratch0_csr.rd_data_o[29]$_DFFE_PN0P_  (.RESET_B(net8272),
    .D(_14377_),
    .Q(_00301_),
    .CLK(clknet_leaf_30__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dscratch0_csr.rd_data_o[2]$_DFFE_PN0P_  (.RESET_B(net8177),
    .D(_14375_),
    .Q(_00302_),
    .CLK(clknet_leaf_25__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dscratch0_csr.rd_data_o[30]$_DFFE_PN0P_  (.RESET_B(net8273),
    .D(_14372_),
    .Q(_00303_),
    .CLK(clknet_leaf_30__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dscratch0_csr.rd_data_o[31]$_DFFE_PN0P_  (.RESET_B(net8272),
    .D(_14370_),
    .Q(_00304_),
    .CLK(clknet_leaf_31__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dscratch0_csr.rd_data_o[3]$_DFFE_PN0P_  (.RESET_B(net8176),
    .D(_14368_),
    .Q(_00305_),
    .CLK(clknet_leaf_22__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dscratch0_csr.rd_data_o[4]$_DFFE_PN0P_  (.RESET_B(net8176),
    .D(_14366_),
    .Q(_00306_),
    .CLK(clknet_leaf_22__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dscratch0_csr.rd_data_o[5]$_DFFE_PN0P_  (.RESET_B(net8186),
    .D(_14364_),
    .Q(_00307_),
    .CLK(clknet_leaf_25__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dscratch0_csr.rd_data_o[6]$_DFFE_PN0P_  (.RESET_B(net8180),
    .D(_14362_),
    .Q(_00308_),
    .CLK(clknet_leaf_26__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dscratch0_csr.rd_data_o[7]$_DFFE_PN0P_  (.RESET_B(net8277),
    .D(_14360_),
    .Q(_00309_),
    .CLK(clknet_leaf_29__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dscratch0_csr.rd_data_o[8]$_DFFE_PN0P_  (.RESET_B(net8179),
    .D(_14357_),
    .Q(_00310_),
    .CLK(clknet_leaf_28__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dscratch0_csr.rd_data_o[9]$_DFFE_PN0P_  (.RESET_B(net8273),
    .D(_14355_),
    .Q(_00311_),
    .CLK(clknet_leaf_30__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dscratch1_csr.rd_data_o[0]$_DFFE_PN0P_  (.RESET_B(net8180),
    .D(_14352_),
    .Q(_00312_),
    .CLK(clknet_leaf_24__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dscratch1_csr.rd_data_o[10]$_DFFE_PN0P_  (.RESET_B(net8274),
    .D(_14349_),
    .Q(_00313_),
    .CLK(clknet_leaf_30__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dscratch1_csr.rd_data_o[11]$_DFFE_PN0P_  (.RESET_B(net8275),
    .D(_14347_),
    .Q(_00314_),
    .CLK(clknet_leaf_29__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dscratch1_csr.rd_data_o[12]$_DFFE_PN0P_  (.RESET_B(net8179),
    .D(_14345_),
    .Q(_00315_),
    .CLK(clknet_leaf_28__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dscratch1_csr.rd_data_o[13]$_DFFE_PN0P_  (.RESET_B(net8272),
    .D(_14343_),
    .Q(_00316_),
    .CLK(clknet_leaf_30__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dscratch1_csr.rd_data_o[14]$_DFFE_PN0P_  (.RESET_B(net8185),
    .D(_14341_),
    .Q(_00317_),
    .CLK(clknet_leaf_28__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dscratch1_csr.rd_data_o[15]$_DFFE_PN0P_  (.RESET_B(net8180),
    .D(_14339_),
    .Q(_00318_),
    .CLK(clknet_leaf_24__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dscratch1_csr.rd_data_o[16]$_DFFE_PN0P_  (.RESET_B(net8278),
    .D(_14336_),
    .Q(_00319_),
    .CLK(clknet_leaf_29__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dscratch1_csr.rd_data_o[17]$_DFFE_PN0P_  (.RESET_B(net8276),
    .D(_14334_),
    .Q(_00320_),
    .CLK(clknet_leaf_30__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dscratch1_csr.rd_data_o[18]$_DFFE_PN0P_  (.RESET_B(net8276),
    .D(_14331_),
    .Q(_00321_),
    .CLK(clknet_leaf_31__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dscratch1_csr.rd_data_o[19]$_DFFE_PN0P_  (.RESET_B(net8277),
    .D(_14329_),
    .Q(_00322_),
    .CLK(clknet_leaf_30__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dscratch1_csr.rd_data_o[1]$_DFFE_PN0P_  (.RESET_B(net8175),
    .D(_14327_),
    .Q(_00323_),
    .CLK(clknet_leaf_24__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dscratch1_csr.rd_data_o[20]$_DFFE_PN0P_  (.RESET_B(net8278),
    .D(_14325_),
    .Q(_00324_),
    .CLK(clknet_leaf_29__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dscratch1_csr.rd_data_o[21]$_DFFE_PN0P_  (.RESET_B(net8185),
    .D(_14323_),
    .Q(_00325_),
    .CLK(clknet_leaf_25__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dscratch1_csr.rd_data_o[22]$_DFFE_PN0P_  (.RESET_B(net8183),
    .D(_14321_),
    .Q(_00326_),
    .CLK(clknet_leaf_29__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dscratch1_csr.rd_data_o[23]$_DFFE_PN0P_  (.RESET_B(net8183),
    .D(_14319_),
    .Q(_00327_),
    .CLK(clknet_leaf_25__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dscratch1_csr.rd_data_o[24]$_DFFE_PN0P_  (.RESET_B(net8183),
    .D(_14317_),
    .Q(_00328_),
    .CLK(clknet_leaf_25__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dscratch1_csr.rd_data_o[25]$_DFFE_PN0P_  (.RESET_B(net8277),
    .D(_14315_),
    .Q(_00329_),
    .CLK(clknet_leaf_29__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dscratch1_csr.rd_data_o[26]$_DFFE_PN0P_  (.RESET_B(net8278),
    .D(_14313_),
    .Q(_00330_),
    .CLK(clknet_leaf_29__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dscratch1_csr.rd_data_o[27]$_DFFE_PN0P_  (.RESET_B(net8179),
    .D(_14311_),
    .Q(_00331_),
    .CLK(clknet_leaf_29__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dscratch1_csr.rd_data_o[28]$_DFFE_PN0P_  (.RESET_B(net8276),
    .D(_14309_),
    .Q(_00332_),
    .CLK(clknet_leaf_31__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dscratch1_csr.rd_data_o[29]$_DFFE_PN0P_  (.RESET_B(net8272),
    .D(_14307_),
    .Q(_00333_),
    .CLK(clknet_leaf_31__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dscratch1_csr.rd_data_o[2]$_DFFE_PN0P_  (.RESET_B(net8180),
    .D(_14305_),
    .Q(_00334_),
    .CLK(clknet_leaf_25__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dscratch1_csr.rd_data_o[30]$_DFFE_PN0P_  (.RESET_B(net8272),
    .D(_14303_),
    .Q(_00335_),
    .CLK(clknet_leaf_31__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dscratch1_csr.rd_data_o[31]$_DFFE_PN0P_  (.RESET_B(net8272),
    .D(_14301_),
    .Q(_00336_),
    .CLK(clknet_leaf_31__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dscratch1_csr.rd_data_o[3]$_DFFE_PN0P_  (.RESET_B(net8175),
    .D(_14298_),
    .Q(_00337_),
    .CLK(clknet_leaf_23__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dscratch1_csr.rd_data_o[4]$_DFFE_PN0P_  (.RESET_B(net8176),
    .D(_14296_),
    .Q(_00338_),
    .CLK(clknet_leaf_24__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dscratch1_csr.rd_data_o[5]$_DFFE_PN0P_  (.RESET_B(net8186),
    .D(_14294_),
    .Q(_00339_),
    .CLK(clknet_leaf_25__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dscratch1_csr.rd_data_o[6]$_DFFE_PN0P_  (.RESET_B(net8175),
    .D(_14292_),
    .Q(_00340_),
    .CLK(clknet_leaf_24__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dscratch1_csr.rd_data_o[7]$_DFFE_PN0P_  (.RESET_B(net8275),
    .D(_14289_),
    .Q(_00341_),
    .CLK(clknet_leaf_28__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dscratch1_csr.rd_data_o[8]$_DFFE_PN0P_  (.RESET_B(net8274),
    .D(_14286_),
    .Q(_00342_),
    .CLK(clknet_leaf_29__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_dscratch1_csr.rd_data_o[9]$_DFFE_PN0P_  (.RESET_B(net8274),
    .D(_14284_),
    .Q(_00343_),
    .CLK(clknet_leaf_30__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mcause_csr.rd_data_o[0]$_DFFE_PN0P_  (.RESET_B(net8249),
    .D(_14281_),
    .Q(_00344_),
    .CLK(clknet_leaf_26__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mcause_csr.rd_data_o[1]$_DFFE_PN0P_  (.RESET_B(net8251),
    .D(_14278_),
    .Q(_00345_),
    .CLK(clknet_leaf_21__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mcause_csr.rd_data_o[2]$_DFFE_PN0P_  (.RESET_B(net8248),
    .D(_14270_),
    .Q(_00346_),
    .CLK(clknet_leaf_21__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mcause_csr.rd_data_o[3]$_DFFE_PN0P_  (.RESET_B(net8248),
    .D(_14263_),
    .Q(_00347_),
    .CLK(clknet_leaf_21__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mcause_csr.rd_data_o[4]$_DFFE_PN0P_  (.RESET_B(net8248),
    .D(_14257_),
    .Q(_00348_),
    .CLK(clknet_leaf_21__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mcause_csr.rd_data_o[5]$_DFFE_PN0P_  (.RESET_B(net8249),
    .D(_14249_),
    .Q(_00349_),
    .CLK(clknet_leaf_26__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mepc_csr.rd_data_o[0]$_DFFE_PN0P_  (.RESET_B(net8251),
    .D(_14245_),
    .Q(_00350_),
    .CLK(clknet_leaf_22__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mepc_csr.rd_data_o[10]$_DFFE_PN0P_  (.RESET_B(net8254),
    .D(_14243_),
    .Q(_00351_),
    .CLK(clknet_leaf_34__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mepc_csr.rd_data_o[11]$_DFFE_PN0P_  (.RESET_B(net8261),
    .D(_14237_),
    .Q(_00352_),
    .CLK(clknet_leaf_35__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mepc_csr.rd_data_o[12]$_DFFE_PN0P_  (.RESET_B(net8258),
    .D(_14233_),
    .Q(_00353_),
    .CLK(clknet_leaf_34__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mepc_csr.rd_data_o[13]$_DFFE_PN0P_  (.RESET_B(net8254),
    .D(_14229_),
    .Q(_00354_),
    .CLK(clknet_leaf_34__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mepc_csr.rd_data_o[14]$_DFFE_PN0P_  (.RESET_B(net8258),
    .D(_14224_),
    .Q(_00355_),
    .CLK(clknet_leaf_39__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mepc_csr.rd_data_o[15]$_DFFE_PN0P_  (.RESET_B(net8247),
    .D(_14220_),
    .Q(_00356_),
    .CLK(clknet_leaf_21__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mepc_csr.rd_data_o[16]$_DFFE_PN0P_  (.RESET_B(net8261),
    .D(_14216_),
    .Q(_00357_),
    .CLK(clknet_leaf_34__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mepc_csr.rd_data_o[17]$_DFFE_PN0P_  (.RESET_B(net8264),
    .D(_14212_),
    .Q(_00358_),
    .CLK(clknet_leaf_32__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mepc_csr.rd_data_o[18]$_DFFE_PN0P_  (.RESET_B(net8263),
    .D(_14208_),
    .Q(_00359_),
    .CLK(clknet_leaf_32__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mepc_csr.rd_data_o[19]$_DFFE_PN0P_  (.RESET_B(net8264),
    .D(_14202_),
    .Q(_00360_),
    .CLK(clknet_leaf_32__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mepc_csr.rd_data_o[1]$_DFFE_PN0P_  (.RESET_B(net8245),
    .D(_14197_),
    .Q(_00361_),
    .CLK(clknet_leaf_21__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mepc_csr.rd_data_o[20]$_DFFE_PN0P_  (.RESET_B(net8259),
    .D(_14187_),
    .Q(_00362_),
    .CLK(clknet_leaf_34__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mepc_csr.rd_data_o[21]$_DFFE_PN0P_  (.RESET_B(net8269),
    .D(_14182_),
    .Q(_00363_),
    .CLK(clknet_leaf_27__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mepc_csr.rd_data_o[22]$_DFFE_PN0P_  (.RESET_B(net8281),
    .D(_14178_),
    .Q(_00364_),
    .CLK(clknet_leaf_27__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mepc_csr.rd_data_o[23]$_DFFE_PN0P_  (.RESET_B(net8281),
    .D(_14174_),
    .Q(_00365_),
    .CLK(clknet_leaf_27__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mepc_csr.rd_data_o[24]$_DFFE_PN0P_  (.RESET_B(net8269),
    .D(_14170_),
    .Q(_00366_),
    .CLK(clknet_leaf_33__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mepc_csr.rd_data_o[25]$_DFFE_PN0P_  (.RESET_B(net8268),
    .D(_14165_),
    .Q(_00367_),
    .CLK(clknet_leaf_33__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mepc_csr.rd_data_o[26]$_DFFE_PN0P_  (.RESET_B(net8268),
    .D(_14160_),
    .Q(_00368_),
    .CLK(clknet_leaf_33__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mepc_csr.rd_data_o[27]$_DFFE_PN0P_  (.RESET_B(net8259),
    .D(_14156_),
    .Q(_00369_),
    .CLK(clknet_leaf_33__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mepc_csr.rd_data_o[28]$_DFFE_PN0P_  (.RESET_B(net8263),
    .D(_14152_),
    .Q(_00370_),
    .CLK(clknet_leaf_32__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mepc_csr.rd_data_o[29]$_DFFE_PN0P_  (.RESET_B(net8263),
    .D(_14146_),
    .Q(_00371_),
    .CLK(clknet_leaf_32__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mepc_csr.rd_data_o[2]$_DFFE_PN0P_  (.RESET_B(net8247),
    .D(_14142_),
    .Q(_00372_),
    .CLK(clknet_leaf_21__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mepc_csr.rd_data_o[30]$_DFFE_PN0P_  (.RESET_B(net8263),
    .D(_14133_),
    .Q(_00373_),
    .CLK(clknet_leaf_32__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mepc_csr.rd_data_o[31]$_DFFE_PN0P_  (.RESET_B(net8261),
    .D(_14128_),
    .Q(_00374_),
    .CLK(clknet_leaf_34__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mepc_csr.rd_data_o[3]$_DFFE_PN0P_  (.RESET_B(net8247),
    .D(_14123_),
    .Q(_00375_),
    .CLK(clknet_leaf_20__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mepc_csr.rd_data_o[4]$_DFFE_PN0P_  (.RESET_B(net8246),
    .D(_14111_),
    .Q(_00376_),
    .CLK(clknet_leaf_20__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mepc_csr.rd_data_o[5]$_DFFE_PN0P_  (.RESET_B(net8282),
    .D(_14099_),
    .Q(_00377_),
    .CLK(clknet_leaf_27__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mepc_csr.rd_data_o[6]$_DFFE_PN0P_  (.RESET_B(net8267),
    .D(_14095_),
    .Q(_00378_),
    .CLK(clknet_leaf_27__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mepc_csr.rd_data_o[7]$_DFFE_PN0P_  (.RESET_B(net8266),
    .D(_14090_),
    .Q(_00379_),
    .CLK(clknet_leaf_34__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mepc_csr.rd_data_o[8]$_DFFE_PN0P_  (.RESET_B(net8260),
    .D(_14084_),
    .Q(_00380_),
    .CLK(clknet_leaf_39__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mepc_csr.rd_data_o[9]$_DFFE_PN0P_  (.RESET_B(net8261),
    .D(_14080_),
    .Q(_00381_),
    .CLK(clknet_leaf_34__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mie_csr.rd_data_o[0]$_DFFE_PN0P_  (.RESET_B(net8269),
    .D(_14073_),
    .Q(_00382_),
    .CLK(clknet_leaf_28__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mie_csr.rd_data_o[10]$_DFFE_PN0P_  (.RESET_B(net8270),
    .D(_14070_),
    .Q(_00383_),
    .CLK(clknet_leaf_32__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mie_csr.rd_data_o[11]$_DFFE_PN0P_  (.RESET_B(net8270),
    .D(_14068_),
    .Q(_00384_),
    .CLK(clknet_leaf_32__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mie_csr.rd_data_o[12]$_DFFE_PN0P_  (.RESET_B(net8270),
    .D(_14066_),
    .Q(_00385_),
    .CLK(clknet_leaf_31__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mie_csr.rd_data_o[13]$_DFFE_PN0P_  (.RESET_B(net8270),
    .D(_14064_),
    .Q(_00386_),
    .CLK(clknet_leaf_31__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mie_csr.rd_data_o[14]$_DFFE_PN0P_  (.RESET_B(net8270),
    .D(_14061_),
    .Q(_00387_),
    .CLK(clknet_leaf_31__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mie_csr.rd_data_o[15]$_DFFE_PN0P_  (.RESET_B(net8270),
    .D(_14058_),
    .Q(_00388_),
    .CLK(clknet_leaf_31__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mie_csr.rd_data_o[16]$_DFFE_PN0P_  (.RESET_B(net8269),
    .D(_14056_),
    .Q(_00389_),
    .CLK(clknet_leaf_28__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mie_csr.rd_data_o[17]$_DFFE_PN0P_  (.RESET_B(net8280),
    .D(_14053_),
    .Q(_00390_),
    .CLK(clknet_leaf_27__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mie_csr.rd_data_o[1]$_DFFE_PN0P_  (.RESET_B(net8270),
    .D(_14051_),
    .Q(_00391_),
    .CLK(clknet_leaf_31__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mie_csr.rd_data_o[2]$_DFFE_PN0P_  (.RESET_B(net8270),
    .D(_14049_),
    .Q(_00392_),
    .CLK(clknet_leaf_31__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mie_csr.rd_data_o[3]$_DFFE_PN0P_  (.RESET_B(net8271),
    .D(_14047_),
    .Q(_00393_),
    .CLK(clknet_leaf_31__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mie_csr.rd_data_o[4]$_DFFE_PN0P_  (.RESET_B(net8273),
    .D(_14045_),
    .Q(_00394_),
    .CLK(clknet_leaf_30__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mie_csr.rd_data_o[5]$_DFFE_PN0P_  (.RESET_B(net8273),
    .D(_14043_),
    .Q(_00395_),
    .CLK(clknet_leaf_28__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mie_csr.rd_data_o[6]$_DFFE_PN0P_  (.RESET_B(net8275),
    .D(_14041_),
    .Q(_00396_),
    .CLK(clknet_leaf_28__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mie_csr.rd_data_o[7]$_DFFE_PN0P_  (.RESET_B(net8275),
    .D(_14039_),
    .Q(_00397_),
    .CLK(clknet_leaf_27__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mie_csr.rd_data_o[8]$_DFFE_PN0P_  (.RESET_B(net8271),
    .D(_14037_),
    .Q(_00398_),
    .CLK(clknet_leaf_31__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mie_csr.rd_data_o[9]$_DFFE_PN0P_  (.RESET_B(net8271),
    .D(_14035_),
    .Q(_00399_),
    .CLK(clknet_leaf_31__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mscratch_csr.rd_data_o[0]$_DFFE_PN0P_  (.RESET_B(net8174),
    .D(_14032_),
    .Q(_00400_),
    .CLK(clknet_leaf_22__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mscratch_csr.rd_data_o[10]$_DFFE_PN0P_  (.RESET_B(net8279),
    .D(_14029_),
    .Q(_00401_),
    .CLK(clknet_leaf_30__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mscratch_csr.rd_data_o[11]$_DFFE_PN0P_  (.RESET_B(net8274),
    .D(_14026_),
    .Q(_00402_),
    .CLK(clknet_leaf_29__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mscratch_csr.rd_data_o[12]$_DFFE_PN0P_  (.RESET_B(net8274),
    .D(_14024_),
    .Q(_00403_),
    .CLK(clknet_leaf_28__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mscratch_csr.rd_data_o[13]$_DFFE_PN0P_  (.RESET_B(net8271),
    .D(_14022_),
    .Q(_00404_),
    .CLK(clknet_leaf_31__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mscratch_csr.rd_data_o[14]$_DFFE_PN0P_  (.RESET_B(net8185),
    .D(_14020_),
    .Q(_00405_),
    .CLK(clknet_leaf_28__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mscratch_csr.rd_data_o[15]$_DFFE_PN0P_  (.RESET_B(net8174),
    .D(_14018_),
    .Q(_00406_),
    .CLK(clknet_leaf_22__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mscratch_csr.rd_data_o[16]$_DFFE_PN0P_  (.RESET_B(net8278),
    .D(_14016_),
    .Q(_00407_),
    .CLK(clknet_leaf_29__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mscratch_csr.rd_data_o[17]$_DFFE_PN0P_  (.RESET_B(net8276),
    .D(_14014_),
    .Q(_00408_),
    .CLK(clknet_leaf_30__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mscratch_csr.rd_data_o[18]$_DFFE_PN0P_  (.RESET_B(net8276),
    .D(_14011_),
    .Q(_00409_),
    .CLK(clknet_leaf_31__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mscratch_csr.rd_data_o[19]$_DFFE_PN0P_  (.RESET_B(net8277),
    .D(_14008_),
    .Q(_00410_),
    .CLK(clknet_leaf_30__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mscratch_csr.rd_data_o[1]$_DFFE_PN0P_  (.RESET_B(net8174),
    .D(_14006_),
    .Q(_00411_),
    .CLK(clknet_leaf_22__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mscratch_csr.rd_data_o[20]$_DFFE_PN0P_  (.RESET_B(net8278),
    .D(_14004_),
    .Q(_00412_),
    .CLK(clknet_leaf_29__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mscratch_csr.rd_data_o[21]$_DFFE_PN0P_  (.RESET_B(net8185),
    .D(_14002_),
    .Q(_00413_),
    .CLK(clknet_leaf_25__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mscratch_csr.rd_data_o[22]$_DFFE_PN0P_  (.RESET_B(net8183),
    .D(_14000_),
    .Q(_00414_),
    .CLK(clknet_leaf_25__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mscratch_csr.rd_data_o[23]$_DFFE_PN0P_  (.RESET_B(net8183),
    .D(_13998_),
    .Q(_00415_),
    .CLK(clknet_leaf_25__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mscratch_csr.rd_data_o[24]$_DFFE_PN0P_  (.RESET_B(net8183),
    .D(_13996_),
    .Q(_00416_),
    .CLK(clknet_leaf_25__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mscratch_csr.rd_data_o[25]$_DFFE_PN0P_  (.RESET_B(net8277),
    .D(_13993_),
    .Q(_00417_),
    .CLK(clknet_leaf_29__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mscratch_csr.rd_data_o[26]$_DFFE_PN0P_  (.RESET_B(net8277),
    .D(_13990_),
    .Q(_00418_),
    .CLK(clknet_leaf_29__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mscratch_csr.rd_data_o[27]$_DFFE_PN0P_  (.RESET_B(net8179),
    .D(_13988_),
    .Q(_00419_),
    .CLK(clknet_leaf_29__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mscratch_csr.rd_data_o[28]$_DFFE_PN0P_  (.RESET_B(net8276),
    .D(_13986_),
    .Q(_00420_),
    .CLK(clknet_leaf_30__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mscratch_csr.rd_data_o[29]$_DFFE_PN0P_  (.RESET_B(net8272),
    .D(_13984_),
    .Q(_00421_),
    .CLK(clknet_leaf_31__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mscratch_csr.rd_data_o[2]$_DFFE_PN0P_  (.RESET_B(net8178),
    .D(_13982_),
    .Q(_00422_),
    .CLK(clknet_leaf_26__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mscratch_csr.rd_data_o[30]$_DFFE_PN0P_  (.RESET_B(net8272),
    .D(_13980_),
    .Q(_00423_),
    .CLK(clknet_leaf_31__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mscratch_csr.rd_data_o[31]$_DFFE_PN0P_  (.RESET_B(net8271),
    .D(_13977_),
    .Q(_00424_),
    .CLK(clknet_leaf_31__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mscratch_csr.rd_data_o[3]$_DFFE_PN0P_  (.RESET_B(net8174),
    .D(_13974_),
    .Q(_00425_),
    .CLK(clknet_leaf_22__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mscratch_csr.rd_data_o[4]$_DFFE_PN0P_  (.RESET_B(net8174),
    .D(_13972_),
    .Q(_00426_),
    .CLK(clknet_leaf_22__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mscratch_csr.rd_data_o[5]$_DFFE_PN0P_  (.RESET_B(net8185),
    .D(_13970_),
    .Q(_00427_),
    .CLK(clknet_leaf_25__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mscratch_csr.rd_data_o[6]$_DFFE_PN0P_  (.RESET_B(net8177),
    .D(_13968_),
    .Q(_00428_),
    .CLK(clknet_leaf_25__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mscratch_csr.rd_data_o[7]$_DFFE_PN0P_  (.RESET_B(net8275),
    .D(_13966_),
    .Q(_00429_),
    .CLK(clknet_leaf_28__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mscratch_csr.rd_data_o[8]$_DFFE_PN0P_  (.RESET_B(net8185),
    .D(_13964_),
    .Q(_00430_),
    .CLK(clknet_leaf_28__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mscratch_csr.rd_data_o[9]$_DFFE_PN0P_  (.RESET_B(net8279),
    .D(_13962_),
    .Q(_00431_),
    .CLK(clknet_leaf_30__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mstack_cause_csr.rd_data_o[0]$_DFFE_PN0P_  (.RESET_B(net8249),
    .D(_13958_),
    .Q(_00432_),
    .CLK(clknet_leaf_26__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mstack_cause_csr.rd_data_o[1]$_DFFE_PN0P_  (.RESET_B(net8250),
    .D(_13957_),
    .Q(_00433_),
    .CLK(clknet_leaf_22__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mstack_cause_csr.rd_data_o[2]$_DFFE_PN0P_  (.RESET_B(net8249),
    .D(_13956_),
    .Q(_00434_),
    .CLK(clknet_leaf_26__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mstack_cause_csr.rd_data_o[3]$_DFFE_PN0P_  (.RESET_B(net8247),
    .D(_13954_),
    .Q(_00435_),
    .CLK(clknet_leaf_20__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mstack_cause_csr.rd_data_o[4]$_DFFE_PN0P_  (.RESET_B(net8248),
    .D(_13952_),
    .Q(_00436_),
    .CLK(clknet_leaf_21__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mstack_cause_csr.rd_data_o[5]$_DFFE_PN0P_  (.RESET_B(net8249),
    .D(_13950_),
    .Q(_00437_),
    .CLK(clknet_leaf_27__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mstack_csr.rd_data_o[0]$_DFFE_PN0P_  (.RESET_B(net8250),
    .D(_13949_),
    .Q(_00438_),
    .CLK(clknet_leaf_22__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mstack_csr.rd_data_o[1]$_DFFE_PN0P_  (.RESET_B(net8247),
    .D(_13948_),
    .Q(_00439_),
    .CLK(clknet_leaf_21__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mstack_csr.rd_data_o[2]$_DFFE_PN1P_  (.RESET_B(net8178),
    .D(_13947_),
    .Q(_00002_),
    .CLK(clknet_leaf_26__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mstack_epc_csr.rd_data_o[0]$_DFFE_PN0P_  (.RESET_B(net8251),
    .D(_13945_),
    .Q(_00440_),
    .CLK(clknet_leaf_22__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mstack_epc_csr.rd_data_o[10]$_DFFE_PN0P_  (.RESET_B(net8253),
    .D(_13944_),
    .Q(_00441_),
    .CLK(clknet_leaf_39__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mstack_epc_csr.rd_data_o[11]$_DFFE_PN0P_  (.RESET_B(net8254),
    .D(_13943_),
    .Q(_00442_),
    .CLK(clknet_leaf_35__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mstack_epc_csr.rd_data_o[12]$_DFFE_PN0P_  (.RESET_B(net8253),
    .D(_13942_),
    .Q(_00443_),
    .CLK(clknet_leaf_39__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mstack_epc_csr.rd_data_o[13]$_DFFE_PN0P_  (.RESET_B(net8256),
    .D(_13941_),
    .Q(_00444_),
    .CLK(clknet_leaf_39__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mstack_epc_csr.rd_data_o[14]$_DFFE_PN0P_  (.RESET_B(net8253),
    .D(_13940_),
    .Q(_00445_),
    .CLK(clknet_leaf_39__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mstack_epc_csr.rd_data_o[15]$_DFFE_PN0P_  (.RESET_B(net8260),
    .D(_13939_),
    .Q(_00446_),
    .CLK(clknet_leaf_40__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mstack_epc_csr.rd_data_o[16]$_DFFE_PN0P_  (.RESET_B(net8266),
    .D(_13938_),
    .Q(_00447_),
    .CLK(clknet_leaf_34__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mstack_epc_csr.rd_data_o[17]$_DFFE_PN0P_  (.RESET_B(net8264),
    .D(_13937_),
    .Q(_00448_),
    .CLK(clknet_leaf_32__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mstack_epc_csr.rd_data_o[18]$_DFFE_PN0P_  (.RESET_B(net8264),
    .D(_13936_),
    .Q(_00449_),
    .CLK(clknet_leaf_32__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mstack_epc_csr.rd_data_o[19]$_DFFE_PN0P_  (.RESET_B(net8264),
    .D(_13935_),
    .Q(_00450_),
    .CLK(clknet_leaf_32__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mstack_epc_csr.rd_data_o[1]$_DFFE_PN0P_  (.RESET_B(net8245),
    .D(_13933_),
    .Q(_00451_),
    .CLK(clknet_leaf_20__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mstack_epc_csr.rd_data_o[20]$_DFFE_PN0P_  (.RESET_B(net8267),
    .D(_13932_),
    .Q(_00452_),
    .CLK(clknet_leaf_27__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mstack_epc_csr.rd_data_o[21]$_DFFE_PN0P_  (.RESET_B(net8259),
    .D(_13931_),
    .Q(_00453_),
    .CLK(clknet_leaf_33__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mstack_epc_csr.rd_data_o[22]$_DFFE_PN0P_  (.RESET_B(net8267),
    .D(_13930_),
    .Q(_00454_),
    .CLK(clknet_leaf_27__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mstack_epc_csr.rd_data_o[23]$_DFFE_PN0P_  (.RESET_B(net8267),
    .D(_13929_),
    .Q(_00455_),
    .CLK(clknet_leaf_27__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mstack_epc_csr.rd_data_o[24]$_DFFE_PN0P_  (.RESET_B(net8259),
    .D(_13928_),
    .Q(_00456_),
    .CLK(clknet_leaf_33__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mstack_epc_csr.rd_data_o[25]$_DFFE_PN0P_  (.RESET_B(net8259),
    .D(_13927_),
    .Q(_00457_),
    .CLK(clknet_leaf_33__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mstack_epc_csr.rd_data_o[26]$_DFFE_PN0P_  (.RESET_B(net8264),
    .D(_13925_),
    .Q(_00458_),
    .CLK(clknet_leaf_33__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mstack_epc_csr.rd_data_o[27]$_DFFE_PN0P_  (.RESET_B(net8259),
    .D(_13924_),
    .Q(_00459_),
    .CLK(clknet_leaf_33__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mstack_epc_csr.rd_data_o[28]$_DFFE_PN0P_  (.RESET_B(net8262),
    .D(_13923_),
    .Q(_00460_),
    .CLK(clknet_leaf_35__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mstack_epc_csr.rd_data_o[29]$_DFFE_PN0P_  (.RESET_B(net8262),
    .D(_13922_),
    .Q(_00461_),
    .CLK(clknet_leaf_35__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mstack_epc_csr.rd_data_o[2]$_DFFE_PN0P_  (.RESET_B(net8247),
    .D(_13921_),
    .Q(_00462_),
    .CLK(clknet_leaf_21__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mstack_epc_csr.rd_data_o[30]$_DFFE_PN0P_  (.RESET_B(net8262),
    .D(_13919_),
    .Q(_00463_),
    .CLK(clknet_leaf_35__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mstack_epc_csr.rd_data_o[31]$_DFFE_PN0P_  (.RESET_B(net8256),
    .D(_13918_),
    .Q(_00464_),
    .CLK(clknet_leaf_34__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mstack_epc_csr.rd_data_o[3]$_DFFE_PN0P_  (.RESET_B(net8247),
    .D(_13917_),
    .Q(_00465_),
    .CLK(clknet_leaf_20__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mstack_epc_csr.rd_data_o[4]$_DFFE_PN0P_  (.RESET_B(net8246),
    .D(_13915_),
    .Q(_00466_),
    .CLK(clknet_leaf_20__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mstack_epc_csr.rd_data_o[5]$_DFFE_PN0P_  (.RESET_B(net8258),
    .D(_13913_),
    .Q(_00467_),
    .CLK(clknet_leaf_40__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mstack_epc_csr.rd_data_o[6]$_DFFE_PN0P_  (.RESET_B(net8260),
    .D(_13912_),
    .Q(_00468_),
    .CLK(clknet_leaf_40__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mstack_epc_csr.rd_data_o[7]$_DFFE_PN0P_  (.RESET_B(net8266),
    .D(_13911_),
    .Q(_00469_),
    .CLK(clknet_leaf_34__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mstack_epc_csr.rd_data_o[8]$_DFFE_PN0P_  (.RESET_B(net8253),
    .D(_13910_),
    .Q(_00470_),
    .CLK(clknet_leaf_39__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mstack_epc_csr.rd_data_o[9]$_DFFE_PN0P_  (.RESET_B(net8254),
    .D(_13909_),
    .Q(_00471_),
    .CLK(clknet_leaf_34__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mstatus_csr.rd_data_o[0]$_DFFE_PN0P_  (.RESET_B(net8177),
    .D(_13908_),
    .Q(\cs_registers_i.csr_mstatus_tw_o ),
    .CLK(clknet_leaf_25__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mstatus_csr.rd_data_o[1]$_DFFE_PN0P_  (.RESET_B(net8274),
    .D(_13905_),
    .Q(_00472_),
    .CLK(clknet_leaf_30__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mstatus_csr.rd_data_o[2]$_DFFE_PN0P_  (.RESET_B(net8250),
    .D(_13903_),
    .Q(_00473_),
    .CLK(clknet_leaf_26__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mstatus_csr.rd_data_o[3]$_DFFE_PN0P_  (.RESET_B(net8250),
    .D(_13900_),
    .Q(_00474_),
    .CLK(clknet_leaf_22__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mstatus_csr.rd_data_o[4]$_DFFE_PN1P_  (.RESET_B(net8178),
    .D(_13894_),
    .Q(_00003_),
    .CLK(clknet_leaf_26__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mstatus_csr.rd_data_o[5]$_DFFE_PN0P_  (.RESET_B(net8178),
    .D(_13884_),
    .Q(\cs_registers_i.csr_mstatus_mie_o ),
    .CLK(clknet_leaf_26__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mtval_csr.rd_data_o[0]$_DFFE_PN0P_  (.RESET_B(net8246),
    .D(_13878_),
    .Q(_00475_),
    .CLK(clknet_leaf_20__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mtval_csr.rd_data_o[10]$_DFFE_PN0P_  (.RESET_B(net8280),
    .D(_13867_),
    .Q(_00476_),
    .CLK(clknet_leaf_27__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mtval_csr.rd_data_o[11]$_DFFE_PN0P_  (.RESET_B(net8175),
    .D(_13859_),
    .Q(_00477_),
    .CLK(clknet_leaf_26__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mtval_csr.rd_data_o[12]$_DFFE_PN0P_  (.RESET_B(net8250),
    .D(_13850_),
    .Q(_00478_),
    .CLK(clknet_leaf_26__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mtval_csr.rd_data_o[13]$_DFFE_PN0P_  (.RESET_B(net8249),
    .D(_13841_),
    .Q(_00479_),
    .CLK(clknet_leaf_26__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mtval_csr.rd_data_o[14]$_DFFE_PN0P_  (.RESET_B(net8280),
    .D(_13828_),
    .Q(_00480_),
    .CLK(clknet_leaf_27__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mtval_csr.rd_data_o[15]$_DFFE_PN0P_  (.RESET_B(net8246),
    .D(_13819_),
    .Q(_00481_),
    .CLK(clknet_leaf_20__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mtval_csr.rd_data_o[16]$_DFFE_PN0P_  (.RESET_B(net8250),
    .D(_13811_),
    .Q(_00482_),
    .CLK(clknet_leaf_22__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mtval_csr.rd_data_o[17]$_DFFE_PN0P_  (.RESET_B(net8177),
    .D(_13802_),
    .Q(_00483_),
    .CLK(clknet_leaf_24__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mtval_csr.rd_data_o[18]$_DFFE_PN0P_  (.RESET_B(net8186),
    .D(_13795_),
    .Q(_00484_),
    .CLK(clknet_leaf_24__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mtval_csr.rd_data_o[19]$_DFFE_PN0P_  (.RESET_B(net8184),
    .D(_13789_),
    .Q(_00485_),
    .CLK(clknet_leaf_24__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mtval_csr.rd_data_o[1]$_DFFE_PN0P_  (.RESET_B(net8251),
    .D(_13782_),
    .Q(_00486_),
    .CLK(clknet_leaf_21__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mtval_csr.rd_data_o[20]$_DFFE_PN0P_  (.RESET_B(net8184),
    .D(_13772_),
    .Q(_00487_),
    .CLK(clknet_leaf_24__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mtval_csr.rd_data_o[21]$_DFFE_PN0P_  (.RESET_B(net8177),
    .D(_13765_),
    .Q(_00488_),
    .CLK(clknet_leaf_26__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mtval_csr.rd_data_o[22]$_DFFE_PN0P_  (.RESET_B(net8200),
    .D(_13758_),
    .Q(_00489_),
    .CLK(clknet_leaf_24__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mtval_csr.rd_data_o[23]$_DFFE_PN0P_  (.RESET_B(net8184),
    .D(_13752_),
    .Q(_00490_),
    .CLK(clknet_leaf_24__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mtval_csr.rd_data_o[24]$_DFFE_PN0P_  (.RESET_B(net8200),
    .D(_13746_),
    .Q(_00491_),
    .CLK(clknet_leaf_24__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mtval_csr.rd_data_o[25]$_DFFE_PN0P_  (.RESET_B(net8184),
    .D(_13738_),
    .Q(_00492_),
    .CLK(clknet_leaf_24__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mtval_csr.rd_data_o[26]$_DFFE_PN0P_  (.RESET_B(net8200),
    .D(_13732_),
    .Q(_00493_),
    .CLK(clknet_leaf_24__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mtval_csr.rd_data_o[27]$_DFFE_PN0P_  (.RESET_B(net8200),
    .D(_13726_),
    .Q(_00494_),
    .CLK(clknet_leaf_24__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mtval_csr.rd_data_o[28]$_DFFE_PN0P_  (.RESET_B(net8186),
    .D(_13719_),
    .Q(_00495_),
    .CLK(clknet_leaf_24__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mtval_csr.rd_data_o[29]$_DFFE_PN0P_  (.RESET_B(net8186),
    .D(_13712_),
    .Q(_00496_),
    .CLK(clknet_leaf_25__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mtval_csr.rd_data_o[2]$_DFFE_PN0P_  (.RESET_B(net8175),
    .D(_13706_),
    .Q(_00497_),
    .CLK(clknet_leaf_26__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mtval_csr.rd_data_o[30]$_DFFE_PN0P_  (.RESET_B(net8274),
    .D(_13694_),
    .Q(_00498_),
    .CLK(clknet_leaf_30__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mtval_csr.rd_data_o[31]$_DFFE_PN0P_  (.RESET_B(net8178),
    .D(_13688_),
    .Q(_00499_),
    .CLK(clknet_leaf_26__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mtval_csr.rd_data_o[3]$_DFFE_PN0P_  (.RESET_B(net8252),
    .D(_13659_),
    .Q(_00500_),
    .CLK(clknet_leaf_22__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mtval_csr.rd_data_o[4]$_DFFE_PN0P_  (.RESET_B(net8251),
    .D(_13648_),
    .Q(_00501_),
    .CLK(clknet_leaf_22__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mtval_csr.rd_data_o[5]$_DFFE_PN0P_  (.RESET_B(net8177),
    .D(_13637_),
    .Q(_00502_),
    .CLK(clknet_leaf_24__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mtval_csr.rd_data_o[6]$_DFFE_PN0P_  (.RESET_B(net8175),
    .D(_13625_),
    .Q(_00503_),
    .CLK(clknet_leaf_26__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mtval_csr.rd_data_o[7]$_DFFE_PN0P_  (.RESET_B(net8250),
    .D(_13613_),
    .Q(_00504_),
    .CLK(clknet_leaf_26__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mtval_csr.rd_data_o[8]$_DFFE_PN0P_  (.RESET_B(net8175),
    .D(_13602_),
    .Q(_00505_),
    .CLK(clknet_leaf_26__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mtval_csr.rd_data_o[9]$_DFFE_PN0P_  (.RESET_B(net8275),
    .D(_13594_),
    .Q(_00506_),
    .CLK(clknet_leaf_28__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mtvec_csr.rd_data_o[10]$_DFFE_PN0P_  (.RESET_B(net8254),
    .D(_13560_),
    .Q(_00507_),
    .CLK(clknet_leaf_34__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mtvec_csr.rd_data_o[11]$_DFFE_PN0P_  (.RESET_B(net8255),
    .D(_13554_),
    .Q(_00508_),
    .CLK(clknet_leaf_35__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mtvec_csr.rd_data_o[12]$_DFFE_PN0P_  (.RESET_B(net8255),
    .D(_13548_),
    .Q(_00509_),
    .CLK(clknet_leaf_35__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mtvec_csr.rd_data_o[13]$_DFFE_PN0P_  (.RESET_B(net8255),
    .D(_13543_),
    .Q(_00510_),
    .CLK(clknet_leaf_35__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mtvec_csr.rd_data_o[14]$_DFFE_PN0P_  (.RESET_B(net8254),
    .D(_13538_),
    .Q(_00511_),
    .CLK(clknet_leaf_34__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mtvec_csr.rd_data_o[15]$_DFFE_PN0P_  (.RESET_B(net8260),
    .D(_13533_),
    .Q(_00512_),
    .CLK(clknet_leaf_40__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mtvec_csr.rd_data_o[16]$_DFFE_PN0P_  (.RESET_B(net8261),
    .D(_13528_),
    .Q(_00513_),
    .CLK(clknet_leaf_34__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mtvec_csr.rd_data_o[17]$_DFFE_PN0P_  (.RESET_B(net8262),
    .D(_13523_),
    .Q(_00514_),
    .CLK(clknet_leaf_35__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mtvec_csr.rd_data_o[18]$_DFFE_PN0P_  (.RESET_B(net8255),
    .D(_13517_),
    .Q(_00515_),
    .CLK(clknet_leaf_35__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mtvec_csr.rd_data_o[19]$_DFFE_PN0P_  (.RESET_B(net8265),
    .D(_13512_),
    .Q(_00516_),
    .CLK(clknet_leaf_35__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mtvec_csr.rd_data_o[20]$_DFFE_PN0P_  (.RESET_B(net8262),
    .D(_13507_),
    .Q(_00517_),
    .CLK(clknet_leaf_35__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mtvec_csr.rd_data_o[21]$_DFFE_PN0P_  (.RESET_B(net8265),
    .D(_13502_),
    .Q(_00518_),
    .CLK(clknet_leaf_35__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mtvec_csr.rd_data_o[22]$_DFFE_PN0P_  (.RESET_B(net8268),
    .D(_13496_),
    .Q(_00519_),
    .CLK(clknet_leaf_33__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mtvec_csr.rd_data_o[23]$_DFFE_PN0P_  (.RESET_B(net8269),
    .D(_13491_),
    .Q(_00520_),
    .CLK(clknet_leaf_33__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mtvec_csr.rd_data_o[24]$_DFFE_PN0P_  (.RESET_B(net8265),
    .D(_13485_),
    .Q(_00521_),
    .CLK(clknet_leaf_35__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mtvec_csr.rd_data_o[25]$_DFFE_PN0P_  (.RESET_B(net8262),
    .D(_13479_),
    .Q(_00522_),
    .CLK(clknet_leaf_35__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mtvec_csr.rd_data_o[26]$_DFFE_PN0P_  (.RESET_B(net8265),
    .D(_13472_),
    .Q(_00523_),
    .CLK(clknet_leaf_35__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mtvec_csr.rd_data_o[27]$_DFFE_PN0P_  (.RESET_B(net8265),
    .D(_13466_),
    .Q(_00524_),
    .CLK(clknet_leaf_35__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mtvec_csr.rd_data_o[28]$_DFFE_PN0P_  (.RESET_B(net8255),
    .D(_13460_),
    .Q(_00525_),
    .CLK(clknet_leaf_35__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mtvec_csr.rd_data_o[29]$_DFFE_PN0P_  (.RESET_B(net8255),
    .D(_13453_),
    .Q(_00526_),
    .CLK(clknet_leaf_36__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mtvec_csr.rd_data_o[30]$_DFFE_PN0P_  (.RESET_B(net8255),
    .D(_13447_),
    .Q(_00527_),
    .CLK(clknet_leaf_35__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mtvec_csr.rd_data_o[31]$_DFFE_PN0P_  (.RESET_B(net8255),
    .D(_13442_),
    .Q(_00528_),
    .CLK(clknet_leaf_36__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mtvec_csr.rd_data_o[8]$_DFFE_PN0P_  (.RESET_B(net8254),
    .D(_13437_),
    .Q(_00529_),
    .CLK(clknet_leaf_34__06563_));
 sg13g2_dfrbpq_1 \cs_registers_i.u_mtvec_csr.rd_data_o[9]$_DFFE_PN0P_  (.RESET_B(net8254),
    .D(_13432_),
    .Q(_00530_),
    .CLK(clknet_leaf_35__06563_));
 sg13g2_buf_16 delaybuf_0_core_clock (.X(delaynet_0_core_clock),
    .A(clk_i));
 sg13g2_buf_16 delaybuf_1_core_clock (.X(delaynet_1_core_clock),
    .A(delaynet_0_core_clock));
 sg13g2_buf_16 delaybuf_2_core_clock (.X(delaynet_2_core_clock),
    .A(delaynet_1_core_clock));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.div_by_zero_q$_DFFE_PN0P_  (.RESET_B(net8151),
    .D(_13416_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.div_by_zero_q ),
    .CLK(clknet_leaf_6__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0]$_DFFE_PN0P_  (.RESET_B(net8170),
    .D(_13413_),
    .Q(_00531_),
    .CLK(clknet_leaf_14__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[1]$_DFFE_PN0P_  (.RESET_B(net8170),
    .D(_13411_),
    .Q(_00532_),
    .CLK(clknet_leaf_15__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[2]$_DFFE_PN0P_  (.RESET_B(net8190),
    .D(_13404_),
    .Q(_00533_),
    .CLK(clknet_leaf_14__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[3]$_DFFE_PN0P_  (.RESET_B(net8170),
    .D(_13400_),
    .Q(_00534_),
    .CLK(clknet_leaf_14__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[4]$_DFFE_PN0P_  (.RESET_B(net8190),
    .D(_13398_),
    .Q(_00535_),
    .CLK(clknet_leaf_14__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[0]$_DFF_PN1_  (.RESET_B(net8161),
    .D(_13392_),
    .Q(_00004_),
    .CLK(clknet_leaf_7__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[1]$_DFF_PN0_  (.RESET_B(net8161),
    .D(_13389_),
    .Q(_00536_),
    .CLK(clknet_leaf_7__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[2]$_DFF_PN0_  (.RESET_B(net8161),
    .D(_13388_),
    .Q(_00537_),
    .CLK(clknet_leaf_7__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[3]$_DFF_PN0_  (.RESET_B(net8162),
    .D(_13385_),
    .Q(_00538_),
    .CLK(clknet_leaf_7__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[0]$_DFF_PN1_  (.RESET_B(net8151),
    .D(_13383_),
    .Q(_00005_),
    .CLK(clknet_leaf_6__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[1]$_DFF_PN0_  (.RESET_B(net8167),
    .D(_13381_),
    .Q(_00539_),
    .CLK(clknet_leaf_9__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[2]$_DFF_PN0_  (.RESET_B(net8167),
    .D(_13379_),
    .Q(_00540_),
    .CLK(clknet_leaf_6__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[3]$_DFF_PN0_  (.RESET_B(net8151),
    .D(_13378_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.div_valid ),
    .CLK(clknet_leaf_6__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[4]$_DFF_PN0_  (.RESET_B(net8151),
    .D(_13374_),
    .Q(_00541_),
    .CLK(clknet_leaf_6__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[5]$_DFF_PN0_  (.RESET_B(net8167),
    .D(_13372_),
    .Q(_00542_),
    .CLK(clknet_leaf_6__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[6]$_DFF_PN0_  (.RESET_B(net8171),
    .D(_13371_),
    .Q(_00543_),
    .CLK(clknet_leaf_10__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[0]$_DFFE_PN0P_  (.RESET_B(net8189),
    .D(_13368_),
    .Q(_00544_),
    .CLK(clknet_leaf_10__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[10]$_DFFE_PN0P_  (.RESET_B(net8166),
    .D(_13363_),
    .Q(_00545_),
    .CLK(clknet_leaf_19__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[11]$_DFFE_PN0P_  (.RESET_B(net8165),
    .D(_13359_),
    .Q(_00546_),
    .CLK(clknet_leaf_9__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[12]$_DFFE_PN0P_  (.RESET_B(net8189),
    .D(_13353_),
    .Q(_00547_),
    .CLK(clknet_leaf_9__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[13]$_DFFE_PN0P_  (.RESET_B(net8189),
    .D(_13348_),
    .Q(_00548_),
    .CLK(clknet_leaf_11__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[14]$_DFFE_PN0P_  (.RESET_B(net8189),
    .D(_13344_),
    .Q(_00549_),
    .CLK(clknet_leaf_11__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[15]$_DFFE_PN0P_  (.RESET_B(net8170),
    .D(_13340_),
    .Q(_00550_),
    .CLK(clknet_leaf_14__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[16]$_DFFE_PN0P_  (.RESET_B(net8166),
    .D(_13336_),
    .Q(_00551_),
    .CLK(clknet_leaf_6__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[17]$_DFFE_PN0P_  (.RESET_B(net8167),
    .D(_13332_),
    .Q(_00552_),
    .CLK(clknet_leaf_10__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[18]$_DFFE_PN0P_  (.RESET_B(net8166),
    .D(_13327_),
    .Q(_00553_),
    .CLK(clknet_leaf_19__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[19]$_DFFE_PN0P_  (.RESET_B(net8166),
    .D(_13322_),
    .Q(_00554_),
    .CLK(clknet_leaf_6__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[1]$_DFFE_PN0P_  (.RESET_B(net8164),
    .D(_13318_),
    .Q(_00555_),
    .CLK(clknet_leaf_9__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[20]$_DFFE_PN0P_  (.RESET_B(net8166),
    .D(_13314_),
    .Q(_00556_),
    .CLK(clknet_leaf_19__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[21]$_DFFE_PN0P_  (.RESET_B(net8166),
    .D(_13310_),
    .Q(_00557_),
    .CLK(clknet_leaf_19__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[22]$_DFFE_PN0P_  (.RESET_B(net8166),
    .D(_13306_),
    .Q(_00558_),
    .CLK(clknet_leaf_19__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[23]$_DFFE_PN0P_  (.RESET_B(net8169),
    .D(_13302_),
    .Q(_00559_),
    .CLK(clknet_leaf_14__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[24]$_DFFE_PN0P_  (.RESET_B(net8168),
    .D(_13298_),
    .Q(_00560_),
    .CLK(clknet_leaf_19__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[25]$_DFFE_PN0P_  (.RESET_B(net8168),
    .D(_13294_),
    .Q(_00561_),
    .CLK(clknet_leaf_19__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[26]$_DFFE_PN0P_  (.RESET_B(net8168),
    .D(_13289_),
    .Q(_00562_),
    .CLK(clknet_leaf_19__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[27]$_DFFE_PN0P_  (.RESET_B(net8170),
    .D(_13285_),
    .Q(_00563_),
    .CLK(clknet_leaf_19__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[28]$_DFFE_PN0P_  (.RESET_B(net8165),
    .D(_13281_),
    .Q(_00564_),
    .CLK(clknet_leaf_9__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[29]$_DFFE_PN0P_  (.RESET_B(net8167),
    .D(_13277_),
    .Q(_00565_),
    .CLK(clknet_leaf_10__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[2]$_DFFE_PN0P_  (.RESET_B(net8164),
    .D(_13273_),
    .Q(_00566_),
    .CLK(clknet_leaf_9__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[30]$_DFFE_PN0P_  (.RESET_B(net8165),
    .D(_13269_),
    .Q(_00567_),
    .CLK(clknet_leaf_10__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[31]$_DFFE_PN0P_  (.RESET_B(net8165),
    .D(_13265_),
    .Q(_00568_),
    .CLK(clknet_leaf_9__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[3]$_DFFE_PN0P_  (.RESET_B(net8169),
    .D(_13262_),
    .Q(_00569_),
    .CLK(clknet_leaf_14__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[4]$_DFFE_PN0P_  (.RESET_B(net8164),
    .D(_13258_),
    .Q(_00570_),
    .CLK(clknet_leaf_10__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[5]$_DFFE_PN0P_  (.RESET_B(net8171),
    .D(_13253_),
    .Q(_00571_),
    .CLK(clknet_leaf_14__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[6]$_DFFE_PN0P_  (.RESET_B(net8164),
    .D(_13248_),
    .Q(_00572_),
    .CLK(clknet_leaf_10__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[7]$_DFFE_PN0P_  (.RESET_B(net8170),
    .D(_13244_),
    .Q(_00573_),
    .CLK(clknet_leaf_14__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[8]$_DFFE_PN0P_  (.RESET_B(net8170),
    .D(_13240_),
    .Q(_00574_),
    .CLK(clknet_leaf_14__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[9]$_DFFE_PN0P_  (.RESET_B(net8166),
    .D(_13236_),
    .Q(_00575_),
    .CLK(clknet_leaf_6__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[0]$_DFFE_PN0P_  (.RESET_B(net8171),
    .D(_13232_),
    .Q(_00576_),
    .CLK(clknet_leaf_10__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[10]$_DFFE_PN0P_  (.RESET_B(net8193),
    .D(_13230_),
    .Q(_00577_),
    .CLK(clknet_leaf_14__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[11]$_DFFE_PN0P_  (.RESET_B(net8192),
    .D(_13228_),
    .Q(_00578_),
    .CLK(clknet_leaf_11__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[12]$_DFFE_PN0P_  (.RESET_B(net8190),
    .D(_13226_),
    .Q(_00579_),
    .CLK(clknet_leaf_11__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[13]$_DFFE_PN0P_  (.RESET_B(net8192),
    .D(_13224_),
    .Q(_00580_),
    .CLK(clknet_leaf_12__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[14]$_DFFE_PN0P_  (.RESET_B(net8192),
    .D(_13222_),
    .Q(_00581_),
    .CLK(clknet_leaf_12__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[15]$_DFFE_PN0P_  (.RESET_B(net8192),
    .D(_13220_),
    .Q(_00582_),
    .CLK(clknet_leaf_12__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[16]$_DFFE_PN0P_  (.RESET_B(net8171),
    .D(_13218_),
    .Q(_00583_),
    .CLK(clknet_leaf_10__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[17]$_DFFE_PN0P_  (.RESET_B(net8206),
    .D(_13216_),
    .Q(_00584_),
    .CLK(clknet_leaf_11__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[18]$_DFFE_PN0P_  (.RESET_B(net8191),
    .D(_13214_),
    .Q(_00585_),
    .CLK(clknet_leaf_11__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[19]$_DFFE_PN0P_  (.RESET_B(net8191),
    .D(_13212_),
    .Q(_00586_),
    .CLK(clknet_leaf_11__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[1]$_DFFE_PN0P_  (.RESET_B(net8164),
    .D(_13210_),
    .Q(_00587_),
    .CLK(clknet_leaf_10__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[20]$_DFFE_PN0P_  (.RESET_B(net8190),
    .D(_13208_),
    .Q(_00588_),
    .CLK(clknet_leaf_10__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[21]$_DFFE_PN0P_  (.RESET_B(net8191),
    .D(_13206_),
    .Q(_00589_),
    .CLK(clknet_leaf_11__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[22]$_DFFE_PN0P_  (.RESET_B(net8191),
    .D(_13204_),
    .Q(_00590_),
    .CLK(clknet_leaf_11__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[23]$_DFFE_PN0P_  (.RESET_B(net8191),
    .D(_13201_),
    .Q(_00591_),
    .CLK(clknet_leaf_11__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[24]$_DFFE_PN0P_  (.RESET_B(net8190),
    .D(_13199_),
    .Q(_00592_),
    .CLK(clknet_leaf_10__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[25]$_DFFE_PN0P_  (.RESET_B(net8191),
    .D(_13197_),
    .Q(_00593_),
    .CLK(clknet_leaf_11__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[26]$_DFFE_PN0P_  (.RESET_B(net8164),
    .D(_13195_),
    .Q(_00594_),
    .CLK(clknet_leaf_10__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[27]$_DFFE_PN0P_  (.RESET_B(net8164),
    .D(_13193_),
    .Q(_00595_),
    .CLK(clknet_leaf_11__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[28]$_DFFE_PN0P_  (.RESET_B(net8193),
    .D(_13191_),
    .Q(_00596_),
    .CLK(clknet_leaf_14__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[29]$_DFFE_PN0P_  (.RESET_B(net8191),
    .D(_13189_),
    .Q(_00597_),
    .CLK(clknet_leaf_11__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[2]$_DFFE_PN0P_  (.RESET_B(net8192),
    .D(_13186_),
    .Q(_00598_),
    .CLK(clknet_leaf_11__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[30]$_DFFE_PN0P_  (.RESET_B(net8164),
    .D(_13184_),
    .Q(_00599_),
    .CLK(clknet_leaf_10__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[31]$_DFFE_PN0P_  (.RESET_B(net8190),
    .D(_13182_),
    .Q(_00600_),
    .CLK(clknet_leaf_14__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[3]$_DFFE_PN0P_  (.RESET_B(net8192),
    .D(_13179_),
    .Q(_00601_),
    .CLK(clknet_leaf_11__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[4]$_DFFE_PN0P_  (.RESET_B(net8190),
    .D(_13176_),
    .Q(_00602_),
    .CLK(clknet_leaf_10__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[5]$_DFFE_PN0P_  (.RESET_B(net8205),
    .D(_13174_),
    .Q(_00603_),
    .CLK(clknet_leaf_11__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[6]$_DFFE_PN0P_  (.RESET_B(net8193),
    .D(_13172_),
    .Q(_00604_),
    .CLK(clknet_leaf_11__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[7]$_DFFE_PN0P_  (.RESET_B(net8193),
    .D(_13170_),
    .Q(_00605_),
    .CLK(clknet_leaf_11__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[8]$_DFFE_PN0P_  (.RESET_B(net8190),
    .D(_13167_),
    .Q(_00606_),
    .CLK(clknet_leaf_11__06563_));
 sg13g2_dfrbpq_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[9]$_DFFE_PN0P_  (.RESET_B(net8192),
    .D(_13165_),
    .Q(_00607_),
    .CLK(clknet_leaf_12__06563_));
 sg13g2_buf_1 fanout8287 (.A(net5859),
    .X(net8286));
 sg13g2_buf_1 fanout8288 (.A(net5859),
    .X(net8287));
 sg13g2_dfrbpq_1 \fetch_enable_q$_DFFE_PN0P_  (.RESET_B(net8242),
    .D(_13156_),
    .Q(fetch_enable_q),
    .CLK(clknet_leaf_38_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[1000]$_DFFE_PN0P_  (.RESET_B(net8091),
    .D(_13155_),
    .Q(_00608_),
    .CLK(clknet_leaf_9_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[1001]$_DFFE_PN0P_  (.RESET_B(net8027),
    .D(_13153_),
    .Q(_00609_),
    .CLK(clknet_leaf_14_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[1002]$_DFFE_PN0P_  (.RESET_B(net8056),
    .D(_13151_),
    .Q(_00610_),
    .CLK(clknet_leaf_2_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[1003]$_DFFE_PN0P_  (.RESET_B(net8024),
    .D(_13149_),
    .Q(_00611_),
    .CLK(clknet_leaf_14_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[1004]$_DFFE_PN0P_  (.RESET_B(net8098),
    .D(_13146_),
    .Q(_00612_),
    .CLK(clknet_leaf_17_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[1005]$_DFFE_PN0P_  (.RESET_B(net8096),
    .D(_13144_),
    .Q(_00613_),
    .CLK(clknet_leaf_24_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[1006]$_DFFE_PN0P_  (.RESET_B(net8067),
    .D(_13142_),
    .Q(_00614_),
    .CLK(clknet_leaf_9_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[1007]$_DFFE_PN0P_  (.RESET_B(net8155),
    .D(_13140_),
    .Q(_00615_),
    .CLK(clknet_leaf_33_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[1008]$_DFFE_PN0P_  (.RESET_B(net8053),
    .D(_13139_),
    .Q(_00616_),
    .CLK(clknet_leaf_4_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[1009]$_DFFE_PN0P_  (.RESET_B(net8038),
    .D(_13137_),
    .Q(_00617_),
    .CLK(clknet_leaf_1_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[100]$_DFFE_PN0P_  (.RESET_B(net8157),
    .D(_13135_),
    .Q(_00618_),
    .CLK(clknet_leaf_31_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[1010]$_DFFE_PN0P_  (.RESET_B(net8055),
    .D(_13133_),
    .Q(_00619_),
    .CLK(clknet_leaf_2_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[1011]$_DFFE_PN0P_  (.RESET_B(net8052),
    .D(_13131_),
    .Q(_00620_),
    .CLK(clknet_leaf_4_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[1012]$_DFFE_PN0P_  (.RESET_B(net8211),
    .D(_13129_),
    .Q(_00621_),
    .CLK(clknet_leaf_41_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[1013]$_DFFE_PN0P_  (.RESET_B(net8140),
    .D(_13127_),
    .Q(_00622_),
    .CLK(clknet_leaf_35_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[1014]$_DFFE_PN0P_  (.RESET_B(net8041),
    .D(_13124_),
    .Q(_00623_),
    .CLK(clknet_leaf_1_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[1015]$_DFFE_PN0P_  (.RESET_B(net8138),
    .D(_13122_),
    .Q(_00624_),
    .CLK(clknet_leaf_35_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[1016]$_DFFE_PN0P_  (.RESET_B(net8064),
    .D(_13119_),
    .Q(_00625_),
    .CLK(clknet_leaf_2_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[1017]$_DFFE_PN0P_  (.RESET_B(net8228),
    .D(_13117_),
    .Q(_00626_),
    .CLK(clknet_leaf_21_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[1018]$_DFFE_PN0P_  (.RESET_B(net8057),
    .D(_13114_),
    .Q(_00627_),
    .CLK(clknet_leaf_2_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[1019]$_DFFE_PN0P_  (.RESET_B(net8097),
    .D(_13111_),
    .Q(_00628_),
    .CLK(clknet_leaf_17_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[101]$_DFFE_PN0P_  (.RESET_B(net8141),
    .D(_13109_),
    .Q(_00629_),
    .CLK(clknet_leaf_22_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[1020]$_DFFE_PN0P_  (.RESET_B(net8110),
    .D(_13107_),
    .Q(_00630_),
    .CLK(clknet_leaf_26_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[1021]$_DFFE_PN0P_  (.RESET_B(net8038),
    .D(_13105_),
    .Q(_00631_),
    .CLK(clknet_leaf_3_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[1022]$_DFFE_PN0P_  (.RESET_B(net8132),
    .D(_13103_),
    .Q(_00632_),
    .CLK(clknet_leaf_22_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[1023]$_DFFE_PN0P_  (.RESET_B(net8157),
    .D(_13100_),
    .Q(_00633_),
    .CLK(clknet_leaf_31_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[102]$_DFFE_PN0P_  (.RESET_B(net8099),
    .D(_13098_),
    .Q(_00634_),
    .CLK(clknet_leaf_18_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[103]$_DFFE_PN0P_  (.RESET_B(net8115),
    .D(_13096_),
    .Q(_00635_),
    .CLK(clknet_leaf_30_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[104]$_DFFE_PN0P_  (.RESET_B(net8208),
    .D(_13094_),
    .Q(_00636_),
    .CLK(clknet_leaf_20_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[105]$_DFFE_PN0P_  (.RESET_B(net8208),
    .D(_13092_),
    .Q(_00637_),
    .CLK(clknet_leaf_19_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[106]$_DFFE_PN0P_  (.RESET_B(net8224),
    .D(_13090_),
    .Q(_00638_),
    .CLK(clknet_leaf_40_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[107]$_DFFE_PN0P_  (.RESET_B(net8083),
    .D(_13088_),
    .Q(_00639_),
    .CLK(clknet_leaf_19_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[108]$_DFFE_PN0P_  (.RESET_B(net8099),
    .D(_13086_),
    .Q(_00640_),
    .CLK(clknet_leaf_18_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[109]$_DFFE_PN0P_  (.RESET_B(net8156),
    .D(_13084_),
    .Q(_00641_),
    .CLK(clknet_leaf_23_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[110]$_DFFE_PN0P_  (.RESET_B(net8210),
    .D(_13082_),
    .Q(_00642_),
    .CLK(clknet_leaf_7_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[111]$_DFFE_PN0P_  (.RESET_B(net8137),
    .D(_13080_),
    .Q(_00643_),
    .CLK(clknet_leaf_37_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[112]$_DFFE_PN0P_  (.RESET_B(net8211),
    .D(_13079_),
    .Q(_00644_),
    .CLK(clknet_leaf_41_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[113]$_DFFE_PN0P_  (.RESET_B(net8220),
    .D(_13077_),
    .Q(_00645_),
    .CLK(clknet_leaf_41_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[114]$_DFFE_PN0P_  (.RESET_B(net8223),
    .D(_13074_),
    .Q(_00646_),
    .CLK(clknet_leaf_40_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[115]$_DFFE_PN0P_  (.RESET_B(net8214),
    .D(_13072_),
    .Q(_00647_),
    .CLK(clknet_leaf_42_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[116]$_DFFE_PN0P_  (.RESET_B(net8234),
    .D(_13070_),
    .Q(_00648_),
    .CLK(clknet_leaf_37_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[117]$_DFFE_PN0P_  (.RESET_B(net8139),
    .D(_13069_),
    .Q(_00649_),
    .CLK(clknet_leaf_36_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[118]$_DFFE_PN0P_  (.RESET_B(net8222),
    .D(_13066_),
    .Q(_00650_),
    .CLK(clknet_leaf_39_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[119]$_DFFE_PN0P_  (.RESET_B(net8134),
    .D(_13064_),
    .Q(_00651_),
    .CLK(clknet_leaf_36_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[120]$_DFFE_PN0P_  (.RESET_B(net8215),
    .D(_13061_),
    .Q(_00652_),
    .CLK(clknet_leaf_42_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[121]$_DFFE_PN0P_  (.RESET_B(net8132),
    .D(_13059_),
    .Q(_00653_),
    .CLK(clknet_leaf_34_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[122]$_DFFE_PN0P_  (.RESET_B(net8214),
    .D(_13056_),
    .Q(_00654_),
    .CLK(clknet_leaf_41_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[123]$_DFFE_PN0P_  (.RESET_B(net8126),
    .D(_13054_),
    .Q(_00655_),
    .CLK(clknet_leaf_23_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[124]$_DFFE_PN0P_  (.RESET_B(net8117),
    .D(_13051_),
    .Q(_00656_),
    .CLK(clknet_leaf_30_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[125]$_DFFE_PN0P_  (.RESET_B(net8221),
    .D(_13049_),
    .Q(_00657_),
    .CLK(clknet_leaf_40_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[126]$_DFFE_PN0P_  (.RESET_B(net8130),
    .D(_13046_),
    .Q(_00658_),
    .CLK(clknet_leaf_34_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[127]$_DFFE_PN0P_  (.RESET_B(net8148),
    .D(_13043_),
    .Q(_00659_),
    .CLK(clknet_leaf_33_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[128]$_DFFE_PN0P_  (.RESET_B(net8221),
    .D(_13041_),
    .Q(_00660_),
    .CLK(clknet_leaf_39_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[129]$_DFFE_PN0P_  (.RESET_B(net8209),
    .D(_13038_),
    .Q(_00661_),
    .CLK(clknet_leaf_7_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[130]$_DFFE_PN0P_  (.RESET_B(net8213),
    .D(_13036_),
    .Q(_00662_),
    .CLK(clknet_leaf_19_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[131]$_DFFE_PN0P_  (.RESET_B(net8087),
    .D(_13034_),
    .Q(_00663_),
    .CLK(clknet_leaf_7_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[132]$_DFFE_PN0P_  (.RESET_B(net8157),
    .D(_13032_),
    .Q(_00664_),
    .CLK(clknet_leaf_31_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[133]$_DFFE_PN0P_  (.RESET_B(net8143),
    .D(_13030_),
    .Q(_00665_),
    .CLK(clknet_leaf_30_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[134]$_DFFE_PN0P_  (.RESET_B(net8083),
    .D(_13028_),
    .Q(_00666_),
    .CLK(clknet_leaf_18_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[135]$_DFFE_PN0P_  (.RESET_B(net8115),
    .D(_13026_),
    .Q(_00667_),
    .CLK(clknet_leaf_31_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[136]$_DFFE_PN0P_  (.RESET_B(net8226),
    .D(_13024_),
    .Q(_00668_),
    .CLK(clknet_leaf_19_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[137]$_DFFE_PN0P_  (.RESET_B(net8226),
    .D(_13021_),
    .Q(_00669_),
    .CLK(clknet_leaf_19_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[138]$_DFFE_PN0P_  (.RESET_B(net8233),
    .D(_13019_),
    .Q(_00670_),
    .CLK(clknet_leaf_40_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[139]$_DFFE_PN0P_  (.RESET_B(net8084),
    .D(_13016_),
    .Q(_00671_),
    .CLK(clknet_leaf_19_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[140]$_DFFE_PN0P_  (.RESET_B(net8100),
    .D(_13014_),
    .Q(_00672_),
    .CLK(clknet_leaf_18_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[141]$_DFFE_PN0P_  (.RESET_B(net8143),
    .D(_13012_),
    .Q(_00673_),
    .CLK(clknet_leaf_27_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[142]$_DFFE_PN0P_  (.RESET_B(net8087),
    .D(_13009_),
    .Q(_00674_),
    .CLK(clknet_leaf_7_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[143]$_DFFE_PN0P_  (.RESET_B(net8135),
    .D(_13007_),
    .Q(_00675_),
    .CLK(clknet_leaf_37_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[144]$_DFFE_PN0P_  (.RESET_B(net8212),
    .D(_13006_),
    .Q(_00676_),
    .CLK(clknet_leaf_6_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[145]$_DFFE_PN0P_  (.RESET_B(net8218),
    .D(_13004_),
    .Q(_00677_),
    .CLK(clknet_leaf_39_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[146]$_DFFE_PN0P_  (.RESET_B(net8223),
    .D(_13002_),
    .Q(_00678_),
    .CLK(clknet_leaf_41_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[147]$_DFFE_PN0P_  (.RESET_B(net8220),
    .D(_13000_),
    .Q(_00679_),
    .CLK(clknet_leaf_41_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[148]$_DFFE_PN0P_  (.RESET_B(net8233),
    .D(_12998_),
    .Q(_00680_),
    .CLK(clknet_leaf_40_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[149]$_DFFE_PN0P_  (.RESET_B(net8229),
    .D(_12996_),
    .Q(_00681_),
    .CLK(clknet_leaf_36_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[150]$_DFFE_PN0P_  (.RESET_B(net8222),
    .D(_12993_),
    .Q(_00682_),
    .CLK(clknet_leaf_39_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[151]$_DFFE_PN0P_  (.RESET_B(net8135),
    .D(_12990_),
    .Q(_00683_),
    .CLK(clknet_leaf_36_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[152]$_DFFE_PN0P_  (.RESET_B(net8216),
    .D(_12986_),
    .Q(_00684_),
    .CLK(clknet_leaf_42_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[153]$_DFFE_PN0P_  (.RESET_B(net8227),
    .D(_12984_),
    .Q(_00685_),
    .CLK(clknet_leaf_35_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[154]$_DFFE_PN0P_  (.RESET_B(net8220),
    .D(_12981_),
    .Q(_00686_),
    .CLK(clknet_leaf_41_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[155]$_DFFE_PN0P_  (.RESET_B(net8128),
    .D(_12979_),
    .Q(_00687_),
    .CLK(clknet_leaf_23_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[156]$_DFFE_PN0P_  (.RESET_B(net8116),
    .D(_12977_),
    .Q(_00688_),
    .CLK(clknet_leaf_29_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[157]$_DFFE_PN0P_  (.RESET_B(net8221),
    .D(_12975_),
    .Q(_00689_),
    .CLK(clknet_leaf_39_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[158]$_DFFE_PN0P_  (.RESET_B(net8141),
    .D(_12973_),
    .Q(_00690_),
    .CLK(clknet_leaf_34_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[159]$_DFFE_PN0P_  (.RESET_B(net8148),
    .D(_12970_),
    .Q(_00691_),
    .CLK(clknet_leaf_34_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[160]$_DFFE_PN0P_  (.RESET_B(net8231),
    .D(_12965_),
    .Q(_00692_),
    .CLK(clknet_leaf_40_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[161]$_DFFE_PN0P_  (.RESET_B(net8209),
    .D(_12962_),
    .Q(_00693_),
    .CLK(clknet_leaf_7_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[162]$_DFFE_PN0P_  (.RESET_B(net8213),
    .D(_12960_),
    .Q(_00694_),
    .CLK(clknet_leaf_19_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[163]$_DFFE_PN0P_  (.RESET_B(net8087),
    .D(_12958_),
    .Q(_00695_),
    .CLK(clknet_leaf_7_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[164]$_DFFE_PN0P_  (.RESET_B(net8157),
    .D(_12956_),
    .Q(_00696_),
    .CLK(clknet_leaf_31_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[165]$_DFFE_PN0P_  (.RESET_B(net8143),
    .D(_12954_),
    .Q(_00697_),
    .CLK(clknet_leaf_30_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[166]$_DFFE_PN0P_  (.RESET_B(net8083),
    .D(_12951_),
    .Q(_00698_),
    .CLK(clknet_leaf_18_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[167]$_DFFE_PN0P_  (.RESET_B(net8115),
    .D(_12949_),
    .Q(_00699_),
    .CLK(clknet_leaf_31_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[168]$_DFFE_PN0P_  (.RESET_B(net8226),
    .D(_12947_),
    .Q(_00700_),
    .CLK(clknet_leaf_19_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[169]$_DFFE_PN0P_  (.RESET_B(net8208),
    .D(_12945_),
    .Q(_00701_),
    .CLK(clknet_leaf_19_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[170]$_DFFE_PN0P_  (.RESET_B(net8232),
    .D(_12943_),
    .Q(_00702_),
    .CLK(clknet_leaf_40_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[171]$_DFFE_PN0P_  (.RESET_B(net8084),
    .D(_12941_),
    .Q(_00703_),
    .CLK(clknet_leaf_19_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[172]$_DFFE_PN0P_  (.RESET_B(net8100),
    .D(_12939_),
    .Q(_00704_),
    .CLK(clknet_leaf_18_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[173]$_DFFE_PN0P_  (.RESET_B(net8156),
    .D(_12937_),
    .Q(_00705_),
    .CLK(clknet_leaf_23_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[174]$_DFFE_PN0P_  (.RESET_B(net8087),
    .D(_12935_),
    .Q(_00706_),
    .CLK(clknet_leaf_7_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[175]$_DFFE_PN0P_  (.RESET_B(net8137),
    .D(_12932_),
    .Q(_00707_),
    .CLK(clknet_leaf_37_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[176]$_DFFE_PN0P_  (.RESET_B(net8212),
    .D(_12931_),
    .Q(_00708_),
    .CLK(clknet_leaf_7_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[177]$_DFFE_PN0P_  (.RESET_B(net8218),
    .D(_12928_),
    .Q(_00709_),
    .CLK(clknet_leaf_39_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[178]$_DFFE_PN0P_  (.RESET_B(net8223),
    .D(_12926_),
    .Q(_00710_),
    .CLK(clknet_leaf_40_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[179]$_DFFE_PN0P_  (.RESET_B(net8220),
    .D(_12923_),
    .Q(_00711_),
    .CLK(clknet_leaf_42_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[180]$_DFFE_PN0P_  (.RESET_B(net8233),
    .D(_12921_),
    .Q(_00712_),
    .CLK(clknet_leaf_37_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[181]$_DFFE_PN0P_  (.RESET_B(net8229),
    .D(_12920_),
    .Q(_00713_),
    .CLK(clknet_leaf_36_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[182]$_DFFE_PN0P_  (.RESET_B(net8222),
    .D(_12917_),
    .Q(_00714_),
    .CLK(clknet_leaf_39_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[183]$_DFFE_PN0P_  (.RESET_B(net8135),
    .D(_12915_),
    .Q(_00715_),
    .CLK(clknet_leaf_36_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[184]$_DFFE_PN0P_  (.RESET_B(net8220),
    .D(_12912_),
    .Q(_00716_),
    .CLK(clknet_leaf_42_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[185]$_DFFE_PN0P_  (.RESET_B(net8227),
    .D(_12910_),
    .Q(_00717_),
    .CLK(clknet_leaf_21_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[186]$_DFFE_PN0P_  (.RESET_B(net8220),
    .D(_12906_),
    .Q(_00718_),
    .CLK(clknet_leaf_41_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[187]$_DFFE_PN0P_  (.RESET_B(net8128),
    .D(_12904_),
    .Q(_00719_),
    .CLK(clknet_leaf_23_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[188]$_DFFE_PN0P_  (.RESET_B(net8116),
    .D(_12901_),
    .Q(_00720_),
    .CLK(clknet_leaf_29_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[189]$_DFFE_PN0P_  (.RESET_B(net8221),
    .D(_12899_),
    .Q(_00721_),
    .CLK(clknet_leaf_39_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[190]$_DFFE_PN0P_  (.RESET_B(net8141),
    .D(_12897_),
    .Q(_00722_),
    .CLK(clknet_leaf_34_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[191]$_DFFE_PN0P_  (.RESET_B(net8148),
    .D(_12893_),
    .Q(_00723_),
    .CLK(clknet_leaf_34_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[192]$_DFFE_PN0P_  (.RESET_B(net8232),
    .D(_12889_),
    .Q(_00724_),
    .CLK(clknet_leaf_39_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[193]$_DFFE_PN0P_  (.RESET_B(net8211),
    .D(_12887_),
    .Q(_00725_),
    .CLK(clknet_leaf_7_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[194]$_DFFE_PN0P_  (.RESET_B(net8213),
    .D(_12885_),
    .Q(_00726_),
    .CLK(clknet_leaf_20_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[195]$_DFFE_PN0P_  (.RESET_B(net8088),
    .D(_12883_),
    .Q(_00727_),
    .CLK(clknet_leaf_7_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[196]$_DFFE_PN0P_  (.RESET_B(net8116),
    .D(_12881_),
    .Q(_00728_),
    .CLK(clknet_leaf_30_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[197]$_DFFE_PN0P_  (.RESET_B(net8143),
    .D(_12879_),
    .Q(_00729_),
    .CLK(clknet_leaf_30_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[198]$_DFFE_PN0P_  (.RESET_B(net8083),
    .D(_12877_),
    .Q(_00730_),
    .CLK(clknet_leaf_18_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[199]$_DFFE_PN0P_  (.RESET_B(net8115),
    .D(_12874_),
    .Q(_00731_),
    .CLK(clknet_leaf_30_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[200]$_DFFE_PN0P_  (.RESET_B(net8226),
    .D(_12871_),
    .Q(_00732_),
    .CLK(clknet_leaf_20_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[201]$_DFFE_PN0P_  (.RESET_B(net8083),
    .D(_12869_),
    .Q(_00733_),
    .CLK(clknet_leaf_19_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[202]$_DFFE_PN0P_  (.RESET_B(net8232),
    .D(_12866_),
    .Q(_00734_),
    .CLK(clknet_leaf_40_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[203]$_DFFE_PN0P_  (.RESET_B(net8101),
    .D(_12864_),
    .Q(_00735_),
    .CLK(clknet_leaf_16_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[204]$_DFFE_PN0P_  (.RESET_B(net8099),
    .D(_12862_),
    .Q(_00736_),
    .CLK(clknet_leaf_18_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[205]$_DFFE_PN0P_  (.RESET_B(net8156),
    .D(_12860_),
    .Q(_00737_),
    .CLK(clknet_leaf_23_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[206]$_DFFE_PN0P_  (.RESET_B(net8087),
    .D(_12858_),
    .Q(_00738_),
    .CLK(clknet_leaf_7_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[207]$_DFFE_PN0P_  (.RESET_B(net8135),
    .D(_12856_),
    .Q(_00739_),
    .CLK(clknet_leaf_37_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[208]$_DFFE_PN0P_  (.RESET_B(net8225),
    .D(_12855_),
    .Q(_00740_),
    .CLK(clknet_leaf_7_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[209]$_DFFE_PN0P_  (.RESET_B(net8218),
    .D(_12853_),
    .Q(_00741_),
    .CLK(clknet_leaf_39_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[210]$_DFFE_PN0P_  (.RESET_B(net8223),
    .D(_12850_),
    .Q(_00742_),
    .CLK(clknet_leaf_41_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[211]$_DFFE_PN0P_  (.RESET_B(net8215),
    .D(_12848_),
    .Q(_00743_),
    .CLK(clknet_leaf_42_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[212]$_DFFE_PN0P_  (.RESET_B(net8233),
    .D(_12845_),
    .Q(_00744_),
    .CLK(clknet_leaf_40_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[213]$_DFFE_PN0P_  (.RESET_B(net8229),
    .D(_12844_),
    .Q(_00745_),
    .CLK(clknet_leaf_36_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[214]$_DFFE_PN0P_  (.RESET_B(net8222),
    .D(_12841_),
    .Q(_00746_),
    .CLK(clknet_leaf_39_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[215]$_DFFE_PN0P_  (.RESET_B(net8135),
    .D(_12839_),
    .Q(_00747_),
    .CLK(clknet_leaf_37_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[216]$_DFFE_PN0P_  (.RESET_B(net8215),
    .D(_12836_),
    .Q(_00748_),
    .CLK(clknet_leaf_42_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[217]$_DFFE_PN0P_  (.RESET_B(net8227),
    .D(_12834_),
    .Q(_00749_),
    .CLK(clknet_leaf_21_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[218]$_DFFE_PN0P_  (.RESET_B(net8214),
    .D(_12831_),
    .Q(_00750_),
    .CLK(clknet_leaf_41_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[219]$_DFFE_PN0P_  (.RESET_B(net8126),
    .D(_12829_),
    .Q(_00751_),
    .CLK(clknet_leaf_23_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[220]$_DFFE_PN0P_  (.RESET_B(net8115),
    .D(_12827_),
    .Q(_00752_),
    .CLK(clknet_leaf_29_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[221]$_DFFE_PN0P_  (.RESET_B(net8221),
    .D(_12825_),
    .Q(_00753_),
    .CLK(clknet_leaf_39_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[222]$_DFFE_PN0P_  (.RESET_B(net8131),
    .D(_12823_),
    .Q(_00754_),
    .CLK(clknet_leaf_34_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[223]$_DFFE_PN0P_  (.RESET_B(net8148),
    .D(_12818_),
    .Q(_00755_),
    .CLK(clknet_leaf_34_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[224]$_DFFE_PN0P_  (.RESET_B(net8232),
    .D(_12814_),
    .Q(_00756_),
    .CLK(clknet_leaf_40_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[225]$_DFFE_PN0P_  (.RESET_B(net8210),
    .D(_12812_),
    .Q(_00757_),
    .CLK(clknet_leaf_20_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[226]$_DFFE_PN0P_  (.RESET_B(net8208),
    .D(_12810_),
    .Q(_00758_),
    .CLK(clknet_leaf_20_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[227]$_DFFE_PN0P_  (.RESET_B(net8210),
    .D(_12808_),
    .Q(_00759_),
    .CLK(clknet_leaf_7_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[228]$_DFFE_PN0P_  (.RESET_B(net8116),
    .D(_12806_),
    .Q(_00760_),
    .CLK(clknet_leaf_30_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[229]$_DFFE_PN0P_  (.RESET_B(net8141),
    .D(_12804_),
    .Q(_00761_),
    .CLK(clknet_leaf_23_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[230]$_DFFE_PN0P_  (.RESET_B(net8083),
    .D(_12802_),
    .Q(_00762_),
    .CLK(clknet_leaf_18_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[231]$_DFFE_PN0P_  (.RESET_B(net8115),
    .D(_12800_),
    .Q(_00763_),
    .CLK(clknet_leaf_30_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[232]$_DFFE_PN0P_  (.RESET_B(net8226),
    .D(_12798_),
    .Q(_00764_),
    .CLK(clknet_leaf_20_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[233]$_DFFE_PN0P_  (.RESET_B(net8285),
    .D(_12795_),
    .Q(_00765_),
    .CLK(clknet_leaf_19_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[234]$_DFFE_PN0P_  (.RESET_B(net8233),
    .D(_12793_),
    .Q(_00766_),
    .CLK(clknet_leaf_40_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[235]$_DFFE_PN0P_  (.RESET_B(net8101),
    .D(_12790_),
    .Q(_00767_),
    .CLK(clknet_leaf_18_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[236]$_DFFE_PN0P_  (.RESET_B(net8099),
    .D(_12787_),
    .Q(_00768_),
    .CLK(clknet_leaf_18_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[237]$_DFFE_PN0P_  (.RESET_B(net8142),
    .D(_12785_),
    .Q(_00769_),
    .CLK(clknet_leaf_23_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[238]$_DFFE_PN0P_  (.RESET_B(net8210),
    .D(_12783_),
    .Q(_00770_),
    .CLK(clknet_leaf_7_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[239]$_DFFE_PN0P_  (.RESET_B(net8136),
    .D(_12780_),
    .Q(_00771_),
    .CLK(clknet_leaf_37_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[240]$_DFFE_PN0P_  (.RESET_B(net8225),
    .D(_12779_),
    .Q(_00772_),
    .CLK(clknet_leaf_42_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[241]$_DFFE_PN0P_  (.RESET_B(net8218),
    .D(_12777_),
    .Q(_00773_),
    .CLK(clknet_leaf_39_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[242]$_DFFE_PN0P_  (.RESET_B(net8224),
    .D(_12775_),
    .Q(_00774_),
    .CLK(clknet_leaf_40_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[243]$_DFFE_PN0P_  (.RESET_B(net8215),
    .D(_12772_),
    .Q(_00775_),
    .CLK(clknet_leaf_42_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[244]$_DFFE_PN0P_  (.RESET_B(net8234),
    .D(_12770_),
    .Q(_00776_),
    .CLK(clknet_leaf_37_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[245]$_DFFE_PN0P_  (.RESET_B(net8139),
    .D(_12769_),
    .Q(_00777_),
    .CLK(clknet_leaf_36_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[246]$_DFFE_PN0P_  (.RESET_B(net8222),
    .D(_12766_),
    .Q(_00778_),
    .CLK(clknet_leaf_39_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[247]$_DFFE_PN0P_  (.RESET_B(net8137),
    .D(_12764_),
    .Q(_00779_),
    .CLK(clknet_leaf_37_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[248]$_DFFE_PN0P_  (.RESET_B(net8215),
    .D(_12761_),
    .Q(_00780_),
    .CLK(clknet_leaf_42_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[249]$_DFFE_PN0P_  (.RESET_B(net8132),
    .D(_12759_),
    .Q(_00781_),
    .CLK(clknet_leaf_34_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[250]$_DFFE_PN0P_  (.RESET_B(net8214),
    .D(_12756_),
    .Q(_00782_),
    .CLK(clknet_leaf_41_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[251]$_DFFE_PN0P_  (.RESET_B(net8126),
    .D(_12754_),
    .Q(_00783_),
    .CLK(clknet_leaf_23_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[252]$_DFFE_PN0P_  (.RESET_B(net8117),
    .D(_12752_),
    .Q(_00784_),
    .CLK(clknet_leaf_29_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[253]$_DFFE_PN0P_  (.RESET_B(net8221),
    .D(_12750_),
    .Q(_00785_),
    .CLK(clknet_leaf_38_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[254]$_DFFE_PN0P_  (.RESET_B(net8130),
    .D(_12748_),
    .Q(_00786_),
    .CLK(clknet_leaf_34_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[255]$_DFFE_PN0P_  (.RESET_B(net8147),
    .D(_12745_),
    .Q(_00787_),
    .CLK(clknet_leaf_33_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[256]$_DFFE_PN0P_  (.RESET_B(net8217),
    .D(_12741_),
    .Q(_00788_),
    .CLK(clknet_leaf_44_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[257]$_DFFE_PN0P_  (.RESET_B(net8088),
    .D(_12739_),
    .Q(_00789_),
    .CLK(clknet_leaf_8_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[258]$_DFFE_PN0P_  (.RESET_B(net8085),
    .D(_12737_),
    .Q(_00790_),
    .CLK(clknet_leaf_8_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[259]$_DFFE_PN0P_  (.RESET_B(net8065),
    .D(_12734_),
    .Q(_00791_),
    .CLK(clknet_leaf_6_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[260]$_DFFE_PN0P_  (.RESET_B(net8114),
    .D(_12732_),
    .Q(_00792_),
    .CLK(clknet_leaf_29_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[261]$_DFFE_PN0P_  (.RESET_B(net8111),
    .D(_12729_),
    .Q(_00793_),
    .CLK(clknet_leaf_27_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[262]$_DFFE_PN0P_  (.RESET_B(net8109),
    .D(_12727_),
    .Q(_00794_),
    .CLK(clknet_leaf_15_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[263]$_DFFE_PN0P_  (.RESET_B(net8114),
    .D(_12725_),
    .Q(_00795_),
    .CLK(clknet_leaf_29_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[264]$_DFFE_PN0P_  (.RESET_B(net8085),
    .D(_12723_),
    .Q(_00796_),
    .CLK(clknet_leaf_8_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[265]$_DFFE_PN0P_  (.RESET_B(net8093),
    .D(_12721_),
    .Q(_00797_),
    .CLK(clknet_leaf_15_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[266]$_DFFE_PN0P_  (.RESET_B(net8216),
    .D(_12719_),
    .Q(_00798_),
    .CLK(clknet_leaf_44_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[267]$_DFFE_PN0P_  (.RESET_B(net8095),
    .D(_12717_),
    .Q(_00799_),
    .CLK(clknet_leaf_15_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[268]$_DFFE_PN0P_  (.RESET_B(net8098),
    .D(_12715_),
    .Q(_00800_),
    .CLK(clknet_leaf_16_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[269]$_DFFE_PN0P_  (.RESET_B(net8123),
    .D(_12713_),
    .Q(_00801_),
    .CLK(clknet_leaf_24_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[270]$_DFFE_PN0P_  (.RESET_B(net8065),
    .D(_12711_),
    .Q(_00802_),
    .CLK(clknet_leaf_8_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[271]$_DFFE_PN0P_  (.RESET_B(net8235),
    .D(_12709_),
    .Q(_00803_),
    .CLK(clknet_leaf_37_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[272]$_DFFE_PN0P_  (.RESET_B(net8069),
    .D(_12708_),
    .Q(_00804_),
    .CLK(clknet_leaf_6_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[273]$_DFFE_PN0P_  (.RESET_B(net8062),
    .D(_12706_),
    .Q(_00805_),
    .CLK(clknet_leaf_46_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[274]$_DFFE_PN0P_  (.RESET_B(net8070),
    .D(_12704_),
    .Q(_00806_),
    .CLK(clknet_leaf_43_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[275]$_DFFE_PN0P_  (.RESET_B(net8068),
    .D(_12702_),
    .Q(_00807_),
    .CLK(clknet_leaf_5_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[276]$_DFFE_PN0P_  (.RESET_B(net8216),
    .D(_12700_),
    .Q(_00808_),
    .CLK(clknet_leaf_43_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[277]$_DFFE_PN0P_  (.RESET_B(net8139),
    .D(_12698_),
    .Q(_00809_),
    .CLK(clknet_leaf_35_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[278]$_DFFE_PN0P_  (.RESET_B(net8071),
    .D(_12695_),
    .Q(_00810_),
    .CLK(clknet_leaf_46_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[279]$_DFFE_PN0P_  (.RESET_B(net8129),
    .D(_12693_),
    .Q(_00811_),
    .CLK(clknet_leaf_34_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[280]$_DFFE_PN0P_  (.RESET_B(net8077),
    .D(_12690_),
    .Q(_00812_),
    .CLK(clknet_leaf_43_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[281]$_DFFE_PN0P_  (.RESET_B(net8127),
    .D(_12688_),
    .Q(_00813_),
    .CLK(clknet_leaf_21_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[282]$_DFFE_PN0P_  (.RESET_B(net8068),
    .D(_12685_),
    .Q(_00814_),
    .CLK(clknet_leaf_5_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[283]$_DFFE_PN0P_  (.RESET_B(net8125),
    .D(_12683_),
    .Q(_00815_),
    .CLK(clknet_leaf_17_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[284]$_DFFE_PN0P_  (.RESET_B(net8111),
    .D(_12681_),
    .Q(_00816_),
    .CLK(clknet_leaf_27_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[285]$_DFFE_PN0P_  (.RESET_B(net8071),
    .D(_12679_),
    .Q(_00817_),
    .CLK(clknet_leaf_43_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[286]$_DFFE_PN0P_  (.RESET_B(net8143),
    .D(_12677_),
    .Q(_00818_),
    .CLK(clknet_leaf_31_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[287]$_DFFE_PN0P_  (.RESET_B(net8163),
    .D(_12674_),
    .Q(_00819_),
    .CLK(clknet_leaf_31_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[288]$_DFFE_PN0P_  (.RESET_B(net8217),
    .D(_12670_),
    .Q(_00820_),
    .CLK(clknet_leaf_44_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[289]$_DFFE_PN0P_  (.RESET_B(net8088),
    .D(_12667_),
    .Q(_00821_),
    .CLK(clknet_leaf_8_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[290]$_DFFE_PN0P_  (.RESET_B(net8085),
    .D(_12665_),
    .Q(_00822_),
    .CLK(clknet_leaf_8_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[291]$_DFFE_PN0P_  (.RESET_B(net8066),
    .D(_12663_),
    .Q(_00823_),
    .CLK(clknet_leaf_7_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[292]$_DFFE_PN0P_  (.RESET_B(net8114),
    .D(_12661_),
    .Q(_00824_),
    .CLK(clknet_leaf_29_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[293]$_DFFE_PN0P_  (.RESET_B(net8111),
    .D(_12658_),
    .Q(_00825_),
    .CLK(clknet_leaf_27_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[294]$_DFFE_PN0P_  (.RESET_B(net8109),
    .D(_12656_),
    .Q(_00826_),
    .CLK(clknet_leaf_15_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[295]$_DFFE_PN0P_  (.RESET_B(net8114),
    .D(_12653_),
    .Q(_00827_),
    .CLK(clknet_leaf_29_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[296]$_DFFE_PN0P_  (.RESET_B(net8085),
    .D(_12651_),
    .Q(_00828_),
    .CLK(clknet_leaf_8_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[297]$_DFFE_PN0P_  (.RESET_B(net8093),
    .D(_12649_),
    .Q(_00829_),
    .CLK(clknet_leaf_15_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[298]$_DFFE_PN0P_  (.RESET_B(net8216),
    .D(_12647_),
    .Q(_00830_),
    .CLK(clknet_leaf_44_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[299]$_DFFE_PN0P_  (.RESET_B(net8095),
    .D(_12645_),
    .Q(_00831_),
    .CLK(clknet_leaf_15_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[300]$_DFFE_PN0P_  (.RESET_B(net8098),
    .D(_12643_),
    .Q(_00832_),
    .CLK(clknet_leaf_16_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[301]$_DFFE_PN0P_  (.RESET_B(net8123),
    .D(_12641_),
    .Q(_00833_),
    .CLK(clknet_leaf_24_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[302]$_DFFE_PN0P_  (.RESET_B(net8066),
    .D(_12639_),
    .Q(_00834_),
    .CLK(clknet_leaf_7_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[303]$_DFFE_PN0P_  (.RESET_B(net8134),
    .D(_12637_),
    .Q(_00835_),
    .CLK(clknet_leaf_38_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[304]$_DFFE_PN0P_  (.RESET_B(net8069),
    .D(_12636_),
    .Q(_00836_),
    .CLK(clknet_leaf_6_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[305]$_DFFE_PN0P_  (.RESET_B(net8076),
    .D(_12633_),
    .Q(_00837_),
    .CLK(clknet_leaf_46_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[306]$_DFFE_PN0P_  (.RESET_B(net8070),
    .D(_12630_),
    .Q(_00838_),
    .CLK(clknet_leaf_43_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[307]$_DFFE_PN0P_  (.RESET_B(net8068),
    .D(_12628_),
    .Q(_00839_),
    .CLK(clknet_leaf_5_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[308]$_DFFE_PN0P_  (.RESET_B(net8216),
    .D(_12626_),
    .Q(_00840_),
    .CLK(clknet_leaf_42_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[309]$_DFFE_PN0P_  (.RESET_B(net8139),
    .D(_12625_),
    .Q(_00841_),
    .CLK(clknet_leaf_36_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[310]$_DFFE_PN0P_  (.RESET_B(net8071),
    .D(_12622_),
    .Q(_00842_),
    .CLK(clknet_leaf_43_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[311]$_DFFE_PN0P_  (.RESET_B(net8129),
    .D(_12620_),
    .Q(_00843_),
    .CLK(clknet_leaf_35_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[312]$_DFFE_PN0P_  (.RESET_B(net8077),
    .D(_12617_),
    .Q(_00844_),
    .CLK(clknet_leaf_43_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[313]$_DFFE_PN0P_  (.RESET_B(net8127),
    .D(_12615_),
    .Q(_00845_),
    .CLK(clknet_leaf_21_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[314]$_DFFE_PN0P_  (.RESET_B(net8068),
    .D(_12612_),
    .Q(_00846_),
    .CLK(clknet_leaf_6_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[315]$_DFFE_PN0P_  (.RESET_B(net437),
    .D(_12610_),
    .Q(_00847_),
    .CLK(clknet_leaf_24_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[316]$_DFFE_PN0P_  (.RESET_B(net8111),
    .D(_12608_),
    .Q(_00848_),
    .CLK(clknet_leaf_27_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[317]$_DFFE_PN0P_  (.RESET_B(net8071),
    .D(_12605_),
    .Q(_00849_),
    .CLK(clknet_leaf_43_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[318]$_DFFE_PN0P_  (.RESET_B(net8143),
    .D(_12602_),
    .Q(_00850_),
    .CLK(clknet_leaf_30_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[319]$_DFFE_PN0P_  (.RESET_B(net8163),
    .D(_12599_),
    .Q(_00851_),
    .CLK(clknet_leaf_31_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[320]$_DFFE_PN0P_  (.RESET_B(net8217),
    .D(_12595_),
    .Q(_00852_),
    .CLK(clknet_leaf_44_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[321]$_DFFE_PN0P_  (.RESET_B(net8088),
    .D(_12593_),
    .Q(_00853_),
    .CLK(clknet_leaf_8_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[322]$_DFFE_PN0P_  (.RESET_B(net8085),
    .D(_12591_),
    .Q(_00854_),
    .CLK(clknet_leaf_19_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[323]$_DFFE_PN0P_  (.RESET_B(net8065),
    .D(_12589_),
    .Q(_00855_),
    .CLK(clknet_leaf_6_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[324]$_DFFE_PN0P_  (.RESET_B(net8114),
    .D(_12587_),
    .Q(_00856_),
    .CLK(clknet_leaf_29_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[325]$_DFFE_PN0P_  (.RESET_B(net8111),
    .D(_12585_),
    .Q(_00857_),
    .CLK(clknet_leaf_26_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[326]$_DFFE_PN0P_  (.RESET_B(net8101),
    .D(_12583_),
    .Q(_00858_),
    .CLK(clknet_leaf_16_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[327]$_DFFE_PN0P_  (.RESET_B(net8114),
    .D(_12581_),
    .Q(_00859_),
    .CLK(clknet_leaf_29_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[328]$_DFFE_PN0P_  (.RESET_B(net8085),
    .D(_12578_),
    .Q(_00860_),
    .CLK(clknet_leaf_8_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[329]$_DFFE_PN0P_  (.RESET_B(net8093),
    .D(_12575_),
    .Q(_00861_),
    .CLK(clknet_leaf_15_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[32]$_DFFE_PN0P_  (.RESET_B(net8224),
    .D(_12573_),
    .Q(_00862_),
    .CLK(clknet_leaf_39_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[330]$_DFFE_PN0P_  (.RESET_B(net8216),
    .D(_12571_),
    .Q(_00863_),
    .CLK(clknet_leaf_43_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[331]$_DFFE_PN0P_  (.RESET_B(net8095),
    .D(_12569_),
    .Q(_00864_),
    .CLK(clknet_leaf_15_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[332]$_DFFE_PN0P_  (.RESET_B(net8098),
    .D(_12567_),
    .Q(_00865_),
    .CLK(clknet_leaf_16_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[333]$_DFFE_PN0P_  (.RESET_B(net8120),
    .D(_12565_),
    .Q(_00866_),
    .CLK(clknet_leaf_24_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[334]$_DFFE_PN0P_  (.RESET_B(net8069),
    .D(_12563_),
    .Q(_00867_),
    .CLK(clknet_leaf_6_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[335]$_DFFE_PN0P_  (.RESET_B(net8134),
    .D(_12561_),
    .Q(_00868_),
    .CLK(clknet_leaf_36_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[336]$_DFFE_PN0P_  (.RESET_B(net8069),
    .D(_12560_),
    .Q(_00869_),
    .CLK(clknet_leaf_6_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[337]$_DFFE_PN0P_  (.RESET_B(net8075),
    .D(_12557_),
    .Q(_00870_),
    .CLK(clknet_leaf_44_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[338]$_DFFE_PN0P_  (.RESET_B(net8070),
    .D(_12555_),
    .Q(_00871_),
    .CLK(clknet_leaf_43_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[339]$_DFFE_PN0P_  (.RESET_B(net8068),
    .D(_12552_),
    .Q(_00872_),
    .CLK(clknet_leaf_5_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[33]$_DFFE_PN0P_  (.RESET_B(net8209),
    .D(_12550_),
    .Q(_00873_),
    .CLK(clknet_leaf_20_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[340]$_DFFE_PN0P_  (.RESET_B(net8216),
    .D(_12548_),
    .Q(_00874_),
    .CLK(clknet_leaf_42_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[341]$_DFFE_PN0P_  (.RESET_B(net8139),
    .D(_12547_),
    .Q(_00875_),
    .CLK(clknet_leaf_36_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[342]$_DFFE_PN0P_  (.RESET_B(net8071),
    .D(_12544_),
    .Q(_00876_),
    .CLK(clknet_leaf_44_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[343]$_DFFE_PN0P_  (.RESET_B(net8129),
    .D(_12541_),
    .Q(_00877_),
    .CLK(clknet_leaf_33_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[344]$_DFFE_PN0P_  (.RESET_B(net8077),
    .D(_12538_),
    .Q(_00878_),
    .CLK(clknet_leaf_43_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[345]$_DFFE_PN0P_  (.RESET_B(net8127),
    .D(_12536_),
    .Q(_00879_),
    .CLK(clknet_leaf_21_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[346]$_DFFE_PN0P_  (.RESET_B(net8212),
    .D(_12532_),
    .Q(_00880_),
    .CLK(clknet_leaf_6_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[347]$_DFFE_PN0P_  (.RESET_B(net437),
    .D(_12530_),
    .Q(_00881_),
    .CLK(clknet_leaf_17_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[348]$_DFFE_PN0P_  (.RESET_B(net8113),
    .D(_12528_),
    .Q(_00882_),
    .CLK(clknet_leaf_27_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[349]$_DFFE_PN0P_  (.RESET_B(net8071),
    .D(_12526_),
    .Q(_00883_),
    .CLK(clknet_leaf_43_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[34]$_DFFE_PN0P_  (.RESET_B(net8237),
    .D(_12524_),
    .Q(_00884_),
    .CLK(clknet_leaf_20_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[350]$_DFFE_PN0P_  (.RESET_B(net8143),
    .D(_12522_),
    .Q(_00885_),
    .CLK(clknet_leaf_31_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[351]$_DFFE_PN0P_  (.RESET_B(net8163),
    .D(_12519_),
    .Q(_00886_),
    .CLK(clknet_leaf_31_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[352]$_DFFE_PN0P_  (.RESET_B(net8218),
    .D(_12515_),
    .Q(_00887_),
    .CLK(clknet_leaf_44_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[353]$_DFFE_PN0P_  (.RESET_B(net8088),
    .D(_12513_),
    .Q(_00888_),
    .CLK(clknet_leaf_8_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[354]$_DFFE_PN0P_  (.RESET_B(net8085),
    .D(_12511_),
    .Q(_00889_),
    .CLK(clknet_leaf_19_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[355]$_DFFE_PN0P_  (.RESET_B(net8069),
    .D(_12509_),
    .Q(_00890_),
    .CLK(clknet_leaf_6_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[356]$_DFFE_PN0P_  (.RESET_B(net8114),
    .D(_12507_),
    .Q(_00891_),
    .CLK(clknet_leaf_29_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[357]$_DFFE_PN0P_  (.RESET_B(net8111),
    .D(_12505_),
    .Q(_00892_),
    .CLK(clknet_leaf_27_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[358]$_DFFE_PN0P_  (.RESET_B(net8023),
    .D(_12503_),
    .Q(_00893_),
    .CLK(clknet_leaf_15_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[359]$_DFFE_PN0P_  (.RESET_B(net8114),
    .D(_12501_),
    .Q(_00894_),
    .CLK(clknet_leaf_29_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[35]$_DFFE_PN0P_  (.RESET_B(net8210),
    .D(_12499_),
    .Q(_00895_),
    .CLK(clknet_leaf_21_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[360]$_DFFE_PN0P_  (.RESET_B(net8085),
    .D(_12497_),
    .Q(_00896_),
    .CLK(clknet_leaf_8_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[361]$_DFFE_PN0P_  (.RESET_B(net8093),
    .D(_12495_),
    .Q(_00897_),
    .CLK(clknet_leaf_19_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[362]$_DFFE_PN0P_  (.RESET_B(net8216),
    .D(_12493_),
    .Q(_00898_),
    .CLK(clknet_leaf_43_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[363]$_DFFE_PN0P_  (.RESET_B(net8095),
    .D(_12491_),
    .Q(_00899_),
    .CLK(clknet_leaf_15_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[364]$_DFFE_PN0P_  (.RESET_B(net8098),
    .D(_12489_),
    .Q(_00900_),
    .CLK(clknet_leaf_16_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[365]$_DFFE_PN0P_  (.RESET_B(net8120),
    .D(_12487_),
    .Q(_00901_),
    .CLK(clknet_leaf_24_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[366]$_DFFE_PN0P_  (.RESET_B(net8069),
    .D(_12485_),
    .Q(_00902_),
    .CLK(clknet_leaf_6_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[367]$_DFFE_PN0P_  (.RESET_B(net8137),
    .D(_12483_),
    .Q(_00903_),
    .CLK(clknet_leaf_37_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[368]$_DFFE_PN0P_  (.RESET_B(net8069),
    .D(_12482_),
    .Q(_00904_),
    .CLK(clknet_leaf_6_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[369]$_DFFE_PN0P_  (.RESET_B(net8075),
    .D(_12480_),
    .Q(_00905_),
    .CLK(clknet_leaf_44_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[36]$_DFFE_PN0P_  (.RESET_B(net8157),
    .D(_12478_),
    .Q(_00906_),
    .CLK(clknet_leaf_31_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[370]$_DFFE_PN0P_  (.RESET_B(net8077),
    .D(_12476_),
    .Q(_00907_),
    .CLK(clknet_leaf_43_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[371]$_DFFE_PN0P_  (.RESET_B(net8068),
    .D(_12474_),
    .Q(_00908_),
    .CLK(clknet_leaf_6_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[372]$_DFFE_PN0P_  (.RESET_B(net8234),
    .D(_12472_),
    .Q(_00909_),
    .CLK(clknet_leaf_37_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[373]$_DFFE_PN0P_  (.RESET_B(net8139),
    .D(_12471_),
    .Q(_00910_),
    .CLK(clknet_leaf_35_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[374]$_DFFE_PN0P_  (.RESET_B(net8076),
    .D(_12468_),
    .Q(_00911_),
    .CLK(clknet_leaf_46_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[375]$_DFFE_PN0P_  (.RESET_B(net8129),
    .D(_12466_),
    .Q(_00912_),
    .CLK(clknet_leaf_35_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[376]$_DFFE_PN0P_  (.RESET_B(net8077),
    .D(_12462_),
    .Q(_00913_),
    .CLK(clknet_leaf_43_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[377]$_DFFE_PN0P_  (.RESET_B(net8130),
    .D(_12460_),
    .Q(_00914_),
    .CLK(clknet_leaf_34_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[378]$_DFFE_PN0P_  (.RESET_B(net8212),
    .D(_12457_),
    .Q(_00915_),
    .CLK(clknet_leaf_6_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[379]$_DFFE_PN0P_  (.RESET_B(net437),
    .D(_12455_),
    .Q(_00916_),
    .CLK(clknet_leaf_24_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[37]$_DFFE_PN0P_  (.RESET_B(net8143),
    .D(_12453_),
    .Q(_00917_),
    .CLK(clknet_leaf_27_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[380]$_DFFE_PN0P_  (.RESET_B(net8112),
    .D(_12451_),
    .Q(_00918_),
    .CLK(clknet_leaf_27_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[381]$_DFFE_PN0P_  (.RESET_B(net8071),
    .D(_12449_),
    .Q(_00919_),
    .CLK(clknet_leaf_43_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[382]$_DFFE_PN0P_  (.RESET_B(net8130),
    .D(_12447_),
    .Q(_00920_),
    .CLK(clknet_leaf_34_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[383]$_DFFE_PN0P_  (.RESET_B(net8163),
    .D(_12444_),
    .Q(_00921_),
    .CLK(clknet_leaf_31_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[384]$_DFFE_PN0P_  (.RESET_B(net8217),
    .D(_12439_),
    .Q(_00922_),
    .CLK(clknet_leaf_44_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[385]$_DFFE_PN0P_  (.RESET_B(net8087),
    .D(_12437_),
    .Q(_00923_),
    .CLK(clknet_leaf_7_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[386]$_DFFE_PN0P_  (.RESET_B(net8092),
    .D(_12435_),
    .Q(_00924_),
    .CLK(clknet_leaf_13_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[387]$_DFFE_PN0P_  (.RESET_B(net8067),
    .D(_12433_),
    .Q(_00925_),
    .CLK(clknet_leaf_8_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[388]$_DFFE_PN0P_  (.RESET_B(net8118),
    .D(_12431_),
    .Q(_00926_),
    .CLK(clknet_leaf_30_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[389]$_DFFE_PN0P_  (.RESET_B(net8111),
    .D(_12428_),
    .Q(_00927_),
    .CLK(clknet_leaf_27_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[38]$_DFFE_PN0P_  (.RESET_B(net8099),
    .D(_12426_),
    .Q(_00928_),
    .CLK(clknet_leaf_24_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[390]$_DFFE_PN0P_  (.RESET_B(net8101),
    .D(_12424_),
    .Q(_00929_),
    .CLK(clknet_leaf_16_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[391]$_DFFE_PN0P_  (.RESET_B(net8113),
    .D(_12422_),
    .Q(_00930_),
    .CLK(clknet_leaf_30_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[392]$_DFFE_PN0P_  (.RESET_B(net8091),
    .D(_12419_),
    .Q(_00931_),
    .CLK(clknet_leaf_9_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[393]$_DFFE_PN0P_  (.RESET_B(net8084),
    .D(_12417_),
    .Q(_00932_),
    .CLK(clknet_leaf_15_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[394]$_DFFE_PN0P_  (.RESET_B(net8219),
    .D(_12414_),
    .Q(_00933_),
    .CLK(clknet_leaf_44_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[395]$_DFFE_PN0P_  (.RESET_B(net8027),
    .D(_12412_),
    .Q(_00934_),
    .CLK(clknet_leaf_14_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[396]$_DFFE_PN0P_  (.RESET_B(net8101),
    .D(_12409_),
    .Q(_00935_),
    .CLK(clknet_leaf_16_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[397]$_DFFE_PN0P_  (.RESET_B(net8124),
    .D(_12407_),
    .Q(_00936_),
    .CLK(clknet_leaf_24_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[398]$_DFFE_PN0P_  (.RESET_B(net8066),
    .D(_12405_),
    .Q(_00937_),
    .CLK(clknet_leaf_4_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[399]$_DFFE_PN0P_  (.RESET_B(net8134),
    .D(_12403_),
    .Q(_00938_),
    .CLK(clknet_leaf_36_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[39]$_DFFE_PN0P_  (.RESET_B(net8115),
    .D(_12401_),
    .Q(_00939_),
    .CLK(clknet_leaf_31_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[400]$_DFFE_PN0P_  (.RESET_B(net8065),
    .D(_12399_),
    .Q(_00940_),
    .CLK(clknet_leaf_6_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[401]$_DFFE_PN0P_  (.RESET_B(net8075),
    .D(_12396_),
    .Q(_00941_),
    .CLK(clknet_leaf_46_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[402]$_DFFE_PN0P_  (.RESET_B(net8072),
    .D(_12394_),
    .Q(_00942_),
    .CLK(clknet_leaf_43_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[403]$_DFFE_PN0P_  (.RESET_B(net8078),
    .D(_12391_),
    .Q(_00943_),
    .CLK(clknet_leaf_5_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[404]$_DFFE_PN0P_  (.RESET_B(net8219),
    .D(_12389_),
    .Q(_00944_),
    .CLK(clknet_leaf_44_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[405]$_DFFE_PN0P_  (.RESET_B(net8236),
    .D(_12387_),
    .Q(_00945_),
    .CLK(clknet_leaf_35_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[406]$_DFFE_PN0P_  (.RESET_B(net8059),
    .D(_12383_),
    .Q(_00946_),
    .CLK(clknet_leaf_46_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[407]$_DFFE_PN0P_  (.RESET_B(net8138),
    .D(_12381_),
    .Q(_00947_),
    .CLK(clknet_leaf_35_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[408]$_DFFE_PN0P_  (.RESET_B(net8070),
    .D(_12378_),
    .Q(_00948_),
    .CLK(clknet_leaf_5_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[409]$_DFFE_PN0P_  (.RESET_B(net8227),
    .D(_12376_),
    .Q(_00949_),
    .CLK(clknet_leaf_21_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[40]$_DFFE_PN0P_  (.RESET_B(net8208),
    .D(_12373_),
    .Q(_00950_),
    .CLK(clknet_leaf_20_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[410]$_DFFE_PN0P_  (.RESET_B(net8077),
    .D(_12371_),
    .Q(_00951_),
    .CLK(clknet_leaf_43_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[411]$_DFFE_PN0P_  (.RESET_B(net8125),
    .D(_12369_),
    .Q(_00952_),
    .CLK(clknet_leaf_18_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[412]$_DFFE_PN0P_  (.RESET_B(net8112),
    .D(_12367_),
    .Q(_00953_),
    .CLK(clknet_leaf_27_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[413]$_DFFE_PN0P_  (.RESET_B(net8062),
    .D(_12365_),
    .Q(_00954_),
    .CLK(clknet_leaf_46_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[414]$_DFFE_PN0P_  (.RESET_B(net8131),
    .D(_12363_),
    .Q(_00955_),
    .CLK(clknet_leaf_22_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[415]$_DFFE_PN0P_  (.RESET_B(net8162),
    .D(_12360_),
    .Q(_00956_),
    .CLK(clknet_leaf_31_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[416]$_DFFE_PN0P_  (.RESET_B(net8217),
    .D(_12356_),
    .Q(_00957_),
    .CLK(clknet_leaf_44_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[417]$_DFFE_PN0P_  (.RESET_B(net8087),
    .D(_12354_),
    .Q(_00958_),
    .CLK(clknet_leaf_7_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[418]$_DFFE_PN0P_  (.RESET_B(net8086),
    .D(_12352_),
    .Q(_00959_),
    .CLK(clknet_leaf_9_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[419]$_DFFE_PN0P_  (.RESET_B(net8067),
    .D(_12350_),
    .Q(_00960_),
    .CLK(clknet_leaf_8_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[41]$_DFFE_PN0P_  (.RESET_B(net8086),
    .D(_12348_),
    .Q(_00961_),
    .CLK(clknet_leaf_19_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[420]$_DFFE_PN0P_  (.RESET_B(net8117),
    .D(_12346_),
    .Q(_00962_),
    .CLK(clknet_leaf_30_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[421]$_DFFE_PN0P_  (.RESET_B(net8112),
    .D(_12344_),
    .Q(_00963_),
    .CLK(clknet_leaf_30_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[422]$_DFFE_PN0P_  (.RESET_B(net8101),
    .D(_12342_),
    .Q(_00964_),
    .CLK(clknet_leaf_16_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[423]$_DFFE_PN0P_  (.RESET_B(net8113),
    .D(_12340_),
    .Q(_00965_),
    .CLK(clknet_leaf_30_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[424]$_DFFE_PN0P_  (.RESET_B(net8090),
    .D(_12338_),
    .Q(_00966_),
    .CLK(clknet_leaf_9_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[425]$_DFFE_PN0P_  (.RESET_B(net8084),
    .D(_12336_),
    .Q(_00967_),
    .CLK(clknet_leaf_15_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[426]$_DFFE_PN0P_  (.RESET_B(net8217),
    .D(_12334_),
    .Q(_00968_),
    .CLK(clknet_leaf_44_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[427]$_DFFE_PN0P_  (.RESET_B(net8094),
    .D(_12332_),
    .Q(_00969_),
    .CLK(clknet_leaf_15_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[428]$_DFFE_PN0P_  (.RESET_B(net8100),
    .D(_12329_),
    .Q(_00970_),
    .CLK(clknet_leaf_18_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[429]$_DFFE_PN0P_  (.RESET_B(net8124),
    .D(_12327_),
    .Q(_00971_),
    .CLK(clknet_leaf_24_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[42]$_DFFE_PN0P_  (.RESET_B(net8224),
    .D(_12325_),
    .Q(_00972_),
    .CLK(clknet_leaf_40_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[430]$_DFFE_PN0P_  (.RESET_B(net8066),
    .D(_12323_),
    .Q(_00973_),
    .CLK(clknet_leaf_10_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[431]$_DFFE_PN0P_  (.RESET_B(net8133),
    .D(_12321_),
    .Q(_00974_),
    .CLK(clknet_leaf_38_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[432]$_DFFE_PN0P_  (.RESET_B(net8065),
    .D(_12320_),
    .Q(_00975_),
    .CLK(clknet_leaf_6_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[433]$_DFFE_PN0P_  (.RESET_B(net8073),
    .D(_12318_),
    .Q(_00976_),
    .CLK(clknet_leaf_46_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[434]$_DFFE_PN0P_  (.RESET_B(net8072),
    .D(_12316_),
    .Q(_00977_),
    .CLK(clknet_leaf_43_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[435]$_DFFE_PN0P_  (.RESET_B(net8068),
    .D(_12314_),
    .Q(_00978_),
    .CLK(clknet_leaf_6_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[436]$_DFFE_PN0P_  (.RESET_B(net8218),
    .D(_12312_),
    .Q(_00979_),
    .CLK(clknet_leaf_44_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[437]$_DFFE_PN0P_  (.RESET_B(net8236),
    .D(_12311_),
    .Q(_00980_),
    .CLK(clknet_leaf_35_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[438]$_DFFE_PN0P_  (.RESET_B(net8059),
    .D(_12308_),
    .Q(_00981_),
    .CLK(clknet_leaf_46_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[439]$_DFFE_PN0P_  (.RESET_B(net8134),
    .D(_12306_),
    .Q(_00982_),
    .CLK(clknet_leaf_35_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[43]$_DFFE_PN0P_  (.RESET_B(net8083),
    .D(_12303_),
    .Q(_00983_),
    .CLK(clknet_leaf_19_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[440]$_DFFE_PN0P_  (.RESET_B(net8070),
    .D(_12301_),
    .Q(_00984_),
    .CLK(clknet_leaf_5_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[441]$_DFFE_PN0P_  (.RESET_B(net8236),
    .D(_12299_),
    .Q(_00985_),
    .CLK(clknet_leaf_35_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[442]$_DFFE_PN0P_  (.RESET_B(net8077),
    .D(_12296_),
    .Q(_00986_),
    .CLK(clknet_leaf_5_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[443]$_DFFE_PN0P_  (.RESET_B(net8125),
    .D(_12294_),
    .Q(_00987_),
    .CLK(clknet_leaf_18_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[444]$_DFFE_PN0P_  (.RESET_B(net8112),
    .D(_12292_),
    .Q(_00988_),
    .CLK(clknet_leaf_27_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[445]$_DFFE_PN0P_  (.RESET_B(net8061),
    .D(_12290_),
    .Q(_00989_),
    .CLK(clknet_leaf_46_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[446]$_DFFE_PN0P_  (.RESET_B(net8132),
    .D(_12288_),
    .Q(_00990_),
    .CLK(clknet_leaf_34_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[447]$_DFFE_PN0P_  (.RESET_B(net8162),
    .D(_12284_),
    .Q(_00991_),
    .CLK(clknet_leaf_31_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[448]$_DFFE_PN0P_  (.RESET_B(net8217),
    .D(_12281_),
    .Q(_00992_),
    .CLK(clknet_leaf_44_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[449]$_DFFE_PN0P_  (.RESET_B(net8088),
    .D(_12279_),
    .Q(_00993_),
    .CLK(clknet_leaf_7_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[44]$_DFFE_PN0P_  (.RESET_B(net8099),
    .D(_12277_),
    .Q(_00994_),
    .CLK(clknet_leaf_18_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[450]$_DFFE_PN0P_  (.RESET_B(net8086),
    .D(_12275_),
    .Q(_00995_),
    .CLK(clknet_leaf_19_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[451]$_DFFE_PN0P_  (.RESET_B(net8067),
    .D(_12273_),
    .Q(_00996_),
    .CLK(clknet_leaf_8_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[452]$_DFFE_PN0P_  (.RESET_B(net8113),
    .D(_12270_),
    .Q(_00997_),
    .CLK(clknet_leaf_29_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[453]$_DFFE_PN0P_  (.RESET_B(net8111),
    .D(_12268_),
    .Q(_00998_),
    .CLK(clknet_leaf_27_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[454]$_DFFE_PN0P_  (.RESET_B(net8100),
    .D(_12266_),
    .Q(_00999_),
    .CLK(clknet_leaf_16_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[455]$_DFFE_PN0P_  (.RESET_B(net8113),
    .D(_12264_),
    .Q(_01000_),
    .CLK(clknet_leaf_29_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[456]$_DFFE_PN0P_  (.RESET_B(net8090),
    .D(_12262_),
    .Q(_01001_),
    .CLK(clknet_leaf_9_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[457]$_DFFE_PN0P_  (.RESET_B(net8084),
    .D(_12260_),
    .Q(_01002_),
    .CLK(clknet_leaf_15_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[458]$_DFFE_PN0P_  (.RESET_B(net8219),
    .D(_12258_),
    .Q(_01003_),
    .CLK(clknet_leaf_44_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[459]$_DFFE_PN0P_  (.RESET_B(net8094),
    .D(_12255_),
    .Q(_01004_),
    .CLK(clknet_leaf_15_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[45]$_DFFE_PN0P_  (.RESET_B(net8142),
    .D(_12253_),
    .Q(_01005_),
    .CLK(clknet_leaf_23_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[460]$_DFFE_PN0P_  (.RESET_B(net8100),
    .D(_12251_),
    .Q(_01006_),
    .CLK(clknet_leaf_18_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[461]$_DFFE_PN0P_  (.RESET_B(net8124),
    .D(_12249_),
    .Q(_01007_),
    .CLK(clknet_leaf_24_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[462]$_DFFE_PN0P_  (.RESET_B(net8066),
    .D(_12247_),
    .Q(_01008_),
    .CLK(clknet_leaf_6_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[463]$_DFFE_PN0P_  (.RESET_B(net8133),
    .D(_12244_),
    .Q(_01009_),
    .CLK(clknet_leaf_38_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[464]$_DFFE_PN0P_  (.RESET_B(net8065),
    .D(_12242_),
    .Q(_01010_),
    .CLK(clknet_leaf_6_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[465]$_DFFE_PN0P_  (.RESET_B(net8075),
    .D(_12240_),
    .Q(_01011_),
    .CLK(clknet_leaf_46_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[466]$_DFFE_PN0P_  (.RESET_B(net8071),
    .D(_12237_),
    .Q(_01012_),
    .CLK(clknet_leaf_43_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[467]$_DFFE_PN0P_  (.RESET_B(net8078),
    .D(_12235_),
    .Q(_01013_),
    .CLK(clknet_leaf_5_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[468]$_DFFE_PN0P_  (.RESET_B(net8219),
    .D(_12233_),
    .Q(_01014_),
    .CLK(clknet_leaf_44_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[469]$_DFFE_PN0P_  (.RESET_B(net8236),
    .D(_12232_),
    .Q(_01015_),
    .CLK(clknet_leaf_35_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[46]$_DFFE_PN0P_  (.RESET_B(net8211),
    .D(_12229_),
    .Q(_01016_),
    .CLK(clknet_leaf_42_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[470]$_DFFE_PN0P_  (.RESET_B(net8059),
    .D(_12226_),
    .Q(_01017_),
    .CLK(clknet_leaf_46_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[471]$_DFFE_PN0P_  (.RESET_B(net8138),
    .D(_12222_),
    .Q(_01018_),
    .CLK(clknet_leaf_35_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[472]$_DFFE_PN0P_  (.RESET_B(net8070),
    .D(_12219_),
    .Q(_01019_),
    .CLK(clknet_leaf_5_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[473]$_DFFE_PN0P_  (.RESET_B(net8227),
    .D(_12217_),
    .Q(_01020_),
    .CLK(clknet_leaf_35_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[474]$_DFFE_PN0P_  (.RESET_B(net8077),
    .D(_12214_),
    .Q(_01021_),
    .CLK(clknet_leaf_43_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[475]$_DFFE_PN0P_  (.RESET_B(net8125),
    .D(_12212_),
    .Q(_01022_),
    .CLK(clknet_leaf_18_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[476]$_DFFE_PN0P_  (.RESET_B(net8112),
    .D(_12210_),
    .Q(_01023_),
    .CLK(clknet_leaf_27_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[477]$_DFFE_PN0P_  (.RESET_B(net8061),
    .D(_12208_),
    .Q(_01024_),
    .CLK(clknet_leaf_46_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[478]$_DFFE_PN0P_  (.RESET_B(net8131),
    .D(_12206_),
    .Q(_01025_),
    .CLK(clknet_leaf_22_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[479]$_DFFE_PN0P_  (.RESET_B(net8162),
    .D(_12203_),
    .Q(_01026_),
    .CLK(clknet_leaf_32_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[47]$_DFFE_PN0P_  (.RESET_B(net8135),
    .D(_12199_),
    .Q(_01027_),
    .CLK(clknet_leaf_37_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[480]$_DFFE_PN0P_  (.RESET_B(net8217),
    .D(_12198_),
    .Q(_01028_),
    .CLK(clknet_leaf_44_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[481]$_DFFE_PN0P_  (.RESET_B(net8088),
    .D(_12196_),
    .Q(_01029_),
    .CLK(clknet_leaf_8_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[482]$_DFFE_PN0P_  (.RESET_B(net8086),
    .D(_12194_),
    .Q(_01030_),
    .CLK(clknet_leaf_9_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[483]$_DFFE_PN0P_  (.RESET_B(net8067),
    .D(_12192_),
    .Q(_01031_),
    .CLK(clknet_leaf_8_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[484]$_DFFE_PN0P_  (.RESET_B(net8117),
    .D(_12189_),
    .Q(_01032_),
    .CLK(clknet_leaf_30_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[485]$_DFFE_PN0P_  (.RESET_B(net8112),
    .D(_12186_),
    .Q(_01033_),
    .CLK(clknet_leaf_30_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[486]$_DFFE_PN0P_  (.RESET_B(net8100),
    .D(_12184_),
    .Q(_01034_),
    .CLK(clknet_leaf_16_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[487]$_DFFE_PN0P_  (.RESET_B(net8113),
    .D(_12182_),
    .Q(_01035_),
    .CLK(clknet_leaf_29_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[488]$_DFFE_PN0P_  (.RESET_B(net8090),
    .D(_12179_),
    .Q(_01036_),
    .CLK(clknet_leaf_9_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[489]$_DFFE_PN0P_  (.RESET_B(net8086),
    .D(_12177_),
    .Q(_01037_),
    .CLK(clknet_leaf_15_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[48]$_DFFE_PN0P_  (.RESET_B(net8211),
    .D(_12175_),
    .Q(_01038_),
    .CLK(clknet_leaf_42_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[490]$_DFFE_PN0P_  (.RESET_B(net8219),
    .D(_12173_),
    .Q(_01039_),
    .CLK(clknet_leaf_44_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[491]$_DFFE_PN0P_  (.RESET_B(net8094),
    .D(_12171_),
    .Q(_01040_),
    .CLK(clknet_leaf_15_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[492]$_DFFE_PN0P_  (.RESET_B(net8100),
    .D(_12169_),
    .Q(_01041_),
    .CLK(clknet_leaf_18_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[493]$_DFFE_PN0P_  (.RESET_B(net8124),
    .D(_12167_),
    .Q(_01042_),
    .CLK(clknet_leaf_24_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[494]$_DFFE_PN0P_  (.RESET_B(net8066),
    .D(_12165_),
    .Q(_01043_),
    .CLK(clknet_leaf_10_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[495]$_DFFE_PN0P_  (.RESET_B(net8133),
    .D(_12163_),
    .Q(_01044_),
    .CLK(clknet_leaf_38_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[496]$_DFFE_PN0P_  (.RESET_B(net8065),
    .D(_12162_),
    .Q(_01045_),
    .CLK(clknet_leaf_6_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[497]$_DFFE_PN0P_  (.RESET_B(net8075),
    .D(_12160_),
    .Q(_01046_),
    .CLK(clknet_leaf_44_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[498]$_DFFE_PN0P_  (.RESET_B(net8070),
    .D(_12158_),
    .Q(_01047_),
    .CLK(clknet_leaf_43_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[499]$_DFFE_PN0P_  (.RESET_B(net8068),
    .D(_12156_),
    .Q(_01048_),
    .CLK(clknet_leaf_6_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[49]$_DFFE_PN0P_  (.RESET_B(net8220),
    .D(_12154_),
    .Q(_01049_),
    .CLK(clknet_leaf_44_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[500]$_DFFE_PN0P_  (.RESET_B(net8219),
    .D(_12152_),
    .Q(_01050_),
    .CLK(clknet_leaf_44_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[501]$_DFFE_PN0P_  (.RESET_B(net8236),
    .D(_12151_),
    .Q(_01051_),
    .CLK(clknet_leaf_35_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[502]$_DFFE_PN0P_  (.RESET_B(net8062),
    .D(_12148_),
    .Q(_01052_),
    .CLK(clknet_leaf_46_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[503]$_DFFE_PN0P_  (.RESET_B(net8134),
    .D(_12146_),
    .Q(_01053_),
    .CLK(clknet_leaf_36_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[504]$_DFFE_PN0P_  (.RESET_B(net8070),
    .D(_12143_),
    .Q(_01054_),
    .CLK(clknet_leaf_43_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[505]$_DFFE_PN0P_  (.RESET_B(net8227),
    .D(_12140_),
    .Q(_01055_),
    .CLK(clknet_leaf_35_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[506]$_DFFE_PN0P_  (.RESET_B(net8078),
    .D(_12136_),
    .Q(_01056_),
    .CLK(clknet_leaf_5_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[507]$_DFFE_PN0P_  (.RESET_B(net8125),
    .D(_12133_),
    .Q(_01057_),
    .CLK(clknet_leaf_18_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[508]$_DFFE_PN0P_  (.RESET_B(net8112),
    .D(_12130_),
    .Q(_01058_),
    .CLK(clknet_leaf_30_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[509]$_DFFE_PN0P_  (.RESET_B(net8061),
    .D(_12128_),
    .Q(_01059_),
    .CLK(clknet_leaf_46_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[50]$_DFFE_PN0P_  (.RESET_B(net8223),
    .D(_12126_),
    .Q(_01060_),
    .CLK(clknet_leaf_41_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[510]$_DFFE_PN0P_  (.RESET_B(net8141),
    .D(_12124_),
    .Q(_01061_),
    .CLK(clknet_leaf_22_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[511]$_DFFE_PN0P_  (.RESET_B(net8162),
    .D(_12121_),
    .Q(_01062_),
    .CLK(clknet_leaf_31_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[512]$_DFFE_PN0P_  (.RESET_B(net8074),
    .D(_12117_),
    .Q(_01063_),
    .CLK(clknet_leaf_45_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[513]$_DFFE_PN0P_  (.RESET_B(net8029),
    .D(_12115_),
    .Q(_01064_),
    .CLK(clknet_leaf_11_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[514]$_DFFE_PN0P_  (.RESET_B(net8090),
    .D(_12113_),
    .Q(_01065_),
    .CLK(clknet_leaf_9_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[515]$_DFFE_PN0P_  (.RESET_B(net8035),
    .D(_12111_),
    .Q(_01066_),
    .CLK(clknet_leaf_10_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[516]$_DFFE_PN0P_  (.RESET_B(net8105),
    .D(_12109_),
    .Q(_01067_),
    .CLK(clknet_leaf_28_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[517]$_DFFE_PN0P_  (.RESET_B(net8142),
    .D(_12107_),
    .Q(_01068_),
    .CLK(clknet_leaf_26_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[518]$_DFFE_PN0P_  (.RESET_B(net8028),
    .D(_12105_),
    .Q(_01069_),
    .CLK(clknet_leaf_14_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[519]$_DFFE_PN0P_  (.RESET_B(net8105),
    .D(_12103_),
    .Q(_01070_),
    .CLK(clknet_leaf_28_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[51]$_DFFE_PN0P_  (.RESET_B(net8214),
    .D(_12101_),
    .Q(_01071_),
    .CLK(clknet_leaf_41_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[520]$_DFFE_PN0P_  (.RESET_B(net8080),
    .D(_12099_),
    .Q(_01072_),
    .CLK(clknet_leaf_9_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[521]$_DFFE_PN0P_  (.RESET_B(net8028),
    .D(_12097_),
    .Q(_01073_),
    .CLK(clknet_leaf_12_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[522]$_DFFE_PN0P_  (.RESET_B(net8075),
    .D(_12095_),
    .Q(_01074_),
    .CLK(clknet_leaf_45_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[523]$_DFFE_PN0P_  (.RESET_B(net8024),
    .D(_12093_),
    .Q(_01075_),
    .CLK(clknet_leaf_14_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[524]$_DFFE_PN0P_  (.RESET_B(net8102),
    .D(_12091_),
    .Q(_01076_),
    .CLK(clknet_leaf_16_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[525]$_DFFE_PN0P_  (.RESET_B(net8103),
    .D(_12089_),
    .Q(_01077_),
    .CLK(clknet_leaf_24_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[526]$_DFFE_PN0P_  (.RESET_B(net8034),
    .D(_12087_),
    .Q(_01078_),
    .CLK(clknet_leaf_11_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[527]$_DFFE_PN0P_  (.RESET_B(net8149),
    .D(_12085_),
    .Q(_01079_),
    .CLK(clknet_leaf_32_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[528]$_DFFE_PN0P_  (.RESET_B(net8043),
    .D(_12084_),
    .Q(_01080_),
    .CLK(clknet_leaf_0_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[529]$_DFFE_PN0P_  (.RESET_B(net8045),
    .D(_12082_),
    .Q(_01081_),
    .CLK(clknet_leaf_48_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[52]$_DFFE_PN0P_  (.RESET_B(net8234),
    .D(_12080_),
    .Q(_01082_),
    .CLK(clknet_leaf_40_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[530]$_DFFE_PN0P_  (.RESET_B(net8047),
    .D(_12079_),
    .Q(_01083_),
    .CLK(clknet_leaf_47_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[531]$_DFFE_PN0P_  (.RESET_B(net8042),
    .D(_12077_),
    .Q(_01084_),
    .CLK(clknet_leaf_1_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[532]$_DFFE_PN0P_  (.RESET_B(net8073),
    .D(_12075_),
    .Q(_01085_),
    .CLK(clknet_leaf_45_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[533]$_DFFE_PN0P_  (.RESET_B(net8236),
    .D(_12073_),
    .Q(_01086_),
    .CLK(clknet_leaf_36_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[534]$_DFFE_PN0P_  (.RESET_B(net8060),
    .D(_12070_),
    .Q(_01087_),
    .CLK(clknet_leaf_45_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[535]$_DFFE_PN0P_  (.RESET_B(net8134),
    .D(_12068_),
    .Q(_01088_),
    .CLK(clknet_leaf_38_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[536]$_DFFE_PN0P_  (.RESET_B(net8044),
    .D(_12065_),
    .Q(_01089_),
    .CLK(clknet_leaf_48_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[537]$_DFFE_PN0P_  (.RESET_B(net8209),
    .D(_12063_),
    .Q(_01090_),
    .CLK(clknet_leaf_21_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[538]$_DFFE_PN0P_  (.RESET_B(net8058),
    .D(_12059_),
    .Q(_01091_),
    .CLK(clknet_leaf_47_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[539]$_DFFE_PN0P_  (.RESET_B(net8107),
    .D(_12057_),
    .Q(_01092_),
    .CLK(clknet_leaf_16_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[53]$_DFFE_PN0P_  (.RESET_B(net8139),
    .D(_12055_),
    .Q(_01093_),
    .CLK(clknet_leaf_36_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[540]$_DFFE_PN0P_  (.RESET_B(net8110),
    .D(_12052_),
    .Q(_01094_),
    .CLK(clknet_leaf_26_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[541]$_DFFE_PN0P_  (.RESET_B(net8074),
    .D(_12050_),
    .Q(_01095_),
    .CLK(clknet_leaf_45_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[542]$_DFFE_PN0P_  (.RESET_B(net8127),
    .D(_12048_),
    .Q(_01096_),
    .CLK(clknet_leaf_22_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[543]$_DFFE_PN0P_  (.RESET_B(net8147),
    .D(_12045_),
    .Q(_01097_),
    .CLK(clknet_leaf_33_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[544]$_DFFE_PN0P_  (.RESET_B(net8074),
    .D(_12041_),
    .Q(_01098_),
    .CLK(clknet_leaf_45_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[545]$_DFFE_PN0P_  (.RESET_B(net8029),
    .D(_12039_),
    .Q(_01099_),
    .CLK(clknet_leaf_11_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[546]$_DFFE_PN0P_  (.RESET_B(net8090),
    .D(_12037_),
    .Q(_01100_),
    .CLK(clknet_leaf_8_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[547]$_DFFE_PN0P_  (.RESET_B(net8035),
    .D(_12035_),
    .Q(_01101_),
    .CLK(clknet_leaf_10_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[548]$_DFFE_PN0P_  (.RESET_B(net8105),
    .D(_12033_),
    .Q(_01102_),
    .CLK(clknet_leaf_28_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[549]$_DFFE_PN0P_  (.RESET_B(net8142),
    .D(_12031_),
    .Q(_01103_),
    .CLK(clknet_leaf_23_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[54]$_DFFE_PN0P_  (.RESET_B(net8222),
    .D(_12029_),
    .Q(_01104_),
    .CLK(clknet_leaf_39_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[550]$_DFFE_PN0P_  (.RESET_B(net8028),
    .D(_12027_),
    .Q(_01105_),
    .CLK(clknet_leaf_14_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[551]$_DFFE_PN0P_  (.RESET_B(net8105),
    .D(_12025_),
    .Q(_01106_),
    .CLK(clknet_leaf_28_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[552]$_DFFE_PN0P_  (.RESET_B(net8080),
    .D(_12022_),
    .Q(_01107_),
    .CLK(clknet_leaf_11_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[553]$_DFFE_PN0P_  (.RESET_B(net8028),
    .D(_12020_),
    .Q(_01108_),
    .CLK(clknet_leaf_12_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[554]$_DFFE_PN0P_  (.RESET_B(net8073),
    .D(_12018_),
    .Q(_01109_),
    .CLK(clknet_leaf_45_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[555]$_DFFE_PN0P_  (.RESET_B(net8024),
    .D(_12016_),
    .Q(_01110_),
    .CLK(clknet_leaf_14_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[556]$_DFFE_PN0P_  (.RESET_B(net8102),
    .D(_12014_),
    .Q(_01111_),
    .CLK(clknet_leaf_16_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[557]$_DFFE_PN0P_  (.RESET_B(net8103),
    .D(_12012_),
    .Q(_01112_),
    .CLK(clknet_leaf_24_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[558]$_DFFE_PN0P_  (.RESET_B(net8035),
    .D(_12010_),
    .Q(_01113_),
    .CLK(clknet_leaf_11_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[559]$_DFFE_PN0P_  (.RESET_B(net8149),
    .D(_12008_),
    .Q(_01114_),
    .CLK(clknet_leaf_32_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[55]$_DFFE_PN0P_  (.RESET_B(net8137),
    .D(_12007_),
    .Q(_01115_),
    .CLK(clknet_leaf_37_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[560]$_DFFE_PN0P_  (.RESET_B(net8049),
    .D(_12004_),
    .Q(_01116_),
    .CLK(clknet_leaf_0_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[561]$_DFFE_PN0P_  (.RESET_B(net8046),
    .D(_12002_),
    .Q(_01117_),
    .CLK(clknet_leaf_47_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[562]$_DFFE_PN0P_  (.RESET_B(net8047),
    .D(_12000_),
    .Q(_01118_),
    .CLK(clknet_leaf_47_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[563]$_DFFE_PN0P_  (.RESET_B(net8042),
    .D(_11998_),
    .Q(_01119_),
    .CLK(clknet_leaf_1_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[564]$_DFFE_PN0P_  (.RESET_B(net8073),
    .D(_11996_),
    .Q(_01120_),
    .CLK(clknet_leaf_45_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[565]$_DFFE_PN0P_  (.RESET_B(net8229),
    .D(_11995_),
    .Q(_01121_),
    .CLK(clknet_leaf_36_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[566]$_DFFE_PN0P_  (.RESET_B(net8060),
    .D(_11992_),
    .Q(_01122_),
    .CLK(clknet_leaf_45_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[567]$_DFFE_PN0P_  (.RESET_B(net8129),
    .D(_11990_),
    .Q(_01123_),
    .CLK(clknet_leaf_33_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[568]$_DFFE_PN0P_  (.RESET_B(net8045),
    .D(_11987_),
    .Q(_01124_),
    .CLK(clknet_leaf_0_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[569]$_DFFE_PN0P_  (.RESET_B(net8209),
    .D(_11985_),
    .Q(_01125_),
    .CLK(clknet_leaf_7_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[56]$_DFFE_PN0P_  (.RESET_B(net8215),
    .D(_11982_),
    .Q(_01126_),
    .CLK(clknet_leaf_42_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[570]$_DFFE_PN0P_  (.RESET_B(net8058),
    .D(_11980_),
    .Q(_01127_),
    .CLK(clknet_leaf_47_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[571]$_DFFE_PN0P_  (.RESET_B(net8107),
    .D(_11978_),
    .Q(_01128_),
    .CLK(clknet_leaf_17_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[572]$_DFFE_PN0P_  (.RESET_B(net8118),
    .D(_11976_),
    .Q(_01129_),
    .CLK(clknet_leaf_26_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[573]$_DFFE_PN0P_  (.RESET_B(net8074),
    .D(_11973_),
    .Q(_01130_),
    .CLK(clknet_leaf_45_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[574]$_DFFE_PN0P_  (.RESET_B(net8127),
    .D(_11971_),
    .Q(_01131_),
    .CLK(clknet_leaf_22_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[575]$_DFFE_PN0P_  (.RESET_B(net8147),
    .D(_11968_),
    .Q(_01132_),
    .CLK(clknet_leaf_33_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[576]$_DFFE_PN0P_  (.RESET_B(net8074),
    .D(_11964_),
    .Q(_01133_),
    .CLK(clknet_leaf_45_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[577]$_DFFE_PN0P_  (.RESET_B(net8029),
    .D(_11962_),
    .Q(_01134_),
    .CLK(clknet_leaf_11_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[578]$_DFFE_PN0P_  (.RESET_B(net8089),
    .D(_11960_),
    .Q(_01135_),
    .CLK(clknet_leaf_8_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[579]$_DFFE_PN0P_  (.RESET_B(net8035),
    .D(_11958_),
    .Q(_01136_),
    .CLK(clknet_leaf_10_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[57]$_DFFE_PN0P_  (.RESET_B(net8228),
    .D(_11956_),
    .Q(_01137_),
    .CLK(clknet_leaf_21_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[580]$_DFFE_PN0P_  (.RESET_B(net8123),
    .D(_11953_),
    .Q(_01138_),
    .CLK(clknet_leaf_28_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[581]$_DFFE_PN0P_  (.RESET_B(net8142),
    .D(_11951_),
    .Q(_01139_),
    .CLK(clknet_leaf_26_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[582]$_DFFE_PN0P_  (.RESET_B(net8028),
    .D(_11949_),
    .Q(_01140_),
    .CLK(clknet_leaf_12_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[583]$_DFFE_PN0P_  (.RESET_B(net8105),
    .D(_11947_),
    .Q(_01141_),
    .CLK(clknet_leaf_28_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[584]$_DFFE_PN0P_  (.RESET_B(net8034),
    .D(_11945_),
    .Q(_01142_),
    .CLK(clknet_leaf_11_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[585]$_DFFE_PN0P_  (.RESET_B(net8033),
    .D(_11943_),
    .Q(_01143_),
    .CLK(clknet_leaf_12_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[586]$_DFFE_PN0P_  (.RESET_B(net8073),
    .D(_11941_),
    .Q(_01144_),
    .CLK(clknet_leaf_46_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[587]$_DFFE_PN0P_  (.RESET_B(net8024),
    .D(_11939_),
    .Q(_01145_),
    .CLK(clknet_leaf_14_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[588]$_DFFE_PN0P_  (.RESET_B(net8102),
    .D(_11937_),
    .Q(_01146_),
    .CLK(clknet_leaf_16_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[589]$_DFFE_PN0P_  (.RESET_B(net8106),
    .D(_11935_),
    .Q(_01147_),
    .CLK(clknet_leaf_25_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[58]$_DFFE_PN0P_  (.RESET_B(net8214),
    .D(_11933_),
    .Q(_01148_),
    .CLK(clknet_leaf_41_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[590]$_DFFE_PN0P_  (.RESET_B(net8034),
    .D(_11930_),
    .Q(_01149_),
    .CLK(clknet_leaf_11_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[591]$_DFFE_PN0P_  (.RESET_B(net8149),
    .D(_11928_),
    .Q(_01150_),
    .CLK(clknet_leaf_32_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[592]$_DFFE_PN0P_  (.RESET_B(net8043),
    .D(_11927_),
    .Q(_01151_),
    .CLK(clknet_leaf_0_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[593]$_DFFE_PN0P_  (.RESET_B(net8046),
    .D(_11925_),
    .Q(_01152_),
    .CLK(clknet_leaf_47_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[594]$_DFFE_PN0P_  (.RESET_B(net8047),
    .D(_11922_),
    .Q(_01153_),
    .CLK(clknet_leaf_47_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[595]$_DFFE_PN0P_  (.RESET_B(net8042),
    .D(_11919_),
    .Q(_01154_),
    .CLK(clknet_leaf_0_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[596]$_DFFE_PN0P_  (.RESET_B(net8073),
    .D(_11917_),
    .Q(_01155_),
    .CLK(clknet_leaf_45_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[597]$_DFFE_PN0P_  (.RESET_B(net8236),
    .D(_11916_),
    .Q(_01156_),
    .CLK(clknet_leaf_36_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[598]$_DFFE_PN0P_  (.RESET_B(net8060),
    .D(_11913_),
    .Q(_01157_),
    .CLK(clknet_leaf_45_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[599]$_DFFE_PN0P_  (.RESET_B(net8129),
    .D(_11911_),
    .Q(_01158_),
    .CLK(clknet_leaf_33_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[59]$_DFFE_PN0P_  (.RESET_B(net8126),
    .D(_11908_),
    .Q(_01159_),
    .CLK(clknet_leaf_23_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[600]$_DFFE_PN0P_  (.RESET_B(net8045),
    .D(_11906_),
    .Q(_01160_),
    .CLK(clknet_leaf_0_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[601]$_DFFE_PN0P_  (.RESET_B(net8209),
    .D(_11904_),
    .Q(_01161_),
    .CLK(clknet_leaf_20_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[602]$_DFFE_PN0P_  (.RESET_B(net8058),
    .D(_11901_),
    .Q(_01162_),
    .CLK(clknet_leaf_47_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[603]$_DFFE_PN0P_  (.RESET_B(net8107),
    .D(_11898_),
    .Q(_01163_),
    .CLK(clknet_leaf_16_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[604]$_DFFE_PN0P_  (.RESET_B(net8110),
    .D(_11895_),
    .Q(_01164_),
    .CLK(clknet_leaf_26_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[605]$_DFFE_PN0P_  (.RESET_B(net8074),
    .D(_11893_),
    .Q(_01165_),
    .CLK(clknet_leaf_45_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[606]$_DFFE_PN0P_  (.RESET_B(net8127),
    .D(_11891_),
    .Q(_01166_),
    .CLK(clknet_leaf_22_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[607]$_DFFE_PN0P_  (.RESET_B(net8147),
    .D(_11888_),
    .Q(_01167_),
    .CLK(clknet_leaf_33_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[608]$_DFFE_PN0P_  (.RESET_B(net8074),
    .D(_11884_),
    .Q(_01168_),
    .CLK(clknet_leaf_45_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[609]$_DFFE_PN0P_  (.RESET_B(net8031),
    .D(_11882_),
    .Q(_01169_),
    .CLK(clknet_leaf_11_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[60]$_DFFE_PN0P_  (.RESET_B(net8117),
    .D(_11880_),
    .Q(_01170_),
    .CLK(clknet_leaf_29_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[610]$_DFFE_PN0P_  (.RESET_B(net8090),
    .D(_11878_),
    .Q(_01171_),
    .CLK(clknet_leaf_9_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[611]$_DFFE_PN0P_  (.RESET_B(net8051),
    .D(_11876_),
    .Q(_01172_),
    .CLK(clknet_leaf_10_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[612]$_DFFE_PN0P_  (.RESET_B(net8123),
    .D(_11874_),
    .Q(_01173_),
    .CLK(clknet_leaf_28_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[613]$_DFFE_PN0P_  (.RESET_B(net8142),
    .D(_11872_),
    .Q(_01174_),
    .CLK(clknet_leaf_26_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[614]$_DFFE_PN0P_  (.RESET_B(net8028),
    .D(_11869_),
    .Q(_01175_),
    .CLK(clknet_leaf_12_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[615]$_DFFE_PN0P_  (.RESET_B(net8105),
    .D(_11867_),
    .Q(_01176_),
    .CLK(clknet_leaf_28_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[616]$_DFFE_PN0P_  (.RESET_B(net8080),
    .D(_11864_),
    .Q(_01177_),
    .CLK(clknet_leaf_10_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[617]$_DFFE_PN0P_  (.RESET_B(net8033),
    .D(_11862_),
    .Q(_01178_),
    .CLK(clknet_leaf_12_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[618]$_DFFE_PN0P_  (.RESET_B(net8073),
    .D(_11860_),
    .Q(_01179_),
    .CLK(clknet_leaf_45_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[619]$_DFFE_PN0P_  (.RESET_B(net8024),
    .D(_11858_),
    .Q(_01180_),
    .CLK(clknet_leaf_14_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[61]$_DFFE_PN0P_  (.RESET_B(net8221),
    .D(_11856_),
    .Q(_01181_),
    .CLK(clknet_leaf_39_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[620]$_DFFE_PN0P_  (.RESET_B(net8102),
    .D(_11854_),
    .Q(_01182_),
    .CLK(clknet_leaf_16_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[621]$_DFFE_PN0P_  (.RESET_B(net8103),
    .D(_11852_),
    .Q(_01183_),
    .CLK(clknet_leaf_25_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[622]$_DFFE_PN0P_  (.RESET_B(net8035),
    .D(_11850_),
    .Q(_01184_),
    .CLK(clknet_leaf_11_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[623]$_DFFE_PN0P_  (.RESET_B(net8149),
    .D(_11848_),
    .Q(_01185_),
    .CLK(clknet_leaf_32_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[624]$_DFFE_PN0P_  (.RESET_B(net8043),
    .D(_11846_),
    .Q(_01186_),
    .CLK(clknet_leaf_0_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[625]$_DFFE_PN0P_  (.RESET_B(net8046),
    .D(_11844_),
    .Q(_01187_),
    .CLK(clknet_leaf_47_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[626]$_DFFE_PN0P_  (.RESET_B(net8047),
    .D(_11841_),
    .Q(_01188_),
    .CLK(clknet_leaf_47_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[627]$_DFFE_PN0P_  (.RESET_B(net8042),
    .D(_11839_),
    .Q(_01189_),
    .CLK(clknet_leaf_1_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[628]$_DFFE_PN0P_  (.RESET_B(net8073),
    .D(_11837_),
    .Q(_01190_),
    .CLK(clknet_leaf_45_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[629]$_DFFE_PN0P_  (.RESET_B(net8229),
    .D(_11836_),
    .Q(_01191_),
    .CLK(clknet_leaf_36_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[62]$_DFFE_PN0P_  (.RESET_B(net8131),
    .D(_11833_),
    .Q(_01192_),
    .CLK(clknet_leaf_34_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[630]$_DFFE_PN0P_  (.RESET_B(net8060),
    .D(_11830_),
    .Q(_01193_),
    .CLK(clknet_leaf_45_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[631]$_DFFE_PN0P_  (.RESET_B(net8129),
    .D(_11828_),
    .Q(_01194_),
    .CLK(clknet_leaf_33_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[632]$_DFFE_PN0P_  (.RESET_B(net8045),
    .D(_11825_),
    .Q(_01195_),
    .CLK(clknet_leaf_48_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[633]$_DFFE_PN0P_  (.RESET_B(net8209),
    .D(_11823_),
    .Q(_01196_),
    .CLK(clknet_leaf_20_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[634]$_DFFE_PN0P_  (.RESET_B(net8058),
    .D(_11819_),
    .Q(_01197_),
    .CLK(clknet_leaf_47_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[635]$_DFFE_PN0P_  (.RESET_B(net8107),
    .D(_11817_),
    .Q(_01198_),
    .CLK(clknet_leaf_17_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[636]$_DFFE_PN0P_  (.RESET_B(net8110),
    .D(_11815_),
    .Q(_01199_),
    .CLK(clknet_leaf_26_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[637]$_DFFE_PN0P_  (.RESET_B(net8074),
    .D(_11812_),
    .Q(_01200_),
    .CLK(clknet_leaf_45_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[638]$_DFFE_PN0P_  (.RESET_B(net8127),
    .D(_11809_),
    .Q(_01201_),
    .CLK(clknet_leaf_22_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[639]$_DFFE_PN0P_  (.RESET_B(net8147),
    .D(_11806_),
    .Q(_01202_),
    .CLK(clknet_leaf_32_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[63]$_DFFE_PN0P_  (.RESET_B(net8148),
    .D(_11802_),
    .Q(_01203_),
    .CLK(clknet_leaf_34_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[640]$_DFFE_PN0P_  (.RESET_B(net8046),
    .D(_11797_),
    .Q(_01204_),
    .CLK(clknet_leaf_47_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[641]$_DFFE_PN0P_  (.RESET_B(net8029),
    .D(_11795_),
    .Q(_01205_),
    .CLK(clknet_leaf_11_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[642]$_DFFE_PN0P_  (.RESET_B(net8090),
    .D(_11793_),
    .Q(_01206_),
    .CLK(clknet_leaf_9_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[643]$_DFFE_PN0P_  (.RESET_B(net8040),
    .D(_11791_),
    .Q(_01207_),
    .CLK(clknet_leaf_10_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[644]$_DFFE_PN0P_  (.RESET_B(net8106),
    .D(_11789_),
    .Q(_01208_),
    .CLK(clknet_leaf_26_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[645]$_DFFE_PN0P_  (.RESET_B(net8207),
    .D(_11787_),
    .Q(_01209_),
    .CLK(clknet_leaf_24_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[646]$_DFFE_PN0P_  (.RESET_B(net8032),
    .D(_11784_),
    .Q(_01210_),
    .CLK(clknet_leaf_13_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[647]$_DFFE_PN0P_  (.RESET_B(net8106),
    .D(_11782_),
    .Q(_01211_),
    .CLK(clknet_leaf_25_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[648]$_DFFE_PN0P_  (.RESET_B(net8034),
    .D(_11779_),
    .Q(_01212_),
    .CLK(clknet_leaf_11_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[649]$_DFFE_PN0P_  (.RESET_B(net8032),
    .D(_11777_),
    .Q(_01213_),
    .CLK(clknet_leaf_12_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[64]$_DFFE_PN0P_  (.RESET_B(net8232),
    .D(_11775_),
    .Q(_01214_),
    .CLK(clknet_leaf_39_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[650]$_DFFE_PN0P_  (.RESET_B(net8061),
    .D(_11773_),
    .Q(_01215_),
    .CLK(clknet_leaf_46_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[651]$_DFFE_PN0P_  (.RESET_B(net8026),
    .D(_11771_),
    .Q(_01216_),
    .CLK(clknet_leaf_13_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[652]$_DFFE_PN0P_  (.RESET_B(net8108),
    .D(_11769_),
    .Q(_01217_),
    .CLK(clknet_leaf_16_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[653]$_DFFE_PN0P_  (.RESET_B(net8103),
    .D(_11767_),
    .Q(_01218_),
    .CLK(clknet_leaf_25_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[654]$_DFFE_PN0P_  (.RESET_B(net8034),
    .D(_11765_),
    .Q(_01219_),
    .CLK(clknet_leaf_11_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[655]$_DFFE_PN0P_  (.RESET_B(net8149),
    .D(_11763_),
    .Q(_01220_),
    .CLK(clknet_leaf_32_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[656]$_DFFE_PN0P_  (.RESET_B(net8043),
    .D(_11762_),
    .Q(_01221_),
    .CLK(clknet_leaf_0_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[657]$_DFFE_PN0P_  (.RESET_B(net8047),
    .D(_11760_),
    .Q(_01222_),
    .CLK(clknet_leaf_48_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[658]$_DFFE_PN0P_  (.RESET_B(net8048),
    .D(_11758_),
    .Q(_01223_),
    .CLK(clknet_leaf_48_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[659]$_DFFE_PN0P_  (.RESET_B(net8049),
    .D(_11755_),
    .Q(_01224_),
    .CLK(clknet_leaf_0_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[65]$_DFFE_PN0P_  (.RESET_B(net8209),
    .D(_11753_),
    .Q(_01225_),
    .CLK(clknet_leaf_21_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[660]$_DFFE_PN0P_  (.RESET_B(net8060),
    .D(_11750_),
    .Q(_01226_),
    .CLK(clknet_leaf_45_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[661]$_DFFE_PN0P_  (.RESET_B(net8235),
    .D(_11749_),
    .Q(_01227_),
    .CLK(clknet_leaf_36_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[662]$_DFFE_PN0P_  (.RESET_B(net8044),
    .D(_11746_),
    .Q(_01228_),
    .CLK(clknet_leaf_47_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[663]$_DFFE_PN0P_  (.RESET_B(net8150),
    .D(_11744_),
    .Q(_01229_),
    .CLK(clknet_leaf_33_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[664]$_DFFE_PN0P_  (.RESET_B(net8049),
    .D(_11741_),
    .Q(_01230_),
    .CLK(clknet_leaf_0_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[665]$_DFFE_PN0P_  (.RESET_B(net8213),
    .D(_11739_),
    .Q(_01231_),
    .CLK(clknet_leaf_20_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[666]$_DFFE_PN0P_  (.RESET_B(net8042),
    .D(_11736_),
    .Q(_01232_),
    .CLK(clknet_leaf_47_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[667]$_DFFE_PN0P_  (.RESET_B(net8102),
    .D(_11734_),
    .Q(_01233_),
    .CLK(clknet_leaf_16_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[668]$_DFFE_PN0P_  (.RESET_B(net8104),
    .D(_11732_),
    .Q(_01234_),
    .CLK(clknet_leaf_25_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[669]$_DFFE_PN0P_  (.RESET_B(net8044),
    .D(_11730_),
    .Q(_01235_),
    .CLK(clknet_leaf_48_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[66]$_DFFE_PN0P_  (.RESET_B(net8208),
    .D(_11727_),
    .Q(_01236_),
    .CLK(clknet_leaf_20_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[670]$_DFFE_PN0P_  (.RESET_B(net8127),
    .D(_11724_),
    .Q(_01237_),
    .CLK(clknet_leaf_22_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[671]$_DFFE_PN0P_  (.RESET_B(net8146),
    .D(_11721_),
    .Q(_01238_),
    .CLK(clknet_leaf_32_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[672]$_DFFE_PN0P_  (.RESET_B(net8046),
    .D(_11717_),
    .Q(_01239_),
    .CLK(clknet_leaf_47_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[673]$_DFFE_PN0P_  (.RESET_B(net8029),
    .D(_11715_),
    .Q(_01240_),
    .CLK(clknet_leaf_11_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[674]$_DFFE_PN0P_  (.RESET_B(net8090),
    .D(_11713_),
    .Q(_01241_),
    .CLK(clknet_leaf_9_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[675]$_DFFE_PN0P_  (.RESET_B(net8040),
    .D(_11711_),
    .Q(_01242_),
    .CLK(clknet_leaf_10_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[676]$_DFFE_PN0P_  (.RESET_B(net8106),
    .D(_11709_),
    .Q(_01243_),
    .CLK(clknet_leaf_25_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[677]$_DFFE_PN0P_  (.RESET_B(net8142),
    .D(_11707_),
    .Q(_01244_),
    .CLK(clknet_leaf_23_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[678]$_DFFE_PN0P_  (.RESET_B(net8032),
    .D(_11705_),
    .Q(_01245_),
    .CLK(clknet_leaf_13_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[679]$_DFFE_PN0P_  (.RESET_B(net8104),
    .D(_11703_),
    .Q(_01246_),
    .CLK(clknet_leaf_25_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[67]$_DFFE_PN0P_  (.RESET_B(net8210),
    .D(_11701_),
    .Q(_01247_),
    .CLK(clknet_leaf_21_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[680]$_DFFE_PN0P_  (.RESET_B(net8035),
    .D(_11699_),
    .Q(_01248_),
    .CLK(clknet_leaf_11_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[681]$_DFFE_PN0P_  (.RESET_B(net8031),
    .D(_11697_),
    .Q(_01249_),
    .CLK(clknet_leaf_13_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[682]$_DFFE_PN0P_  (.RESET_B(net8061),
    .D(_11695_),
    .Q(_01250_),
    .CLK(clknet_leaf_46_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[683]$_DFFE_PN0P_  (.RESET_B(net8025),
    .D(_11693_),
    .Q(_01251_),
    .CLK(clknet_leaf_13_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[684]$_DFFE_PN0P_  (.RESET_B(net8109),
    .D(_11691_),
    .Q(_01252_),
    .CLK(clknet_leaf_16_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[685]$_DFFE_PN0P_  (.RESET_B(net8104),
    .D(_11689_),
    .Q(_01253_),
    .CLK(clknet_leaf_25_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[686]$_DFFE_PN0P_  (.RESET_B(net8034),
    .D(_11687_),
    .Q(_01254_),
    .CLK(clknet_leaf_11_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[687]$_DFFE_PN0P_  (.RESET_B(net8149),
    .D(_11685_),
    .Q(_01255_),
    .CLK(clknet_leaf_32_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[688]$_DFFE_PN0P_  (.RESET_B(net8043),
    .D(_11683_),
    .Q(_01256_),
    .CLK(clknet_leaf_0_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[689]$_DFFE_PN0P_  (.RESET_B(net8045),
    .D(_11680_),
    .Q(_01257_),
    .CLK(clknet_leaf_48_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[68]$_DFFE_PN0P_  (.RESET_B(net8157),
    .D(_11677_),
    .Q(_01258_),
    .CLK(clknet_leaf_31_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[690]$_DFFE_PN0P_  (.RESET_B(net8048),
    .D(_11675_),
    .Q(_01259_),
    .CLK(clknet_leaf_0_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[691]$_DFFE_PN0P_  (.RESET_B(net8049),
    .D(_11673_),
    .Q(_01260_),
    .CLK(clknet_leaf_0_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[692]$_DFFE_PN0P_  (.RESET_B(net8060),
    .D(_11671_),
    .Q(_01261_),
    .CLK(clknet_leaf_45_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[693]$_DFFE_PN0P_  (.RESET_B(net8235),
    .D(_11670_),
    .Q(_01262_),
    .CLK(clknet_leaf_37_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[694]$_DFFE_PN0P_  (.RESET_B(net8044),
    .D(_11667_),
    .Q(_01263_),
    .CLK(clknet_leaf_48_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[695]$_DFFE_PN0P_  (.RESET_B(net8150),
    .D(_11664_),
    .Q(_01264_),
    .CLK(clknet_leaf_33_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[696]$_DFFE_PN0P_  (.RESET_B(net8048),
    .D(_11661_),
    .Q(_01265_),
    .CLK(clknet_leaf_0_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[697]$_DFFE_PN0P_  (.RESET_B(net8213),
    .D(_11658_),
    .Q(_01266_),
    .CLK(clknet_leaf_20_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[698]$_DFFE_PN0P_  (.RESET_B(net8042),
    .D(_11655_),
    .Q(_01267_),
    .CLK(clknet_leaf_47_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[699]$_DFFE_PN0P_  (.RESET_B(net8102),
    .D(_11653_),
    .Q(_01268_),
    .CLK(clknet_leaf_16_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[69]$_DFFE_PN0P_  (.RESET_B(net8141),
    .D(_11651_),
    .Q(_01269_),
    .CLK(clknet_leaf_27_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[700]$_DFFE_PN0P_  (.RESET_B(net8104),
    .D(_11649_),
    .Q(_01270_),
    .CLK(clknet_leaf_25_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[701]$_DFFE_PN0P_  (.RESET_B(net8044),
    .D(_11646_),
    .Q(_01271_),
    .CLK(clknet_leaf_48_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[702]$_DFFE_PN0P_  (.RESET_B(net8128),
    .D(_11644_),
    .Q(_01272_),
    .CLK(clknet_leaf_23_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[703]$_DFFE_PN0P_  (.RESET_B(net8144),
    .D(_11641_),
    .Q(_01273_),
    .CLK(clknet_leaf_32_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[704]$_DFFE_PN0P_  (.RESET_B(net8046),
    .D(_11637_),
    .Q(_01274_),
    .CLK(clknet_leaf_47_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[705]$_DFFE_PN0P_  (.RESET_B(net8029),
    .D(_11635_),
    .Q(_01275_),
    .CLK(clknet_leaf_11_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[706]$_DFFE_PN0P_  (.RESET_B(net8089),
    .D(_11633_),
    .Q(_01276_),
    .CLK(clknet_leaf_8_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[707]$_DFFE_PN0P_  (.RESET_B(net8040),
    .D(_11631_),
    .Q(_01277_),
    .CLK(clknet_leaf_10_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[708]$_DFFE_PN0P_  (.RESET_B(net8106),
    .D(_11629_),
    .Q(_01278_),
    .CLK(clknet_leaf_26_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[709]$_DFFE_PN0P_  (.RESET_B(net8207),
    .D(_11626_),
    .Q(_01279_),
    .CLK(clknet_leaf_24_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[70]$_DFFE_PN0P_  (.RESET_B(net8099),
    .D(_11624_),
    .Q(_01280_),
    .CLK(clknet_leaf_18_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[710]$_DFFE_PN0P_  (.RESET_B(net8028),
    .D(_11621_),
    .Q(_01281_),
    .CLK(clknet_leaf_14_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[711]$_DFFE_PN0P_  (.RESET_B(net8105),
    .D(_11619_),
    .Q(_01282_),
    .CLK(clknet_leaf_28_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[712]$_DFFE_PN0P_  (.RESET_B(net8081),
    .D(_11617_),
    .Q(_01283_),
    .CLK(clknet_leaf_11_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[713]$_DFFE_PN0P_  (.RESET_B(net8032),
    .D(_11615_),
    .Q(_01284_),
    .CLK(clknet_leaf_12_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[714]$_DFFE_PN0P_  (.RESET_B(net8061),
    .D(_11613_),
    .Q(_01285_),
    .CLK(clknet_leaf_46_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[715]$_DFFE_PN0P_  (.RESET_B(net8025),
    .D(_11611_),
    .Q(_01286_),
    .CLK(clknet_leaf_14_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[716]$_DFFE_PN0P_  (.RESET_B(net8108),
    .D(_11609_),
    .Q(_01287_),
    .CLK(clknet_leaf_16_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[717]$_DFFE_PN0P_  (.RESET_B(net8104),
    .D(_11607_),
    .Q(_01288_),
    .CLK(clknet_leaf_25_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[718]$_DFFE_PN0P_  (.RESET_B(net8034),
    .D(_11605_),
    .Q(_01289_),
    .CLK(clknet_leaf_11_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[719]$_DFFE_PN0P_  (.RESET_B(net8154),
    .D(_11603_),
    .Q(_01290_),
    .CLK(clknet_leaf_32_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[71]$_DFFE_PN0P_  (.RESET_B(net8115),
    .D(_11601_),
    .Q(_01291_),
    .CLK(clknet_leaf_31_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[720]$_DFFE_PN0P_  (.RESET_B(net8043),
    .D(_11599_),
    .Q(_01292_),
    .CLK(clknet_leaf_0_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[721]$_DFFE_PN0P_  (.RESET_B(net8045),
    .D(_11596_),
    .Q(_01293_),
    .CLK(clknet_leaf_48_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[722]$_DFFE_PN0P_  (.RESET_B(net8048),
    .D(_11594_),
    .Q(_01294_),
    .CLK(clknet_leaf_0_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[723]$_DFFE_PN0P_  (.RESET_B(net8049),
    .D(_11592_),
    .Q(_01295_),
    .CLK(clknet_leaf_0_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[724]$_DFFE_PN0P_  (.RESET_B(net8060),
    .D(_11590_),
    .Q(_01296_),
    .CLK(clknet_leaf_45_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[725]$_DFFE_PN0P_  (.RESET_B(net8235),
    .D(_11589_),
    .Q(_01297_),
    .CLK(clknet_leaf_37_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[726]$_DFFE_PN0P_  (.RESET_B(net8044),
    .D(_11586_),
    .Q(_01298_),
    .CLK(clknet_leaf_48_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[727]$_DFFE_PN0P_  (.RESET_B(net8149),
    .D(_11584_),
    .Q(_01299_),
    .CLK(clknet_leaf_33_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[728]$_DFFE_PN0P_  (.RESET_B(net8048),
    .D(_11581_),
    .Q(_01300_),
    .CLK(clknet_leaf_0_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[729]$_DFFE_PN0P_  (.RESET_B(net8213),
    .D(_11579_),
    .Q(_01301_),
    .CLK(clknet_leaf_19_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[72]$_DFFE_PN0P_  (.RESET_B(net8208),
    .D(_11576_),
    .Q(_01302_),
    .CLK(clknet_leaf_20_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[730]$_DFFE_PN0P_  (.RESET_B(net8042),
    .D(_11573_),
    .Q(_01303_),
    .CLK(clknet_leaf_0_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[731]$_DFFE_PN0P_  (.RESET_B(net8102),
    .D(_11570_),
    .Q(_01304_),
    .CLK(clknet_leaf_16_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[732]$_DFFE_PN0P_  (.RESET_B(net8104),
    .D(_11568_),
    .Q(_01305_),
    .CLK(clknet_leaf_25_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[733]$_DFFE_PN0P_  (.RESET_B(net8044),
    .D(_11566_),
    .Q(_01306_),
    .CLK(clknet_leaf_48_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[734]$_DFFE_PN0P_  (.RESET_B(net8128),
    .D(_11564_),
    .Q(_01307_),
    .CLK(clknet_leaf_22_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[735]$_DFFE_PN0P_  (.RESET_B(net8144),
    .D(_11561_),
    .Q(_01308_),
    .CLK(clknet_leaf_32_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[736]$_DFFE_PN0P_  (.RESET_B(net8046),
    .D(_11557_),
    .Q(_01309_),
    .CLK(clknet_leaf_47_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[737]$_DFFE_PN0P_  (.RESET_B(net8031),
    .D(_11555_),
    .Q(_01310_),
    .CLK(clknet_leaf_11_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[738]$_DFFE_PN0P_  (.RESET_B(net8089),
    .D(_11553_),
    .Q(_01311_),
    .CLK(clknet_leaf_8_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[739]$_DFFE_PN0P_  (.RESET_B(net8040),
    .D(_11551_),
    .Q(_01312_),
    .CLK(clknet_leaf_10_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[73]$_DFFE_PN0P_  (.RESET_B(net8208),
    .D(_11548_),
    .Q(_01313_),
    .CLK(clknet_leaf_19_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[740]$_DFFE_PN0P_  (.RESET_B(net8106),
    .D(_11546_),
    .Q(_01314_),
    .CLK(clknet_leaf_25_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[741]$_DFFE_PN0P_  (.RESET_B(net8128),
    .D(_11543_),
    .Q(_01315_),
    .CLK(clknet_leaf_24_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[742]$_DFFE_PN0P_  (.RESET_B(net8033),
    .D(_11541_),
    .Q(_01316_),
    .CLK(clknet_leaf_12_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[743]$_DFFE_PN0P_  (.RESET_B(net8105),
    .D(_11539_),
    .Q(_01317_),
    .CLK(clknet_leaf_26_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[744]$_DFFE_PN0P_  (.RESET_B(net8034),
    .D(_11537_),
    .Q(_01318_),
    .CLK(clknet_leaf_11_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[745]$_DFFE_PN0P_  (.RESET_B(net8031),
    .D(_11535_),
    .Q(_01319_),
    .CLK(clknet_leaf_12_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[746]$_DFFE_PN0P_  (.RESET_B(net8061),
    .D(_11533_),
    .Q(_01320_),
    .CLK(clknet_leaf_46_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[747]$_DFFE_PN0P_  (.RESET_B(net8025),
    .D(_11531_),
    .Q(_01321_),
    .CLK(clknet_leaf_14_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[748]$_DFFE_PN0P_  (.RESET_B(net8108),
    .D(_11529_),
    .Q(_01322_),
    .CLK(clknet_leaf_16_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[749]$_DFFE_PN0P_  (.RESET_B(net8104),
    .D(_11527_),
    .Q(_01323_),
    .CLK(clknet_leaf_25_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[74]$_DFFE_PN0P_  (.RESET_B(net8224),
    .D(_11525_),
    .Q(_01324_),
    .CLK(clknet_leaf_40_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[750]$_DFFE_PN0P_  (.RESET_B(net8035),
    .D(_11522_),
    .Q(_01325_),
    .CLK(clknet_leaf_11_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[751]$_DFFE_PN0P_  (.RESET_B(net8154),
    .D(_11519_),
    .Q(_01326_),
    .CLK(clknet_leaf_32_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[752]$_DFFE_PN0P_  (.RESET_B(net8043),
    .D(_11518_),
    .Q(_01327_),
    .CLK(clknet_leaf_0_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[753]$_DFFE_PN0P_  (.RESET_B(net8045),
    .D(_11516_),
    .Q(_01328_),
    .CLK(clknet_leaf_48_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[754]$_DFFE_PN0P_  (.RESET_B(net8047),
    .D(_11514_),
    .Q(_01329_),
    .CLK(clknet_leaf_0_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[755]$_DFFE_PN0P_  (.RESET_B(net8049),
    .D(_11512_),
    .Q(_01330_),
    .CLK(clknet_leaf_0_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[756]$_DFFE_PN0P_  (.RESET_B(net8060),
    .D(_11510_),
    .Q(_01331_),
    .CLK(clknet_leaf_45_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[757]$_DFFE_PN0P_  (.RESET_B(net8229),
    .D(_11509_),
    .Q(_01332_),
    .CLK(clknet_leaf_37_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[758]$_DFFE_PN0P_  (.RESET_B(net8046),
    .D(_11506_),
    .Q(_01333_),
    .CLK(clknet_leaf_47_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[759]$_DFFE_PN0P_  (.RESET_B(net8149),
    .D(_11504_),
    .Q(_01334_),
    .CLK(clknet_leaf_33_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[75]$_DFFE_PN0P_  (.RESET_B(net8083),
    .D(_11501_),
    .Q(_01335_),
    .CLK(clknet_leaf_19_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[760]$_DFFE_PN0P_  (.RESET_B(net8045),
    .D(_11499_),
    .Q(_01336_),
    .CLK(clknet_leaf_0_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[761]$_DFFE_PN0P_  (.RESET_B(net8213),
    .D(_11497_),
    .Q(_01337_),
    .CLK(clknet_leaf_20_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[762]$_DFFE_PN0P_  (.RESET_B(net8042),
    .D(_11494_),
    .Q(_01338_),
    .CLK(clknet_leaf_47_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[763]$_DFFE_PN0P_  (.RESET_B(net8102),
    .D(_11492_),
    .Q(_01339_),
    .CLK(clknet_leaf_16_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[764]$_DFFE_PN0P_  (.RESET_B(net8104),
    .D(_11490_),
    .Q(_01340_),
    .CLK(clknet_leaf_25_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[765]$_DFFE_PN0P_  (.RESET_B(net8044),
    .D(_11488_),
    .Q(_01341_),
    .CLK(clknet_leaf_47_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[766]$_DFFE_PN0P_  (.RESET_B(net8128),
    .D(_11486_),
    .Q(_01342_),
    .CLK(clknet_leaf_22_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[767]$_DFFE_PN0P_  (.RESET_B(net8144),
    .D(_11483_),
    .Q(_01343_),
    .CLK(clknet_leaf_32_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[768]$_DFFE_PN0P_  (.RESET_B(net8041),
    .D(_11476_),
    .Q(_01344_),
    .CLK(clknet_leaf_1_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[769]$_DFFE_PN0P_  (.RESET_B(net8030),
    .D(_11473_),
    .Q(_01345_),
    .CLK(clknet_leaf_13_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[76]$_DFFE_PN0P_  (.RESET_B(net8099),
    .D(_11471_),
    .Q(_01346_),
    .CLK(clknet_leaf_18_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[770]$_DFFE_PN0P_  (.RESET_B(net8092),
    .D(_11469_),
    .Q(_01347_),
    .CLK(clknet_leaf_13_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[771]$_DFFE_PN0P_  (.RESET_B(net8079),
    .D(_11467_),
    .Q(_01348_),
    .CLK(clknet_leaf_10_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[772]$_DFFE_PN0P_  (.RESET_B(net8121),
    .D(_11465_),
    .Q(_01349_),
    .CLK(clknet_leaf_28_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[773]$_DFFE_PN0P_  (.RESET_B(net8110),
    .D(_11463_),
    .Q(_01350_),
    .CLK(clknet_leaf_26_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[774]$_DFFE_PN0P_  (.RESET_B(net8082),
    .D(_11461_),
    .Q(_01351_),
    .CLK(clknet_leaf_13_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[775]$_DFFE_PN0P_  (.RESET_B(net8121),
    .D(_11459_),
    .Q(_01352_),
    .CLK(clknet_leaf_28_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[776]$_DFFE_PN0P_  (.RESET_B(net8030),
    .D(_11457_),
    .Q(_01353_),
    .CLK(clknet_leaf_9_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[777]$_DFFE_PN0P_  (.RESET_B(net8027),
    .D(_11455_),
    .Q(_01354_),
    .CLK(clknet_leaf_14_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[778]$_DFFE_PN0P_  (.RESET_B(net8056),
    .D(_11453_),
    .Q(_01355_),
    .CLK(clknet_leaf_2_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[779]$_DFFE_PN0P_  (.RESET_B(net8025),
    .D(_11451_),
    .Q(_01356_),
    .CLK(clknet_leaf_13_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[77]$_DFFE_PN0P_  (.RESET_B(net8156),
    .D(_11449_),
    .Q(_01357_),
    .CLK(clknet_leaf_23_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[780]$_DFFE_PN0P_  (.RESET_B(net8103),
    .D(_11447_),
    .Q(_01358_),
    .CLK(clknet_leaf_17_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[781]$_DFFE_PN0P_  (.RESET_B(net8096),
    .D(_11445_),
    .Q(_01359_),
    .CLK(clknet_leaf_25_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[782]$_DFFE_PN0P_  (.RESET_B(net8079),
    .D(_11443_),
    .Q(_01360_),
    .CLK(clknet_leaf_10_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[783]$_DFFE_PN0P_  (.RESET_B(net8144),
    .D(_11441_),
    .Q(_01361_),
    .CLK(clknet_leaf_32_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[784]$_DFFE_PN0P_  (.RESET_B(net8052),
    .D(_11440_),
    .Q(_01362_),
    .CLK(clknet_leaf_4_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[785]$_DFFE_PN0P_  (.RESET_B(net8041),
    .D(_11438_),
    .Q(_01363_),
    .CLK(clknet_leaf_1_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[786]$_DFFE_PN0P_  (.RESET_B(net8038),
    .D(_11436_),
    .Q(_01364_),
    .CLK(clknet_leaf_3_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[787]$_DFFE_PN0P_  (.RESET_B(net8063),
    .D(_11434_),
    .Q(_01365_),
    .CLK(clknet_leaf_4_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[788]$_DFFE_PN0P_  (.RESET_B(net8072),
    .D(_11431_),
    .Q(_01366_),
    .CLK(clknet_leaf_5_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[789]$_DFFE_PN0P_  (.RESET_B(net8132),
    .D(_11430_),
    .Q(_01367_),
    .CLK(clknet_leaf_34_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[78]$_DFFE_PN0P_  (.RESET_B(net8211),
    .D(_11426_),
    .Q(_01368_),
    .CLK(clknet_leaf_42_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[790]$_DFFE_PN0P_  (.RESET_B(net8058),
    .D(_11424_),
    .Q(_01369_),
    .CLK(clknet_leaf_1_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[791]$_DFFE_PN0P_  (.RESET_B(net8150),
    .D(_11422_),
    .Q(_01370_),
    .CLK(clknet_leaf_33_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[792]$_DFFE_PN0P_  (.RESET_B(net8064),
    .D(_11419_),
    .Q(_01371_),
    .CLK(clknet_leaf_2_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[793]$_DFFE_PN0P_  (.RESET_B(net8228),
    .D(_11417_),
    .Q(_01372_),
    .CLK(clknet_leaf_21_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[794]$_DFFE_PN0P_  (.RESET_B(net8057),
    .D(_11413_),
    .Q(_01373_),
    .CLK(clknet_leaf_4_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[795]$_DFFE_PN0P_  (.RESET_B(net8103),
    .D(_11411_),
    .Q(_01374_),
    .CLK(clknet_leaf_17_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[796]$_DFFE_PN0P_  (.RESET_B(net8120),
    .D(_11409_),
    .Q(_01375_),
    .CLK(clknet_leaf_25_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[797]$_DFFE_PN0P_  (.RESET_B(net8038),
    .D(_11407_),
    .Q(_01376_),
    .CLK(clknet_leaf_2_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[798]$_DFFE_PN0P_  (.RESET_B(net8126),
    .D(_11405_),
    .Q(_01377_),
    .CLK(clknet_leaf_23_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[799]$_DFFE_PN0P_  (.RESET_B(net8144),
    .D(_11402_),
    .Q(_01378_),
    .CLK(clknet_leaf_32_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[79]$_DFFE_PN0P_  (.RESET_B(net8135),
    .D(_11397_),
    .Q(_01379_),
    .CLK(clknet_leaf_37_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[800]$_DFFE_PN0P_  (.RESET_B(net8041),
    .D(_11396_),
    .Q(_01380_),
    .CLK(clknet_leaf_1_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[801]$_DFFE_PN0P_  (.RESET_B(net8030),
    .D(_11394_),
    .Q(_01381_),
    .CLK(clknet_leaf_12_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[802]$_DFFE_PN0P_  (.RESET_B(net8092),
    .D(_11392_),
    .Q(_01382_),
    .CLK(clknet_leaf_13_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[803]$_DFFE_PN0P_  (.RESET_B(net8051),
    .D(_11390_),
    .Q(_01383_),
    .CLK(clknet_leaf_10_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[804]$_DFFE_PN0P_  (.RESET_B(net8122),
    .D(_11388_),
    .Q(_01384_),
    .CLK(clknet_leaf_28_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[805]$_DFFE_PN0P_  (.RESET_B(net8110),
    .D(_11386_),
    .Q(_01385_),
    .CLK(clknet_leaf_26_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[806]$_DFFE_PN0P_  (.RESET_B(net8082),
    .D(_11384_),
    .Q(_01386_),
    .CLK(clknet_leaf_14_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[807]$_DFFE_PN0P_  (.RESET_B(net8123),
    .D(_11382_),
    .Q(_01387_),
    .CLK(clknet_leaf_28_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[808]$_DFFE_PN0P_  (.RESET_B(net8030),
    .D(_11380_),
    .Q(_01388_),
    .CLK(clknet_leaf_9_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[809]$_DFFE_PN0P_  (.RESET_B(net8027),
    .D(_11378_),
    .Q(_01389_),
    .CLK(clknet_leaf_14_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[80]$_DFFE_PN0P_  (.RESET_B(net8211),
    .D(_11376_),
    .Q(_01390_),
    .CLK(clknet_leaf_42_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[810]$_DFFE_PN0P_  (.RESET_B(net8056),
    .D(_11374_),
    .Q(_01391_),
    .CLK(clknet_leaf_2_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[811]$_DFFE_PN0P_  (.RESET_B(net8025),
    .D(_11372_),
    .Q(_01392_),
    .CLK(clknet_leaf_14_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[812]$_DFFE_PN0P_  (.RESET_B(net8103),
    .D(_11370_),
    .Q(_01393_),
    .CLK(clknet_leaf_17_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[813]$_DFFE_PN0P_  (.RESET_B(net8096),
    .D(_11368_),
    .Q(_01394_),
    .CLK(clknet_leaf_25_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[814]$_DFFE_PN0P_  (.RESET_B(net8079),
    .D(_11365_),
    .Q(_01395_),
    .CLK(clknet_leaf_9_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[815]$_DFFE_PN0P_  (.RESET_B(net8146),
    .D(_11363_),
    .Q(_01396_),
    .CLK(clknet_leaf_32_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[816]$_DFFE_PN0P_  (.RESET_B(net8052),
    .D(_11362_),
    .Q(_01397_),
    .CLK(clknet_leaf_4_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[817]$_DFFE_PN0P_  (.RESET_B(net8054),
    .D(_11360_),
    .Q(_01398_),
    .CLK(clknet_leaf_1_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[818]$_DFFE_PN0P_  (.RESET_B(net8039),
    .D(_11358_),
    .Q(_01399_),
    .CLK(clknet_leaf_3_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[819]$_DFFE_PN0P_  (.RESET_B(net8063),
    .D(_11356_),
    .Q(_01400_),
    .CLK(clknet_leaf_4_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[81]$_DFFE_PN0P_  (.RESET_B(net8220),
    .D(_11354_),
    .Q(_01401_),
    .CLK(clknet_leaf_41_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[820]$_DFFE_PN0P_  (.RESET_B(net8072),
    .D(_11351_),
    .Q(_01402_),
    .CLK(clknet_leaf_2_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[821]$_DFFE_PN0P_  (.RESET_B(net8132),
    .D(_11350_),
    .Q(_01403_),
    .CLK(clknet_leaf_34_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[822]$_DFFE_PN0P_  (.RESET_B(net8058),
    .D(_11347_),
    .Q(_01404_),
    .CLK(clknet_leaf_47_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[823]$_DFFE_PN0P_  (.RESET_B(net8150),
    .D(_11345_),
    .Q(_01405_),
    .CLK(clknet_leaf_33_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[824]$_DFFE_PN0P_  (.RESET_B(net8055),
    .D(_11342_),
    .Q(_01406_),
    .CLK(clknet_leaf_3_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[825]$_DFFE_PN0P_  (.RESET_B(net8237),
    .D(_11340_),
    .Q(_01407_),
    .CLK(clknet_leaf_21_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[826]$_DFFE_PN0P_  (.RESET_B(net8063),
    .D(_11337_),
    .Q(_01408_),
    .CLK(clknet_leaf_4_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[827]$_DFFE_PN0P_  (.RESET_B(net8103),
    .D(_11335_),
    .Q(_01409_),
    .CLK(clknet_leaf_17_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[828]$_DFFE_PN0P_  (.RESET_B(net8120),
    .D(_11333_),
    .Q(_01410_),
    .CLK(clknet_leaf_26_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[829]$_DFFE_PN0P_  (.RESET_B(net8055),
    .D(_11331_),
    .Q(_01411_),
    .CLK(clknet_leaf_3_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[82]$_DFFE_PN0P_  (.RESET_B(net8223),
    .D(_11329_),
    .Q(_01412_),
    .CLK(clknet_leaf_40_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[830]$_DFFE_PN0P_  (.RESET_B(net8126),
    .D(_11327_),
    .Q(_01413_),
    .CLK(clknet_leaf_23_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[831]$_DFFE_PN0P_  (.RESET_B(net8144),
    .D(_11324_),
    .Q(_01414_),
    .CLK(clknet_leaf_32_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[832]$_DFFE_PN0P_  (.RESET_B(net8054),
    .D(_11320_),
    .Q(_01415_),
    .CLK(clknet_leaf_1_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[833]$_DFFE_PN0P_  (.RESET_B(net8031),
    .D(_11318_),
    .Q(_01416_),
    .CLK(clknet_leaf_13_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[834]$_DFFE_PN0P_  (.RESET_B(net8086),
    .D(_11316_),
    .Q(_01417_),
    .CLK(clknet_leaf_13_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[835]$_DFFE_PN0P_  (.RESET_B(net8051),
    .D(_11314_),
    .Q(_01418_),
    .CLK(clknet_leaf_10_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[836]$_DFFE_PN0P_  (.RESET_B(net8121),
    .D(_11312_),
    .Q(_01419_),
    .CLK(clknet_leaf_28_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[837]$_DFFE_PN0P_  (.RESET_B(net8119),
    .D(_11310_),
    .Q(_01420_),
    .CLK(clknet_leaf_27_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[838]$_DFFE_PN0P_  (.RESET_B(net8082),
    .D(_11308_),
    .Q(_01421_),
    .CLK(clknet_leaf_14_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[839]$_DFFE_PN0P_  (.RESET_B(net8122),
    .D(_11306_),
    .Q(_01422_),
    .CLK(clknet_leaf_28_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[83]$_DFFE_PN0P_  (.RESET_B(net8214),
    .D(_11303_),
    .Q(_01423_),
    .CLK(clknet_leaf_41_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[840]$_DFFE_PN0P_  (.RESET_B(net8030),
    .D(_11301_),
    .Q(_01424_),
    .CLK(clknet_leaf_13_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[841]$_DFFE_PN0P_  (.RESET_B(net8026),
    .D(_11299_),
    .Q(_01425_),
    .CLK(clknet_leaf_13_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[842]$_DFFE_PN0P_  (.RESET_B(net8062),
    .D(_11297_),
    .Q(_01426_),
    .CLK(clknet_leaf_2_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[843]$_DFFE_PN0P_  (.RESET_B(net8025),
    .D(_11295_),
    .Q(_01427_),
    .CLK(clknet_leaf_13_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[844]$_DFFE_PN0P_  (.RESET_B(net8107),
    .D(_11292_),
    .Q(_01428_),
    .CLK(clknet_leaf_17_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[845]$_DFFE_PN0P_  (.RESET_B(net8096),
    .D(_11290_),
    .Q(_01429_),
    .CLK(clknet_leaf_24_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[846]$_DFFE_PN0P_  (.RESET_B(net8079),
    .D(_11288_),
    .Q(_01430_),
    .CLK(clknet_leaf_9_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[847]$_DFFE_PN0P_  (.RESET_B(net8146),
    .D(_11286_),
    .Q(_01431_),
    .CLK(clknet_leaf_32_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[848]$_DFFE_PN0P_  (.RESET_B(net8052),
    .D(_11285_),
    .Q(_01432_),
    .CLK(clknet_leaf_4_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[849]$_DFFE_PN0P_  (.RESET_B(net8054),
    .D(_11283_),
    .Q(_01433_),
    .CLK(clknet_leaf_1_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[84]$_DFFE_PN0P_  (.RESET_B(net8234),
    .D(_11280_),
    .Q(_01434_),
    .CLK(clknet_leaf_40_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[850]$_DFFE_PN0P_  (.RESET_B(net8054),
    .D(_11279_),
    .Q(_01435_),
    .CLK(clknet_leaf_2_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[851]$_DFFE_PN0P_  (.RESET_B(net8052),
    .D(_11277_),
    .Q(_01436_),
    .CLK(clknet_leaf_4_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[852]$_DFFE_PN0P_  (.RESET_B(net8072),
    .D(_11275_),
    .Q(_01437_),
    .CLK(clknet_leaf_5_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[853]$_DFFE_PN0P_  (.RESET_B(net8132),
    .D(_11273_),
    .Q(_01438_),
    .CLK(clknet_leaf_34_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[854]$_DFFE_PN0P_  (.RESET_B(net8059),
    .D(_11269_),
    .Q(_01439_),
    .CLK(clknet_leaf_46_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[855]$_DFFE_PN0P_  (.RESET_B(net8148),
    .D(_11267_),
    .Q(_01440_),
    .CLK(clknet_leaf_33_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[856]$_DFFE_PN0P_  (.RESET_B(net8064),
    .D(_11264_),
    .Q(_01441_),
    .CLK(clknet_leaf_3_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[857]$_DFFE_PN0P_  (.RESET_B(net8228),
    .D(_11262_),
    .Q(_01442_),
    .CLK(clknet_leaf_21_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[858]$_DFFE_PN0P_  (.RESET_B(net8063),
    .D(_11259_),
    .Q(_01443_),
    .CLK(clknet_leaf_4_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[859]$_DFFE_PN0P_  (.RESET_B(net8097),
    .D(_11257_),
    .Q(_01444_),
    .CLK(clknet_leaf_17_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[85]$_DFFE_PN0P_  (.RESET_B(net8229),
    .D(_11255_),
    .Q(_01445_),
    .CLK(clknet_leaf_36_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[860]$_DFFE_PN0P_  (.RESET_B(net8119),
    .D(_11252_),
    .Q(_01446_),
    .CLK(clknet_leaf_25_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[861]$_DFFE_PN0P_  (.RESET_B(net8054),
    .D(_11250_),
    .Q(_01447_),
    .CLK(clknet_leaf_2_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[862]$_DFFE_PN0P_  (.RESET_B(net8126),
    .D(_11248_),
    .Q(_01448_),
    .CLK(clknet_leaf_22_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[863]$_DFFE_PN0P_  (.RESET_B(net8144),
    .D(_11245_),
    .Q(_01449_),
    .CLK(clknet_leaf_32_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[864]$_DFFE_PN0P_  (.RESET_B(net8041),
    .D(_11241_),
    .Q(_01450_),
    .CLK(clknet_leaf_1_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[865]$_DFFE_PN0P_  (.RESET_B(net8030),
    .D(_11239_),
    .Q(_01451_),
    .CLK(clknet_leaf_12_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[866]$_DFFE_PN0P_  (.RESET_B(net8092),
    .D(_11237_),
    .Q(_01452_),
    .CLK(clknet_leaf_13_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[867]$_DFFE_PN0P_  (.RESET_B(net8051),
    .D(_11235_),
    .Q(_01453_),
    .CLK(clknet_leaf_10_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[868]$_DFFE_PN0P_  (.RESET_B(net8121),
    .D(_11233_),
    .Q(_01454_),
    .CLK(clknet_leaf_28_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[869]$_DFFE_PN0P_  (.RESET_B(net8119),
    .D(_11231_),
    .Q(_01455_),
    .CLK(clknet_leaf_27_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[86]$_DFFE_PN0P_  (.RESET_B(net8222),
    .D(_11229_),
    .Q(_01456_),
    .CLK(clknet_leaf_39_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[870]$_DFFE_PN0P_  (.RESET_B(net8082),
    .D(_11227_),
    .Q(_01457_),
    .CLK(clknet_leaf_14_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[871]$_DFFE_PN0P_  (.RESET_B(net8122),
    .D(_11225_),
    .Q(_01458_),
    .CLK(clknet_leaf_29_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[872]$_DFFE_PN0P_  (.RESET_B(net8030),
    .D(_11222_),
    .Q(_01459_),
    .CLK(clknet_leaf_12_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[873]$_DFFE_PN0P_  (.RESET_B(net8026),
    .D(_11220_),
    .Q(_01460_),
    .CLK(clknet_leaf_14_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[874]$_DFFE_PN0P_  (.RESET_B(net8062),
    .D(_11218_),
    .Q(_01461_),
    .CLK(clknet_leaf_2_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[875]$_DFFE_PN0P_  (.RESET_B(net8025),
    .D(_11216_),
    .Q(_01462_),
    .CLK(clknet_leaf_14_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[876]$_DFFE_PN0P_  (.RESET_B(net8107),
    .D(_11214_),
    .Q(_01463_),
    .CLK(clknet_leaf_17_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[877]$_DFFE_PN0P_  (.RESET_B(net8096),
    .D(_11212_),
    .Q(_01464_),
    .CLK(clknet_leaf_24_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[878]$_DFFE_PN0P_  (.RESET_B(net8067),
    .D(_11210_),
    .Q(_01465_),
    .CLK(clknet_leaf_10_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[879]$_DFFE_PN0P_  (.RESET_B(net8146),
    .D(_11208_),
    .Q(_01466_),
    .CLK(clknet_leaf_32_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[87]$_DFFE_PN0P_  (.RESET_B(net8135),
    .D(_11207_),
    .Q(_01467_),
    .CLK(clknet_leaf_37_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[880]$_DFFE_PN0P_  (.RESET_B(net8052),
    .D(_11203_),
    .Q(_01468_),
    .CLK(clknet_leaf_4_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[881]$_DFFE_PN0P_  (.RESET_B(net8054),
    .D(_11201_),
    .Q(_01469_),
    .CLK(clknet_leaf_1_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[882]$_DFFE_PN0P_  (.RESET_B(net8054),
    .D(_11199_),
    .Q(_01470_),
    .CLK(clknet_leaf_2_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[883]$_DFFE_PN0P_  (.RESET_B(net8063),
    .D(_11197_),
    .Q(_01471_),
    .CLK(clknet_leaf_4_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[884]$_DFFE_PN0P_  (.RESET_B(net8072),
    .D(_11195_),
    .Q(_01472_),
    .CLK(clknet_leaf_5_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[885]$_DFFE_PN0P_  (.RESET_B(net8132),
    .D(_11193_),
    .Q(_01473_),
    .CLK(clknet_leaf_35_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[886]$_DFFE_PN0P_  (.RESET_B(net8058),
    .D(_11190_),
    .Q(_01474_),
    .CLK(clknet_leaf_47_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[887]$_DFFE_PN0P_  (.RESET_B(net8150),
    .D(_11188_),
    .Q(_01475_),
    .CLK(clknet_leaf_33_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[888]$_DFFE_PN0P_  (.RESET_B(net8064),
    .D(_11185_),
    .Q(_01476_),
    .CLK(clknet_leaf_3_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[889]$_DFFE_PN0P_  (.RESET_B(net8228),
    .D(_11183_),
    .Q(_01477_),
    .CLK(clknet_leaf_21_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[88]$_DFFE_PN0P_  (.RESET_B(net8215),
    .D(_11179_),
    .Q(_01478_),
    .CLK(clknet_leaf_42_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[890]$_DFFE_PN0P_  (.RESET_B(net8063),
    .D(_11177_),
    .Q(_01479_),
    .CLK(clknet_leaf_4_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[891]$_DFFE_PN0P_  (.RESET_B(net8097),
    .D(_11175_),
    .Q(_01480_),
    .CLK(clknet_leaf_17_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[892]$_DFFE_PN0P_  (.RESET_B(net8119),
    .D(_11173_),
    .Q(_01481_),
    .CLK(clknet_leaf_25_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[893]$_DFFE_PN0P_  (.RESET_B(net8055),
    .D(_11170_),
    .Q(_01482_),
    .CLK(clknet_leaf_2_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[894]$_DFFE_PN0P_  (.RESET_B(net8140),
    .D(_11167_),
    .Q(_01483_),
    .CLK(clknet_leaf_22_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[895]$_DFFE_PN0P_  (.RESET_B(net8144),
    .D(_11163_),
    .Q(_01484_),
    .CLK(clknet_leaf_32_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[896]$_DFFE_PN0P_  (.RESET_B(net8041),
    .D(_11157_),
    .Q(_01485_),
    .CLK(clknet_leaf_1_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[897]$_DFFE_PN0P_  (.RESET_B(net8029),
    .D(_11155_),
    .Q(_01486_),
    .CLK(clknet_leaf_12_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[898]$_DFFE_PN0P_  (.RESET_B(net8091),
    .D(_11153_),
    .Q(_01487_),
    .CLK(clknet_leaf_12_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[899]$_DFFE_PN0P_  (.RESET_B(net8051),
    .D(_11151_),
    .Q(_01488_),
    .CLK(clknet_leaf_4_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[89]$_DFFE_PN0P_  (.RESET_B(net8227),
    .D(_11148_),
    .Q(_01489_),
    .CLK(clknet_leaf_21_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[900]$_DFFE_PN0P_  (.RESET_B(net8122),
    .D(_11144_),
    .Q(_01490_),
    .CLK(clknet_leaf_29_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[901]$_DFFE_PN0P_  (.RESET_B(net8110),
    .D(_11142_),
    .Q(_01491_),
    .CLK(clknet_leaf_27_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[902]$_DFFE_PN0P_  (.RESET_B(net8023),
    .D(_11140_),
    .Q(_01492_),
    .CLK(clknet_leaf_15_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[903]$_DFFE_PN0P_  (.RESET_B(net8122),
    .D(_11138_),
    .Q(_01493_),
    .CLK(clknet_leaf_29_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[904]$_DFFE_PN0P_  (.RESET_B(net8033),
    .D(_11135_),
    .Q(_01494_),
    .CLK(clknet_leaf_11_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[905]$_DFFE_PN0P_  (.RESET_B(net8026),
    .D(_11133_),
    .Q(_01495_),
    .CLK(clknet_leaf_15_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[906]$_DFFE_PN0P_  (.RESET_B(net8056),
    .D(_11131_),
    .Q(_01496_),
    .CLK(clknet_leaf_2_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[907]$_DFFE_PN0P_  (.RESET_B(net8024),
    .D(_11129_),
    .Q(_01497_),
    .CLK(clknet_leaf_14_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[908]$_DFFE_PN0P_  (.RESET_B(net8098),
    .D(_11127_),
    .Q(_01498_),
    .CLK(clknet_leaf_17_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[909]$_DFFE_PN0P_  (.RESET_B(net8120),
    .D(_11124_),
    .Q(_01499_),
    .CLK(clknet_leaf_25_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[90]$_DFFE_PN0P_  (.RESET_B(net8214),
    .D(_11122_),
    .Q(_01500_),
    .CLK(clknet_leaf_41_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[910]$_DFFE_PN0P_  (.RESET_B(net8080),
    .D(_11120_),
    .Q(_01501_),
    .CLK(clknet_leaf_10_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[911]$_DFFE_PN0P_  (.RESET_B(net8155),
    .D(_11118_),
    .Q(_01502_),
    .CLK(clknet_leaf_33_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[912]$_DFFE_PN0P_  (.RESET_B(net8053),
    .D(_11117_),
    .Q(_01503_),
    .CLK(clknet_leaf_4_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[913]$_DFFE_PN0P_  (.RESET_B(net8050),
    .D(_11115_),
    .Q(_01504_),
    .CLK(clknet_leaf_1_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[914]$_DFFE_PN0P_  (.RESET_B(net8039),
    .D(_11113_),
    .Q(_01505_),
    .CLK(clknet_leaf_3_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[915]$_DFFE_PN0P_  (.RESET_B(net8057),
    .D(_11111_),
    .Q(_01506_),
    .CLK(clknet_leaf_5_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[916]$_DFFE_PN0P_  (.RESET_B(net8076),
    .D(_11109_),
    .Q(_01507_),
    .CLK(clknet_leaf_5_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[917]$_DFFE_PN0P_  (.RESET_B(net8140),
    .D(_11107_),
    .Q(_01508_),
    .CLK(clknet_leaf_35_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[918]$_DFFE_PN0P_  (.RESET_B(net8059),
    .D(_11104_),
    .Q(_01509_),
    .CLK(clknet_leaf_1_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[919]$_DFFE_PN0P_  (.RESET_B(net8130),
    .D(_11101_),
    .Q(_01510_),
    .CLK(clknet_leaf_34_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[91]$_DFFE_PN0P_  (.RESET_B(net8126),
    .D(_11098_),
    .Q(_01511_),
    .CLK(clknet_leaf_23_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[920]$_DFFE_PN0P_  (.RESET_B(net8055),
    .D(_11096_),
    .Q(_01512_),
    .CLK(clknet_leaf_3_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[921]$_DFFE_PN0P_  (.RESET_B(net8237),
    .D(_11094_),
    .Q(_01513_),
    .CLK(clknet_leaf_22_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[922]$_DFFE_PN0P_  (.RESET_B(net8056),
    .D(_11091_),
    .Q(_01514_),
    .CLK(clknet_leaf_2_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[923]$_DFFE_PN0P_  (.RESET_B(net8097),
    .D(_11088_),
    .Q(_01515_),
    .CLK(clknet_leaf_17_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[924]$_DFFE_PN0P_  (.RESET_B(net8120),
    .D(_11086_),
    .Q(_01516_),
    .CLK(clknet_leaf_25_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[925]$_DFFE_PN0P_  (.RESET_B(net8038),
    .D(_11083_),
    .Q(_01517_),
    .CLK(clknet_leaf_3_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[926]$_DFFE_PN0P_  (.RESET_B(net8141),
    .D(_11081_),
    .Q(_01518_),
    .CLK(clknet_leaf_22_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[927]$_DFFE_PN0P_  (.RESET_B(net8163),
    .D(_11078_),
    .Q(_01519_),
    .CLK(clknet_leaf_31_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[928]$_DFFE_PN0P_  (.RESET_B(net8041),
    .D(_11073_),
    .Q(_01520_),
    .CLK(clknet_leaf_1_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[929]$_DFFE_PN0P_  (.RESET_B(net8031),
    .D(_11071_),
    .Q(_01521_),
    .CLK(clknet_leaf_12_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[92]$_DFFE_PN0P_  (.RESET_B(net8117),
    .D(_11069_),
    .Q(_01522_),
    .CLK(clknet_leaf_29_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[930]$_DFFE_PN0P_  (.RESET_B(net8091),
    .D(_11067_),
    .Q(_01523_),
    .CLK(clknet_leaf_13_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[931]$_DFFE_PN0P_  (.RESET_B(net8053),
    .D(_11065_),
    .Q(_01524_),
    .CLK(clknet_leaf_4_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[932]$_DFFE_PN0P_  (.RESET_B(net8122),
    .D(_11062_),
    .Q(_01525_),
    .CLK(clknet_leaf_29_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[933]$_DFFE_PN0P_  (.RESET_B(net8119),
    .D(_11059_),
    .Q(_01526_),
    .CLK(clknet_leaf_27_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[934]$_DFFE_PN0P_  (.RESET_B(net8023),
    .D(_11057_),
    .Q(_01527_),
    .CLK(clknet_leaf_15_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[935]$_DFFE_PN0P_  (.RESET_B(net8122),
    .D(_11055_),
    .Q(_01528_),
    .CLK(clknet_leaf_29_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[936]$_DFFE_PN0P_  (.RESET_B(net8030),
    .D(_11053_),
    .Q(_01529_),
    .CLK(clknet_leaf_11_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[937]$_DFFE_PN0P_  (.RESET_B(net8026),
    .D(_11051_),
    .Q(_01530_),
    .CLK(clknet_leaf_15_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[938]$_DFFE_PN0P_  (.RESET_B(net8056),
    .D(_11049_),
    .Q(_01531_),
    .CLK(clknet_leaf_2_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[939]$_DFFE_PN0P_  (.RESET_B(net8024),
    .D(_11047_),
    .Q(_01532_),
    .CLK(clknet_leaf_14_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[93]$_DFFE_PN0P_  (.RESET_B(net8221),
    .D(_11044_),
    .Q(_01533_),
    .CLK(clknet_leaf_39_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[940]$_DFFE_PN0P_  (.RESET_B(net8098),
    .D(_11042_),
    .Q(_01534_),
    .CLK(clknet_leaf_17_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[941]$_DFFE_PN0P_  (.RESET_B(net8120),
    .D(_11039_),
    .Q(_01535_),
    .CLK(clknet_leaf_25_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[942]$_DFFE_PN0P_  (.RESET_B(net8079),
    .D(_11037_),
    .Q(_01536_),
    .CLK(clknet_leaf_10_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[943]$_DFFE_PN0P_  (.RESET_B(net8155),
    .D(_11035_),
    .Q(_01537_),
    .CLK(clknet_leaf_33_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[944]$_DFFE_PN0P_  (.RESET_B(net8053),
    .D(_11034_),
    .Q(_01538_),
    .CLK(clknet_leaf_4_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[945]$_DFFE_PN0P_  (.RESET_B(net8050),
    .D(_11032_),
    .Q(_01539_),
    .CLK(clknet_leaf_1_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[946]$_DFFE_PN0P_  (.RESET_B(net8039),
    .D(_11030_),
    .Q(_01540_),
    .CLK(clknet_leaf_3_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[947]$_DFFE_PN0P_  (.RESET_B(net8057),
    .D(_11028_),
    .Q(_01541_),
    .CLK(clknet_leaf_5_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[948]$_DFFE_PN0P_  (.RESET_B(net8076),
    .D(_11026_),
    .Q(_01542_),
    .CLK(clknet_leaf_5_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[949]$_DFFE_PN0P_  (.RESET_B(net8139),
    .D(_11025_),
    .Q(_01543_),
    .CLK(clknet_leaf_35_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[94]$_DFFE_PN0P_  (.RESET_B(net8131),
    .D(_11021_),
    .Q(_01544_),
    .CLK(clknet_leaf_34_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[950]$_DFFE_PN0P_  (.RESET_B(net8059),
    .D(_11018_),
    .Q(_01545_),
    .CLK(clknet_leaf_2_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[951]$_DFFE_PN0P_  (.RESET_B(net8129),
    .D(_11015_),
    .Q(_01546_),
    .CLK(clknet_leaf_34_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[952]$_DFFE_PN0P_  (.RESET_B(net8055),
    .D(_11012_),
    .Q(_01547_),
    .CLK(clknet_leaf_3_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[953]$_DFFE_PN0P_  (.RESET_B(net8237),
    .D(_11010_),
    .Q(_01548_),
    .CLK(clknet_leaf_22_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[954]$_DFFE_PN0P_  (.RESET_B(net8057),
    .D(_11007_),
    .Q(_01549_),
    .CLK(clknet_leaf_2_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[955]$_DFFE_PN0P_  (.RESET_B(net8097),
    .D(_11005_),
    .Q(_01550_),
    .CLK(clknet_leaf_17_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[956]$_DFFE_PN0P_  (.RESET_B(net8119),
    .D(_11003_),
    .Q(_01551_),
    .CLK(clknet_leaf_26_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[957]$_DFFE_PN0P_  (.RESET_B(net8038),
    .D(_11000_),
    .Q(_01552_),
    .CLK(clknet_leaf_3_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[958]$_DFFE_PN0P_  (.RESET_B(net8141),
    .D(_10997_),
    .Q(_01553_),
    .CLK(clknet_leaf_22_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[959]$_DFFE_PN0P_  (.RESET_B(net8163),
    .D(_10994_),
    .Q(_01554_),
    .CLK(clknet_leaf_31_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[95]$_DFFE_PN0P_  (.RESET_B(net8147),
    .D(_10988_),
    .Q(_01555_),
    .CLK(clknet_leaf_33_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[960]$_DFFE_PN0P_  (.RESET_B(net8041),
    .D(_10983_),
    .Q(_01556_),
    .CLK(clknet_leaf_0_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[961]$_DFFE_PN0P_  (.RESET_B(net8029),
    .D(_10979_),
    .Q(_01557_),
    .CLK(clknet_leaf_12_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[962]$_DFFE_PN0P_  (.RESET_B(net8091),
    .D(_10977_),
    .Q(_01558_),
    .CLK(clknet_leaf_13_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[963]$_DFFE_PN0P_  (.RESET_B(net8051),
    .D(_10975_),
    .Q(_01559_),
    .CLK(clknet_leaf_10_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[964]$_DFFE_PN0P_  (.RESET_B(net8121),
    .D(_10972_),
    .Q(_01560_),
    .CLK(clknet_leaf_28_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[965]$_DFFE_PN0P_  (.RESET_B(net8119),
    .D(_10969_),
    .Q(_01561_),
    .CLK(clknet_leaf_26_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[966]$_DFFE_PN0P_  (.RESET_B(net8023),
    .D(_10967_),
    .Q(_01562_),
    .CLK(clknet_leaf_15_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[967]$_DFFE_PN0P_  (.RESET_B(net8121),
    .D(_10965_),
    .Q(_01563_),
    .CLK(clknet_leaf_28_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[968]$_DFFE_PN0P_  (.RESET_B(net8091),
    .D(_10963_),
    .Q(_01564_),
    .CLK(clknet_leaf_9_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[969]$_DFFE_PN0P_  (.RESET_B(net8026),
    .D(_10930_),
    .Q(_01565_),
    .CLK(clknet_leaf_13_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[96]$_DFFE_PN0P_  (.RESET_B(net8231),
    .D(_10896_),
    .Q(_01566_),
    .CLK(clknet_leaf_40_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[970]$_DFFE_PN0P_  (.RESET_B(net8056),
    .D(_10894_),
    .Q(_01567_),
    .CLK(clknet_leaf_2_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[971]$_DFFE_PN0P_  (.RESET_B(net8024),
    .D(_10859_),
    .Q(_01568_),
    .CLK(clknet_leaf_14_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[972]$_DFFE_PN0P_  (.RESET_B(net8098),
    .D(_10823_),
    .Q(_01569_),
    .CLK(clknet_leaf_17_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[973]$_DFFE_PN0P_  (.RESET_B(net8096),
    .D(_10791_),
    .Q(_01570_),
    .CLK(clknet_leaf_24_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[974]$_DFFE_PN0P_  (.RESET_B(net8067),
    .D(_10759_),
    .Q(_01571_),
    .CLK(clknet_leaf_9_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[975]$_DFFE_PN0P_  (.RESET_B(net8155),
    .D(_10725_),
    .Q(_01572_),
    .CLK(clknet_leaf_33_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[976]$_DFFE_PN0P_  (.RESET_B(net8051),
    .D(_10694_),
    .Q(_01573_),
    .CLK(clknet_leaf_4_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[977]$_DFFE_PN0P_  (.RESET_B(net8038),
    .D(_10653_),
    .Q(_01574_),
    .CLK(clknet_leaf_1_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[978]$_DFFE_PN0P_  (.RESET_B(net8039),
    .D(_10616_),
    .Q(_01575_),
    .CLK(clknet_leaf_3_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[979]$_DFFE_PN0P_  (.RESET_B(net8057),
    .D(_10573_),
    .Q(_01576_),
    .CLK(clknet_leaf_5_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[97]$_DFFE_PN0P_  (.RESET_B(net8210),
    .D(_10535_),
    .Q(_01577_),
    .CLK(clknet_leaf_20_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[980]$_DFFE_PN0P_  (.RESET_B(net8212),
    .D(_10533_),
    .Q(_01578_),
    .CLK(clknet_leaf_42_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[981]$_DFFE_PN0P_  (.RESET_B(net8140),
    .D(_10495_),
    .Q(_01579_),
    .CLK(clknet_leaf_35_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[982]$_DFFE_PN0P_  (.RESET_B(net8059),
    .D(_10457_),
    .Q(_01580_),
    .CLK(clknet_leaf_1_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[983]$_DFFE_PN0P_  (.RESET_B(net8138),
    .D(_10418_),
    .Q(_01581_),
    .CLK(clknet_leaf_35_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[984]$_DFFE_PN0P_  (.RESET_B(net8055),
    .D(_10374_),
    .Q(_01582_),
    .CLK(clknet_leaf_3_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[985]$_DFFE_PN0P_  (.RESET_B(net8228),
    .D(_10343_),
    .Q(_01583_),
    .CLK(clknet_leaf_21_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[986]$_DFFE_PN0P_  (.RESET_B(net8057),
    .D(_10309_),
    .Q(_01584_),
    .CLK(clknet_leaf_2_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[987]$_DFFE_PN0P_  (.RESET_B(net8097),
    .D(_10270_),
    .Q(_01585_),
    .CLK(clknet_leaf_17_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[988]$_DFFE_PN0P_  (.RESET_B(net8110),
    .D(_10237_),
    .Q(_01586_),
    .CLK(clknet_leaf_26_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[989]$_DFFE_PN0P_  (.RESET_B(net8038),
    .D(_10205_),
    .Q(_01587_),
    .CLK(clknet_leaf_3_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[98]$_DFFE_PN0P_  (.RESET_B(net8237),
    .D(_10168_),
    .Q(_01588_),
    .CLK(clknet_leaf_20_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[990]$_DFFE_PN0P_  (.RESET_B(net8131),
    .D(_10166_),
    .Q(_01589_),
    .CLK(clknet_leaf_22_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[991]$_DFFE_PN0P_  (.RESET_B(net8157),
    .D(_10133_),
    .Q(_01590_),
    .CLK(clknet_leaf_31_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[992]$_DFFE_PN0P_  (.RESET_B(net8050),
    .D(_10090_),
    .Q(_01591_),
    .CLK(clknet_leaf_0_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[993]$_DFFE_PN0P_  (.RESET_B(net8031),
    .D(_10024_),
    .Q(_01592_),
    .CLK(clknet_leaf_12_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[994]$_DFFE_PN0P_  (.RESET_B(net8091),
    .D(_09963_),
    .Q(_01593_),
    .CLK(clknet_leaf_12_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[995]$_DFFE_PN0P_  (.RESET_B(net8051),
    .D(_09906_),
    .Q(_01594_),
    .CLK(clknet_leaf_4_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[996]$_DFFE_PN0P_  (.RESET_B(net8121),
    .D(_09904_),
    .Q(_01595_),
    .CLK(clknet_leaf_28_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[997]$_DFFE_PN0P_  (.RESET_B(net8119),
    .D(_09843_),
    .Q(_01596_),
    .CLK(clknet_leaf_26_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[998]$_DFFE_PN0P_  (.RESET_B(net8023),
    .D(_09776_),
    .Q(_01597_),
    .CLK(clknet_leaf_14_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[999]$_DFFE_PN0P_  (.RESET_B(net8121),
    .D(_09688_),
    .Q(_01598_),
    .CLK(clknet_leaf_28_clk_i_regs));
 sg13g2_dfrbpq_1 \gen_regfile_ff.register_file_i.rf_reg[99]$_DFFE_PN0P_  (.RESET_B(net8210),
    .D(_09613_),
    .Q(_01599_),
    .CLK(clknet_leaf_21_clk_i_regs));
 sg13g2_dfrbpq_1 \id_stage_i.branch_set$_DFF_PN0_  (.RESET_B(net8238),
    .D(_07040_),
    .Q(\id_stage_i.branch_set ),
    .CLK(clknet_leaf_41__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.controller_i.ctrl_fsm_cs[0]$_DFF_PN1_  (.RESET_B(net8242),
    .D(net16),
    .Q(_00006_),
    .CLK(clknet_leaf_41__06563_));
 sg13g2_tiehi \id_stage_i.controller_i.ctrl_fsm_cs[0]$_DFF_PN1__17  (.L_HI(net16));
 sg13g2_dfrbpq_1 \id_stage_i.controller_i.ctrl_fsm_cs[1]$_DFF_PN0_  (.RESET_B(net8253),
    .D(_09359_),
    .Q(_01600_),
    .CLK(clknet_leaf_40__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.controller_i.ctrl_fsm_cs[2]$_DFF_PN0_  (.RESET_B(net8241),
    .D(_09357_),
    .Q(_01601_),
    .CLK(clknet_leaf_38__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.controller_i.ctrl_fsm_cs[3]$_DFF_PN0_  (.RESET_B(net8241),
    .D(_09353_),
    .Q(_01602_),
    .CLK(clknet_leaf_38__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.controller_i.ctrl_fsm_cs[4]$_DFF_PN0_  (.RESET_B(net8241),
    .D(_07021_),
    .Q(_01603_),
    .CLK(clknet_leaf_40__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.controller_i.ctrl_fsm_cs[5]$_DFF_PN0_  (.RESET_B(net8241),
    .D(_02251_),
    .Q(_01604_),
    .CLK(clknet_leaf_38__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.controller_i.ctrl_fsm_cs[6]$_DFF_PN0_  (.RESET_B(net8257),
    .D(_09352_),
    .Q(_01605_),
    .CLK(clknet_leaf_40__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.controller_i.ctrl_fsm_cs[7]$_DFF_PN0_  (.RESET_B(net8241),
    .D(_09351_),
    .Q(\id_stage_i.controller_i.controller_run_o ),
    .CLK(clknet_leaf_40__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.controller_i.ctrl_fsm_cs[8]$_DFF_PN0_  (.RESET_B(net8241),
    .D(_09343_),
    .Q(_01606_),
    .CLK(clknet_leaf_39__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.controller_i.ctrl_fsm_cs[9]$_DFF_PN0_  (.RESET_B(net8256),
    .D(_09341_),
    .Q(\id_stage_i.controller_i.nmi_mode_d ),
    .CLK(clknet_leaf_40__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.controller_i.debug_mode_o$_DFFE_PN0P_  (.RESET_B(net8256),
    .D(_09338_),
    .Q(\cs_registers_i.debug_mode_i ),
    .CLK(clknet_leaf_40__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.controller_i.exc_req_q$_DFF_PN0_  (.RESET_B(net8257),
    .D(_09334_),
    .Q(\id_stage_i.controller_i.exc_req_q ),
    .CLK(clknet_leaf_40__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.controller_i.illegal_insn_q$_DFF_PN0_  (.RESET_B(net8257),
    .D(_09333_),
    .Q(\id_stage_i.controller_i.illegal_insn_q ),
    .CLK(clknet_leaf_40__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.controller_i.load_err_q$_DFF_PN0_  (.RESET_B(net8242),
    .D(_09327_),
    .Q(\id_stage_i.controller_i.load_err_q ),
    .CLK(clknet_leaf_42__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.controller_i.nmi_mode_o$_DFFE_PN0P_  (.RESET_B(net8253),
    .D(_09326_),
    .Q(\cs_registers_i.nmi_mode_i ),
    .CLK(clknet_leaf_40__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.controller_i.store_err_q$_DFF_PN0_  (.RESET_B(net8242),
    .D(_09319_),
    .Q(\id_stage_i.controller_i.store_err_q ),
    .CLK(clknet_leaf_42__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.id_fsm_q$_DFFE_PN0P_  (.RESET_B(net8238),
    .D(_09318_),
    .Q(\id_stage_i.id_fsm_q ),
    .CLK(clknet_leaf_41__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.imd_val_q_ex_o[0]$_DFFE_PN0P_  (.RESET_B(net8136),
    .D(_09311_),
    .Q(_01607_),
    .CLK(clknet_leaf_3__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.imd_val_q_ex_o[10]$_DFFE_PN0P_  (.RESET_B(net8136),
    .D(_09306_),
    .Q(_01608_),
    .CLK(clknet_leaf_5__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.imd_val_q_ex_o[11]$_DFFE_PN0P_  (.RESET_B(net8136),
    .D(_09301_),
    .Q(_01609_),
    .CLK(clknet_leaf_5__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.imd_val_q_ex_o[12]$_DFFE_PN0P_  (.RESET_B(net8133),
    .D(_09297_),
    .Q(_01610_),
    .CLK(clknet_leaf_5__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.imd_val_q_ex_o[13]$_DFFE_PN0P_  (.RESET_B(net8153),
    .D(_09293_),
    .Q(_01611_),
    .CLK(clknet_leaf_5__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.imd_val_q_ex_o[14]$_DFFE_PN0P_  (.RESET_B(net8153),
    .D(_09287_),
    .Q(_01612_),
    .CLK(clknet_leaf_5__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.imd_val_q_ex_o[15]$_DFFE_PN0P_  (.RESET_B(net8152),
    .D(_09283_),
    .Q(_01613_),
    .CLK(clknet_leaf_5__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.imd_val_q_ex_o[16]$_DFFE_PN0P_  (.RESET_B(net8133),
    .D(_09278_),
    .Q(_01614_),
    .CLK(clknet_leaf_5__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.imd_val_q_ex_o[17]$_DFFE_PN0P_  (.RESET_B(net8133),
    .D(_09272_),
    .Q(_01615_),
    .CLK(clknet_leaf_5__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.imd_val_q_ex_o[18]$_DFFE_PN0P_  (.RESET_B(net8136),
    .D(_09268_),
    .Q(_01616_),
    .CLK(clknet_leaf_5__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.imd_val_q_ex_o[19]$_DFFE_PN0P_  (.RESET_B(net8151),
    .D(_09264_),
    .Q(_01617_),
    .CLK(clknet_leaf_6__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.imd_val_q_ex_o[1]$_DFFE_PN0P_  (.RESET_B(net8133),
    .D(_09258_),
    .Q(_01618_),
    .CLK(clknet_leaf_5__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.imd_val_q_ex_o[20]$_DFFE_PN0P_  (.RESET_B(net8145),
    .D(_09253_),
    .Q(_01619_),
    .CLK(clknet_leaf_7__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.imd_val_q_ex_o[21]$_DFFE_PN0P_  (.RESET_B(net8145),
    .D(_09248_),
    .Q(_01620_),
    .CLK(clknet_leaf_7__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.imd_val_q_ex_o[22]$_DFFE_PN0P_  (.RESET_B(net8152),
    .D(_09242_),
    .Q(_01621_),
    .CLK(clknet_leaf_6__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.imd_val_q_ex_o[23]$_DFFE_PN0P_  (.RESET_B(net8145),
    .D(_09238_),
    .Q(_01622_),
    .CLK(clknet_leaf_7__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.imd_val_q_ex_o[24]$_DFFE_PN0P_  (.RESET_B(net8152),
    .D(_09233_),
    .Q(_01623_),
    .CLK(clknet_leaf_6__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.imd_val_q_ex_o[25]$_DFFE_PN0P_  (.RESET_B(net8154),
    .D(_09228_),
    .Q(_01624_),
    .CLK(clknet_leaf_7__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.imd_val_q_ex_o[26]$_DFFE_PN0P_  (.RESET_B(net8151),
    .D(_09224_),
    .Q(_01625_),
    .CLK(clknet_leaf_6__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.imd_val_q_ex_o[27]$_DFFE_PN0P_  (.RESET_B(net8153),
    .D(_09219_),
    .Q(_01626_),
    .CLK(clknet_leaf_5__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.imd_val_q_ex_o[28]$_DFFE_PN0P_  (.RESET_B(net8153),
    .D(_09215_),
    .Q(_01627_),
    .CLK(clknet_leaf_5__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.imd_val_q_ex_o[29]$_DFFE_PN0P_  (.RESET_B(net8146),
    .D(_09211_),
    .Q(_01628_),
    .CLK(clknet_leaf_7__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.imd_val_q_ex_o[2]$_DFFE_PN0P_  (.RESET_B(net8136),
    .D(_09207_),
    .Q(_01629_),
    .CLK(clknet_leaf_2__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.imd_val_q_ex_o[30]$_DFFE_PN0P_  (.RESET_B(net8145),
    .D(_09203_),
    .Q(_01630_),
    .CLK(clknet_leaf_7__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.imd_val_q_ex_o[31]$_DFFE_PN0P_  (.RESET_B(net8145),
    .D(_09199_),
    .Q(_01631_),
    .CLK(clknet_leaf_7__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.imd_val_q_ex_o[34]$_DFFE_PN0P_  (.RESET_B(net8161),
    .D(_09196_),
    .Q(_01632_),
    .CLK(clknet_leaf_8__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.imd_val_q_ex_o[35]$_DFFE_PN0P_  (.RESET_B(net8158),
    .D(_09141_),
    .Q(_01633_),
    .CLK(clknet_leaf_8__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.imd_val_q_ex_o[36]$_DFFE_PN0P_  (.RESET_B(net8158),
    .D(_09127_),
    .Q(_01634_),
    .CLK(clknet_leaf_8__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.imd_val_q_ex_o[37]$_DFFE_PN0P_  (.RESET_B(net8158),
    .D(_09117_),
    .Q(_01635_),
    .CLK(clknet_leaf_8__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.imd_val_q_ex_o[38]$_DFFE_PN0P_  (.RESET_B(net8158),
    .D(_09107_),
    .Q(_01636_),
    .CLK(clknet_leaf_8__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.imd_val_q_ex_o[39]$_DFFE_PN0P_  (.RESET_B(net8159),
    .D(_09096_),
    .Q(_01637_),
    .CLK(clknet_leaf_8__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.imd_val_q_ex_o[3]$_DFFE_PN0P_  (.RESET_B(net8136),
    .D(_09086_),
    .Q(_01638_),
    .CLK(clknet_leaf_2__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.imd_val_q_ex_o[40]$_DFFE_PN0P_  (.RESET_B(net8159),
    .D(_09082_),
    .Q(_01639_),
    .CLK(clknet_leaf_8__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.imd_val_q_ex_o[41]$_DFFE_PN0P_  (.RESET_B(net8159),
    .D(_09071_),
    .Q(_01640_),
    .CLK(clknet_leaf_8__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.imd_val_q_ex_o[42]$_DFFE_PN0P_  (.RESET_B(net8161),
    .D(_09058_),
    .Q(_01641_),
    .CLK(clknet_leaf_8__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.imd_val_q_ex_o[43]$_DFFE_PN0P_  (.RESET_B(net8158),
    .D(_09048_),
    .Q(_01642_),
    .CLK(clknet_leaf_8__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.imd_val_q_ex_o[44]$_DFFE_PN0P_  (.RESET_B(net8145),
    .D(_09036_),
    .Q(_01643_),
    .CLK(clknet_leaf_7__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.imd_val_q_ex_o[45]$_DFFE_PN0P_  (.RESET_B(net8161),
    .D(_09022_),
    .Q(_01644_),
    .CLK(clknet_leaf_7__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.imd_val_q_ex_o[46]$_DFFE_PN0P_  (.RESET_B(net8158),
    .D(_09010_),
    .Q(_01645_),
    .CLK(clknet_leaf_7__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.imd_val_q_ex_o[47]$_DFFE_PN0P_  (.RESET_B(net8159),
    .D(_08996_),
    .Q(_01646_),
    .CLK(clknet_leaf_8__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.imd_val_q_ex_o[48]$_DFFE_PN0P_  (.RESET_B(net8160),
    .D(_08984_),
    .Q(_01647_),
    .CLK(clknet_leaf_8__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.imd_val_q_ex_o[49]$_DFFE_PN0P_  (.RESET_B(net8159),
    .D(_08968_),
    .Q(_01648_),
    .CLK(clknet_leaf_8__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.imd_val_q_ex_o[4]$_DFFE_PN0P_  (.RESET_B(net8145),
    .D(_08954_),
    .Q(_01649_),
    .CLK(clknet_leaf_7__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.imd_val_q_ex_o[50]$_DFFE_PN0P_  (.RESET_B(net8160),
    .D(_08950_),
    .Q(_01650_),
    .CLK(clknet_leaf_8__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.imd_val_q_ex_o[51]$_DFFE_PN0P_  (.RESET_B(net8159),
    .D(_08935_),
    .Q(_01651_),
    .CLK(clknet_leaf_9__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.imd_val_q_ex_o[52]$_DFFE_PN0P_  (.RESET_B(net8160),
    .D(_08925_),
    .Q(_01652_),
    .CLK(clknet_leaf_8__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.imd_val_q_ex_o[53]$_DFFE_PN0P_  (.RESET_B(net8189),
    .D(_08913_),
    .Q(_01653_),
    .CLK(clknet_leaf_9__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.imd_val_q_ex_o[54]$_DFFE_PN0P_  (.RESET_B(net8188),
    .D(_08900_),
    .Q(_01654_),
    .CLK(clknet_leaf_11__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.imd_val_q_ex_o[55]$_DFFE_PN0P_  (.RESET_B(net8188),
    .D(_08886_),
    .Q(_01655_),
    .CLK(clknet_leaf_11__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.imd_val_q_ex_o[56]$_DFFE_PN0P_  (.RESET_B(net8171),
    .D(_08875_),
    .Q(_01656_),
    .CLK(clknet_leaf_10__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.imd_val_q_ex_o[57]$_DFFE_PN0P_  (.RESET_B(net8189),
    .D(_08862_),
    .Q(_01657_),
    .CLK(clknet_leaf_11__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.imd_val_q_ex_o[58]$_DFFE_PN0P_  (.RESET_B(net8165),
    .D(_08848_),
    .Q(_01658_),
    .CLK(clknet_leaf_9__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.imd_val_q_ex_o[59]$_DFFE_PN0P_  (.RESET_B(net8189),
    .D(_08833_),
    .Q(_01659_),
    .CLK(clknet_leaf_9__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.imd_val_q_ex_o[5]$_DFFE_PN0P_  (.RESET_B(net8152),
    .D(_08821_),
    .Q(_01660_),
    .CLK(clknet_leaf_6__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.imd_val_q_ex_o[60]$_DFFE_PN0P_  (.RESET_B(net8165),
    .D(_08816_),
    .Q(_01661_),
    .CLK(clknet_leaf_9__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.imd_val_q_ex_o[61]$_DFFE_PN0P_  (.RESET_B(net8189),
    .D(_08803_),
    .Q(_01662_),
    .CLK(clknet_leaf_9__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.imd_val_q_ex_o[62]$_DFFE_PN0P_  (.RESET_B(net8160),
    .D(_08788_),
    .Q(_01663_),
    .CLK(clknet_leaf_8__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.imd_val_q_ex_o[63]$_DFFE_PN0P_  (.RESET_B(net8165),
    .D(_08770_),
    .Q(_01664_),
    .CLK(clknet_leaf_9__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.imd_val_q_ex_o[64]$_DFFE_PN0P_  (.RESET_B(net8206),
    .D(_08756_),
    .Q(_01665_),
    .CLK(clknet_leaf_9__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.imd_val_q_ex_o[65]$_DFFE_PN0P_  (.RESET_B(net8160),
    .D(_08741_),
    .Q(_01666_),
    .CLK(clknet_leaf_8__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.imd_val_q_ex_o[66]$_DFFE_PN0P_  (.RESET_B(net8160),
    .D(_08719_),
    .Q(_01667_),
    .CLK(clknet_leaf_8__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.imd_val_q_ex_o[67]$_DFFE_PN0P_  (.RESET_B(net8206),
    .D(_08713_),
    .Q(_01668_),
    .CLK(clknet_leaf_9__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.imd_val_q_ex_o[6]$_DFFE_PN0P_  (.RESET_B(net8154),
    .D(_08684_),
    .Q(_01669_),
    .CLK(clknet_leaf_7__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.imd_val_q_ex_o[7]$_DFFE_PN0P_  (.RESET_B(net8151),
    .D(_08679_),
    .Q(_01670_),
    .CLK(clknet_leaf_6__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.imd_val_q_ex_o[8]$_DFFE_PN0P_  (.RESET_B(net8133),
    .D(_08675_),
    .Q(_01671_),
    .CLK(clknet_leaf_5__06563_));
 sg13g2_dfrbpq_1 \id_stage_i.imd_val_q_ex_o[9]$_DFFE_PN0P_  (.RESET_B(net8136),
    .D(_08670_),
    .Q(_01672_),
    .CLK(clknet_leaf_5__06563_));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[0]$_DFF_PN0_  (.RESET_B(net8239),
    .D(_08656_),
    .Q(_01673_),
    .CLK(clknet_leaf_44__06563_));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[1]$_DFF_PN0_  (.RESET_B(net8239),
    .D(_08651_),
    .Q(_01674_),
    .CLK(clknet_leaf_44__06563_));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_q$_DFF_PN0_  (.RESET_B(net8239),
    .D(_08647_),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_q ),
    .CLK(clknet_leaf_44__06563_));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[10]$_DFFE_PP_  (.RESET_B(net17),
    .D(_08646_),
    .Q(_01675_),
    .CLK(clknet_leaf_46__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[10]$_DFFE_PP__18  (.L_HI(net17));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[11]$_DFFE_PP_  (.RESET_B(net18),
    .D(_08644_),
    .Q(_01676_),
    .CLK(clknet_leaf_37__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[11]$_DFFE_PP__19  (.L_HI(net18));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[12]$_DFFE_PP_  (.RESET_B(net19),
    .D(_08642_),
    .Q(_01677_),
    .CLK(clknet_leaf_46__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[12]$_DFFE_PP__20  (.L_HI(net19));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[13]$_DFFE_PP_  (.RESET_B(net20),
    .D(_08640_),
    .Q(_01678_),
    .CLK(clknet_leaf_46__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[13]$_DFFE_PP__21  (.L_HI(net20));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[14]$_DFFE_PP_  (.RESET_B(net21),
    .D(_08637_),
    .Q(_01679_),
    .CLK(clknet_leaf_45__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[14]$_DFFE_PP__22  (.L_HI(net21));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[15]$_DFFE_PP_  (.RESET_B(net22),
    .D(_08635_),
    .Q(_01680_),
    .CLK(clknet_leaf_45__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[15]$_DFFE_PP__23  (.L_HI(net22));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[16]$_DFFE_PP_  (.RESET_B(net23),
    .D(_08633_),
    .Q(_01681_),
    .CLK(clknet_leaf_46__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[16]$_DFFE_PP__24  (.L_HI(net23));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[17]$_DFFE_PP_  (.RESET_B(net24),
    .D(_08632_),
    .Q(_01682_),
    .CLK(clknet_leaf_46__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[17]$_DFFE_PP__25  (.L_HI(net24));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[18]$_DFFE_PP_  (.RESET_B(net25),
    .D(_08628_),
    .Q(_01683_),
    .CLK(clknet_leaf_46__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[18]$_DFFE_PP__26  (.L_HI(net25));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[19]$_DFFE_PP_  (.RESET_B(net26),
    .D(_08626_),
    .Q(_01684_),
    .CLK(clknet_leaf_46__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[19]$_DFFE_PP__27  (.L_HI(net26));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[20]$_DFFE_PP_  (.RESET_B(net27),
    .D(_08624_),
    .Q(_01685_),
    .CLK(clknet_leaf_46__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[20]$_DFFE_PP__28  (.L_HI(net27));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[21]$_DFFE_PP_  (.RESET_B(net28),
    .D(_08621_),
    .Q(_01686_),
    .CLK(clknet_leaf_37__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[21]$_DFFE_PP__29  (.L_HI(net28));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[22]$_DFFE_PP_  (.RESET_B(net29),
    .D(_08620_),
    .Q(_01687_),
    .CLK(clknet_leaf_37__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[22]$_DFFE_PP__30  (.L_HI(net29));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[23]$_DFFE_PP_  (.RESET_B(net30),
    .D(_08619_),
    .Q(_01688_),
    .CLK(clknet_leaf_37__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[23]$_DFFE_PP__31  (.L_HI(net30));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[24]$_DFFE_PP_  (.RESET_B(net31),
    .D(_08617_),
    .Q(_01689_),
    .CLK(clknet_leaf_37__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[24]$_DFFE_PP__32  (.L_HI(net31));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[25]$_DFFE_PP_  (.RESET_B(net32),
    .D(_08615_),
    .Q(_01690_),
    .CLK(clknet_leaf_37__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[25]$_DFFE_PP__33  (.L_HI(net32));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[26]$_DFFE_PP_  (.RESET_B(net33),
    .D(_08613_),
    .Q(_01691_),
    .CLK(clknet_leaf_37__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[26]$_DFFE_PP__34  (.L_HI(net33));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[27]$_DFFE_PP_  (.RESET_B(net34),
    .D(_08612_),
    .Q(_01692_),
    .CLK(clknet_leaf_36__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[27]$_DFFE_PP__35  (.L_HI(net34));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[28]$_DFFE_PP_  (.RESET_B(net35),
    .D(_08610_),
    .Q(_01693_),
    .CLK(clknet_leaf_36__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[28]$_DFFE_PP__36  (.L_HI(net35));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[29]$_DFFE_PP_  (.RESET_B(net36),
    .D(_08609_),
    .Q(_01694_),
    .CLK(clknet_leaf_36__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[29]$_DFFE_PP__37  (.L_HI(net36));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[2]$_DFFE_PP_  (.RESET_B(net37),
    .D(_08608_),
    .Q(_01695_),
    .CLK(clknet_leaf_45__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[2]$_DFFE_PP__38  (.L_HI(net37));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[30]$_DFFE_PP_  (.RESET_B(net38),
    .D(_08607_),
    .Q(_01696_),
    .CLK(clknet_leaf_36__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[30]$_DFFE_PP__39  (.L_HI(net38));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[31]$_DFFE_PP_  (.RESET_B(net39),
    .D(_08603_),
    .Q(_01697_),
    .CLK(clknet_leaf_47__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[31]$_DFFE_PP__40  (.L_HI(net39));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[3]$_DFFE_PP_  (.RESET_B(net40),
    .D(_08565_),
    .Q(_01698_),
    .CLK(clknet_leaf_44__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[3]$_DFFE_PP__41  (.L_HI(net40));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[4]$_DFFE_PP_  (.RESET_B(net41),
    .D(_08564_),
    .Q(_01699_),
    .CLK(clknet_leaf_44__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[4]$_DFFE_PP__42  (.L_HI(net41));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[5]$_DFFE_PP_  (.RESET_B(net42),
    .D(_08562_),
    .Q(_01700_),
    .CLK(clknet_leaf_45__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[5]$_DFFE_PP__43  (.L_HI(net42));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[6]$_DFFE_PP_  (.RESET_B(net43),
    .D(_08560_),
    .Q(_01701_),
    .CLK(clknet_leaf_45__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[6]$_DFFE_PP__44  (.L_HI(net43));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[7]$_DFFE_PP_  (.RESET_B(net44),
    .D(_08559_),
    .Q(_01702_),
    .CLK(clknet_leaf_45__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[7]$_DFFE_PP__45  (.L_HI(net44));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[8]$_DFFE_PP_  (.RESET_B(net45),
    .D(_08558_),
    .Q(_01703_),
    .CLK(clknet_leaf_45__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[8]$_DFFE_PP__46  (.L_HI(net45));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[9]$_DFFE_PP_  (.RESET_B(net46),
    .D(_08556_),
    .Q(_01704_),
    .CLK(clknet_leaf_46__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[9]$_DFFE_PP__47  (.L_HI(net46));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[0]$_DFFE_PP_  (.RESET_B(net47),
    .D(_08547_),
    .Q(_01705_),
    .CLK(clknet_leaf_47__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[0]$_DFFE_PP__48  (.L_HI(net47));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[1]$_DFFE_PP_  (.RESET_B(net48),
    .D(_08544_),
    .Q(_01706_),
    .CLK(clknet_leaf_47__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[1]$_DFFE_PP__49  (.L_HI(net48));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[2]$_DFFE_PP_  (.RESET_B(net49),
    .D(_08539_),
    .Q(_01707_),
    .CLK(clknet_leaf_47__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[2]$_DFFE_PP__50  (.L_HI(net49));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[10]$_DFFE_PP_  (.RESET_B(net50),
    .D(_08537_),
    .Q(_01708_),
    .CLK(clknet_leaf_38__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[10]$_DFFE_PP__51  (.L_HI(net50));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[11]$_DFFE_PP_  (.RESET_B(net51),
    .D(_08535_),
    .Q(_01709_),
    .CLK(clknet_leaf_37__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[11]$_DFFE_PP__52  (.L_HI(net51));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[12]$_DFFE_PP_  (.RESET_B(net52),
    .D(_08532_),
    .Q(_01710_),
    .CLK(clknet_leaf_45__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[12]$_DFFE_PP__53  (.L_HI(net52));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[13]$_DFFE_PP_  (.RESET_B(net53),
    .D(_08528_),
    .Q(_01711_),
    .CLK(clknet_leaf_38__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[13]$_DFFE_PP__54  (.L_HI(net53));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[14]$_DFFE_PP_  (.RESET_B(net54),
    .D(_08521_),
    .Q(_01712_),
    .CLK(clknet_leaf_38__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[14]$_DFFE_PP__55  (.L_HI(net54));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[15]$_DFFE_PP_  (.RESET_B(net55),
    .D(_08518_),
    .Q(_01713_),
    .CLK(clknet_leaf_38__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[15]$_DFFE_PP__56  (.L_HI(net55));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[16]$_DFFE_PP_  (.RESET_B(net56),
    .D(_08514_),
    .Q(_01714_),
    .CLK(clknet_leaf_38__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[16]$_DFFE_PP__57  (.L_HI(net56));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[17]$_DFFE_PP_  (.RESET_B(net57),
    .D(_08509_),
    .Q(_01715_),
    .CLK(clknet_leaf_38__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[17]$_DFFE_PP__58  (.L_HI(net57));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[18]$_DFFE_PP_  (.RESET_B(net58),
    .D(_08504_),
    .Q(_01716_),
    .CLK(clknet_leaf_36__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[18]$_DFFE_PP__59  (.L_HI(net58));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[19]$_DFFE_PP_  (.RESET_B(net59),
    .D(_08501_),
    .Q(_01717_),
    .CLK(clknet_leaf_37__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[19]$_DFFE_PP__60  (.L_HI(net59));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[1]$_DFFE_PP_  (.RESET_B(net60),
    .D(_08496_),
    .Q(_01718_),
    .CLK(clknet_leaf_45__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[1]$_DFFE_PP__61  (.L_HI(net60));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[20]$_DFFE_PP_  (.RESET_B(net61),
    .D(_08491_),
    .Q(_01719_),
    .CLK(clknet_leaf_36__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[20]$_DFFE_PP__62  (.L_HI(net61));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[21]$_DFFE_PP_  (.RESET_B(net62),
    .D(_08487_),
    .Q(_01720_),
    .CLK(clknet_leaf_38__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[21]$_DFFE_PP__63  (.L_HI(net62));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[22]$_DFFE_PP_  (.RESET_B(net63),
    .D(_08483_),
    .Q(_01721_),
    .CLK(clknet_leaf_37__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[22]$_DFFE_PP__64  (.L_HI(net63));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[23]$_DFFE_PP_  (.RESET_B(net64),
    .D(_08478_),
    .Q(_01722_),
    .CLK(clknet_leaf_37__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[23]$_DFFE_PP__65  (.L_HI(net64));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[24]$_DFFE_PP_  (.RESET_B(net65),
    .D(_08474_),
    .Q(_01723_),
    .CLK(clknet_leaf_36__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[24]$_DFFE_PP__66  (.L_HI(net65));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[25]$_DFFE_PP_  (.RESET_B(net66),
    .D(_08471_),
    .Q(_01724_),
    .CLK(clknet_leaf_36__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[25]$_DFFE_PP__67  (.L_HI(net66));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[26]$_DFFE_PP_  (.RESET_B(net67),
    .D(_08466_),
    .Q(_01725_),
    .CLK(clknet_leaf_36__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[26]$_DFFE_PP__68  (.L_HI(net67));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[27]$_DFFE_PP_  (.RESET_B(net68),
    .D(_08463_),
    .Q(_01726_),
    .CLK(clknet_leaf_36__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[27]$_DFFE_PP__69  (.L_HI(net68));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[28]$_DFFE_PP_  (.RESET_B(net69),
    .D(_08458_),
    .Q(_01727_),
    .CLK(clknet_leaf_36__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[28]$_DFFE_PP__70  (.L_HI(net69));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[29]$_DFFE_PP_  (.RESET_B(net70),
    .D(_08453_),
    .Q(_01728_),
    .CLK(clknet_leaf_36__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[29]$_DFFE_PP__71  (.L_HI(net70));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[2]$_DFFE_PP_  (.RESET_B(net71),
    .D(_08449_),
    .Q(_01729_),
    .CLK(clknet_leaf_45__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[2]$_DFFE_PP__72  (.L_HI(net71));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[30]$_DFFE_PP_  (.RESET_B(net72),
    .D(_08445_),
    .Q(_01730_),
    .CLK(clknet_leaf_36__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[30]$_DFFE_PP__73  (.L_HI(net72));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[31]$_DFFE_PP_  (.RESET_B(net73),
    .D(_08441_),
    .Q(_01731_),
    .CLK(clknet_leaf_36__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[31]$_DFFE_PP__74  (.L_HI(net73));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[3]$_DFFE_PP_  (.RESET_B(net74),
    .D(_08422_),
    .Q(_01732_),
    .CLK(clknet_leaf_45__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[3]$_DFFE_PP__75  (.L_HI(net74));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[4]$_DFFE_PP_  (.RESET_B(net75),
    .D(_08419_),
    .Q(_01733_),
    .CLK(clknet_leaf_45__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[4]$_DFFE_PP__76  (.L_HI(net75));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[5]$_DFFE_PP_  (.RESET_B(net76),
    .D(_08413_),
    .Q(_01734_),
    .CLK(clknet_leaf_38__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[5]$_DFFE_PP__77  (.L_HI(net76));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[6]$_DFFE_PP_  (.RESET_B(net77),
    .D(_08408_),
    .Q(_01735_),
    .CLK(clknet_leaf_38__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[6]$_DFFE_PP__78  (.L_HI(net77));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[7]$_DFFE_PP_  (.RESET_B(net78),
    .D(_08406_),
    .Q(_01736_),
    .CLK(clknet_leaf_38__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[7]$_DFFE_PP__79  (.L_HI(net78));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[8]$_DFFE_PP_  (.RESET_B(net79),
    .D(_08404_),
    .Q(_01737_),
    .CLK(clknet_leaf_45__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[8]$_DFFE_PP__80  (.L_HI(net79));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[9]$_DFFE_PP_  (.RESET_B(net80),
    .D(_08399_),
    .Q(_01738_),
    .CLK(clknet_leaf_45__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[9]$_DFFE_PP__81  (.L_HI(net80));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[0]$_DFFE_PP_  (.RESET_B(net81),
    .D(_08390_),
    .Q(_01739_),
    .CLK(clknet_leaf_47__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[0]$_DFFE_PP__82  (.L_HI(net81));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[10]$_DFFE_PP_  (.RESET_B(net82),
    .D(_08386_),
    .Q(_01740_),
    .CLK(clknet_leaf_49__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[10]$_DFFE_PP__83  (.L_HI(net82));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[11]$_DFFE_PP_  (.RESET_B(net83),
    .D(_08382_),
    .Q(_01741_),
    .CLK(clknet_leaf_49__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[11]$_DFFE_PP__84  (.L_HI(net83));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[12]$_DFFE_PP_  (.RESET_B(net84),
    .D(_08380_),
    .Q(_01742_),
    .CLK(clknet_leaf_49__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[12]$_DFFE_PP__85  (.L_HI(net84));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[13]$_DFFE_PP_  (.RESET_B(net85),
    .D(_08378_),
    .Q(_01743_),
    .CLK(clknet_leaf_48__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[13]$_DFFE_PP__86  (.L_HI(net85));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[14]$_DFFE_PP_  (.RESET_B(net86),
    .D(_08375_),
    .Q(_01744_),
    .CLK(clknet_leaf_48__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[14]$_DFFE_PP__87  (.L_HI(net86));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[15]$_DFFE_PP_  (.RESET_B(net87),
    .D(_08374_),
    .Q(_01745_),
    .CLK(clknet_leaf_49__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[15]$_DFFE_PP__88  (.L_HI(net87));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[16]$_DFFE_PP_  (.RESET_B(net88),
    .D(_08372_),
    .Q(_01746_),
    .CLK(clknet_leaf_47__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[16]$_DFFE_PP__89  (.L_HI(net88));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[17]$_DFFE_PP_  (.RESET_B(net89),
    .D(_08368_),
    .Q(_01747_),
    .CLK(clknet_leaf_47__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[17]$_DFFE_PP__90  (.L_HI(net89));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[18]$_DFFE_PP_  (.RESET_B(net90),
    .D(_08364_),
    .Q(_01748_),
    .CLK(clknet_leaf_50__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[18]$_DFFE_PP__91  (.L_HI(net90));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[19]$_DFFE_PP_  (.RESET_B(net91),
    .D(_08360_),
    .Q(_01749_),
    .CLK(clknet_leaf_49__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[19]$_DFFE_PP__92  (.L_HI(net91));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[1]$_DFFE_PP_  (.RESET_B(net92),
    .D(_08356_),
    .Q(_01750_),
    .CLK(clknet_leaf_48__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[1]$_DFFE_PP__93  (.L_HI(net92));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[20]$_DFFE_PP_  (.RESET_B(net93),
    .D(_08355_),
    .Q(_01751_),
    .CLK(clknet_leaf_50__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[20]$_DFFE_PP__94  (.L_HI(net93));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[21]$_DFFE_PP_  (.RESET_B(net94),
    .D(_08351_),
    .Q(_01752_),
    .CLK(clknet_leaf_0__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[21]$_DFFE_PP__95  (.L_HI(net94));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[22]$_DFFE_PP_  (.RESET_B(net95),
    .D(_08346_),
    .Q(_01753_),
    .CLK(clknet_leaf_0__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[22]$_DFFE_PP__96  (.L_HI(net95));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[23]$_DFFE_PP_  (.RESET_B(net96),
    .D(_08342_),
    .Q(_01754_),
    .CLK(clknet_leaf_0__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[23]$_DFFE_PP__97  (.L_HI(net96));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[24]$_DFFE_PP_  (.RESET_B(net97),
    .D(_08338_),
    .Q(_01755_),
    .CLK(clknet_leaf_0__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[24]$_DFFE_PP__98  (.L_HI(net97));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[25]$_DFFE_PP_  (.RESET_B(net98),
    .D(_08333_),
    .Q(_01756_),
    .CLK(clknet_leaf_48__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[25]$_DFFE_PP__99  (.L_HI(net98));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[26]$_DFFE_PP_  (.RESET_B(net99),
    .D(_08329_),
    .Q(_01757_),
    .CLK(clknet_leaf_50__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[26]$_DFFE_PP__100  (.L_HI(net99));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[27]$_DFFE_PP_  (.RESET_B(net100),
    .D(_08324_),
    .Q(_01758_),
    .CLK(clknet_leaf_49__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[27]$_DFFE_PP__101  (.L_HI(net100));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[28]$_DFFE_PP_  (.RESET_B(net101),
    .D(_08319_),
    .Q(_01759_),
    .CLK(clknet_leaf_49__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[28]$_DFFE_PP__102  (.L_HI(net101));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[29]$_DFFE_PP_  (.RESET_B(net102),
    .D(_08314_),
    .Q(_01760_),
    .CLK(clknet_leaf_48__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[29]$_DFFE_PP__103  (.L_HI(net102));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[2]$_DFFE_PP_  (.RESET_B(net103),
    .D(_08308_),
    .Q(_01761_),
    .CLK(clknet_leaf_0__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[2]$_DFFE_PP__104  (.L_HI(net103));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[30]$_DFFE_PP_  (.RESET_B(net104),
    .D(_08304_),
    .Q(_01762_),
    .CLK(clknet_leaf_49__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[30]$_DFFE_PP__105  (.L_HI(net104));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[31]$_DFFE_PP_  (.RESET_B(net105),
    .D(_08299_),
    .Q(_01763_),
    .CLK(clknet_leaf_49__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[31]$_DFFE_PP__106  (.L_HI(net105));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[32]$_DFFE_PP_  (.RESET_B(net106),
    .D(_08294_),
    .Q(_01764_),
    .CLK(clknet_leaf_47__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[32]$_DFFE_PP__107  (.L_HI(net106));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[33]$_DFFE_PP_  (.RESET_B(net107),
    .D(_08287_),
    .Q(_01765_),
    .CLK(clknet_leaf_48__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[33]$_DFFE_PP__108  (.L_HI(net107));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[34]$_DFFE_PP_  (.RESET_B(net108),
    .D(_08281_),
    .Q(_01766_),
    .CLK(clknet_leaf_51__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[34]$_DFFE_PP__109  (.L_HI(net108));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[35]$_DFFE_PP_  (.RESET_B(net109),
    .D(_08276_),
    .Q(_01767_),
    .CLK(clknet_leaf_50__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[35]$_DFFE_PP__110  (.L_HI(net109));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[36]$_DFFE_PP_  (.RESET_B(net110),
    .D(_08272_),
    .Q(_01768_),
    .CLK(clknet_leaf_50__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[36]$_DFFE_PP__111  (.L_HI(net110));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[37]$_DFFE_PP_  (.RESET_B(net111),
    .D(_08268_),
    .Q(_01769_),
    .CLK(clknet_leaf_51__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[37]$_DFFE_PP__112  (.L_HI(net111));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[38]$_DFFE_PP_  (.RESET_B(net112),
    .D(_08264_),
    .Q(_01770_),
    .CLK(clknet_leaf_0__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[38]$_DFFE_PP__113  (.L_HI(net112));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[39]$_DFFE_PP_  (.RESET_B(net113),
    .D(_08260_),
    .Q(_01771_),
    .CLK(clknet_leaf_0__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[39]$_DFFE_PP__114  (.L_HI(net113));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[3]$_DFFE_PP_  (.RESET_B(net114),
    .D(_08256_),
    .Q(_01772_),
    .CLK(clknet_leaf_49__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[3]$_DFFE_PP__115  (.L_HI(net114));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[40]$_DFFE_PP_  (.RESET_B(net115),
    .D(_08253_),
    .Q(_01773_),
    .CLK(clknet_leaf_0__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[40]$_DFFE_PP__116  (.L_HI(net115));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[41]$_DFFE_PP_  (.RESET_B(net116),
    .D(_08246_),
    .Q(_01774_),
    .CLK(clknet_leaf_48__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[41]$_DFFE_PP__117  (.L_HI(net116));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[42]$_DFFE_PP_  (.RESET_B(net117),
    .D(_08241_),
    .Q(_01775_),
    .CLK(clknet_leaf_50__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[42]$_DFFE_PP__118  (.L_HI(net117));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[43]$_DFFE_PP_  (.RESET_B(net118),
    .D(_08235_),
    .Q(_01776_),
    .CLK(clknet_leaf_50__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[43]$_DFFE_PP__119  (.L_HI(net118));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[44]$_DFFE_PP_  (.RESET_B(net119),
    .D(_08230_),
    .Q(_01777_),
    .CLK(clknet_leaf_49__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[44]$_DFFE_PP__120  (.L_HI(net119));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[45]$_DFFE_PP_  (.RESET_B(net120),
    .D(_08224_),
    .Q(_01778_),
    .CLK(clknet_leaf_48__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[45]$_DFFE_PP__121  (.L_HI(net120));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[46]$_DFFE_PP_  (.RESET_B(net121),
    .D(_08219_),
    .Q(_01779_),
    .CLK(clknet_leaf_49__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[46]$_DFFE_PP__122  (.L_HI(net121));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[47]$_DFFE_PP_  (.RESET_B(net122),
    .D(_08215_),
    .Q(_01780_),
    .CLK(clknet_leaf_50__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[47]$_DFFE_PP__123  (.L_HI(net122));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[48]$_DFFE_PP_  (.RESET_B(net123),
    .D(_08210_),
    .Q(_01781_),
    .CLK(clknet_leaf_47__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[48]$_DFFE_PP__124  (.L_HI(net123));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[49]$_DFFE_PP_  (.RESET_B(net124),
    .D(_08204_),
    .Q(_01782_),
    .CLK(clknet_leaf_48__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[49]$_DFFE_PP__125  (.L_HI(net124));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[4]$_DFFE_PP_  (.RESET_B(net125),
    .D(_08199_),
    .Q(_01783_),
    .CLK(clknet_leaf_0__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[4]$_DFFE_PP__126  (.L_HI(net125));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[50]$_DFFE_PP_  (.RESET_B(net126),
    .D(_08197_),
    .Q(_01784_),
    .CLK(clknet_leaf_51__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[50]$_DFFE_PP__127  (.L_HI(net126));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[51]$_DFFE_PP_  (.RESET_B(net127),
    .D(_08192_),
    .Q(_01785_),
    .CLK(clknet_leaf_49__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[51]$_DFFE_PP__128  (.L_HI(net127));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[52]$_DFFE_PP_  (.RESET_B(net128),
    .D(_08188_),
    .Q(_01786_),
    .CLK(clknet_leaf_50__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[52]$_DFFE_PP__129  (.L_HI(net128));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[53]$_DFFE_PP_  (.RESET_B(net129),
    .D(_08183_),
    .Q(_01787_),
    .CLK(clknet_leaf_51__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[53]$_DFFE_PP__130  (.L_HI(net129));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[54]$_DFFE_PP_  (.RESET_B(net130),
    .D(_08178_),
    .Q(_01788_),
    .CLK(clknet_leaf_51__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[54]$_DFFE_PP__131  (.L_HI(net130));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[55]$_DFFE_PP_  (.RESET_B(net131),
    .D(_08172_),
    .Q(_01789_),
    .CLK(clknet_leaf_0__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[55]$_DFFE_PP__132  (.L_HI(net131));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[56]$_DFFE_PP_  (.RESET_B(net132),
    .D(_08167_),
    .Q(_01790_),
    .CLK(clknet_leaf_51__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[56]$_DFFE_PP__133  (.L_HI(net132));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[57]$_DFFE_PP_  (.RESET_B(net133),
    .D(_08162_),
    .Q(_01791_),
    .CLK(clknet_leaf_48__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[57]$_DFFE_PP__134  (.L_HI(net133));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[58]$_DFFE_PP_  (.RESET_B(net134),
    .D(_08156_),
    .Q(_01792_),
    .CLK(clknet_leaf_51__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[58]$_DFFE_PP__135  (.L_HI(net134));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[59]$_DFFE_PP_  (.RESET_B(net135),
    .D(_08150_),
    .Q(_01793_),
    .CLK(clknet_leaf_50__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[59]$_DFFE_PP__136  (.L_HI(net135));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[5]$_DFFE_PP_  (.RESET_B(net136),
    .D(_08146_),
    .Q(_01794_),
    .CLK(clknet_leaf_51__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[5]$_DFFE_PP__137  (.L_HI(net136));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[60]$_DFFE_PP_  (.RESET_B(net137),
    .D(_08144_),
    .Q(_01795_),
    .CLK(clknet_leaf_49__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[60]$_DFFE_PP__138  (.L_HI(net137));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[61]$_DFFE_PP_  (.RESET_B(net138),
    .D(_08139_),
    .Q(_01796_),
    .CLK(clknet_leaf_48__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[61]$_DFFE_PP__139  (.L_HI(net138));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[62]$_DFFE_PP_  (.RESET_B(net139),
    .D(_08134_),
    .Q(_01797_),
    .CLK(clknet_leaf_49__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[62]$_DFFE_PP__140  (.L_HI(net139));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[63]$_DFFE_PP_  (.RESET_B(net140),
    .D(_08128_),
    .Q(_01798_),
    .CLK(clknet_leaf_50__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[63]$_DFFE_PP__141  (.L_HI(net140));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[64]$_DFFE_PP_  (.RESET_B(net141),
    .D(_08120_),
    .Q(_01799_),
    .CLK(clknet_leaf_47__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[64]$_DFFE_PP__142  (.L_HI(net141));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[65]$_DFFE_PP_  (.RESET_B(net142),
    .D(_08119_),
    .Q(_01800_),
    .CLK(clknet_leaf_48__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[65]$_DFFE_PP__143  (.L_HI(net142));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[66]$_DFFE_PP_  (.RESET_B(net143),
    .D(_08118_),
    .Q(_01801_),
    .CLK(clknet_leaf_51__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[66]$_DFFE_PP__144  (.L_HI(net143));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[67]$_DFFE_PP_  (.RESET_B(net144),
    .D(_08117_),
    .Q(_01802_),
    .CLK(clknet_leaf_50__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[67]$_DFFE_PP__145  (.L_HI(net144));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[68]$_DFFE_PP_  (.RESET_B(net145),
    .D(_08116_),
    .Q(_01803_),
    .CLK(clknet_leaf_50__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[68]$_DFFE_PP__146  (.L_HI(net145));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[69]$_DFFE_PP_  (.RESET_B(net146),
    .D(_08115_),
    .Q(_01804_),
    .CLK(clknet_leaf_51__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[69]$_DFFE_PP__147  (.L_HI(net146));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[6]$_DFFE_PP_  (.RESET_B(net147),
    .D(_08114_),
    .Q(_01805_),
    .CLK(clknet_leaf_0__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[6]$_DFFE_PP__148  (.L_HI(net147));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[70]$_DFFE_PP_  (.RESET_B(net148),
    .D(_08113_),
    .Q(_01806_),
    .CLK(clknet_leaf_51__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[70]$_DFFE_PP__149  (.L_HI(net148));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[71]$_DFFE_PP_  (.RESET_B(net149),
    .D(_08112_),
    .Q(_01807_),
    .CLK(clknet_leaf_0__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[71]$_DFFE_PP__150  (.L_HI(net149));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[72]$_DFFE_PP_  (.RESET_B(net150),
    .D(_08111_),
    .Q(_01808_),
    .CLK(clknet_leaf_51__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[72]$_DFFE_PP__151  (.L_HI(net150));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[73]$_DFFE_PP_  (.RESET_B(net151),
    .D(_08110_),
    .Q(_01809_),
    .CLK(clknet_leaf_48__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[73]$_DFFE_PP__152  (.L_HI(net151));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[74]$_DFFE_PP_  (.RESET_B(net152),
    .D(_08109_),
    .Q(_01810_),
    .CLK(clknet_leaf_50__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[74]$_DFFE_PP__153  (.L_HI(net152));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[75]$_DFFE_PP_  (.RESET_B(net153),
    .D(_08107_),
    .Q(_01811_),
    .CLK(clknet_leaf_50__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[75]$_DFFE_PP__154  (.L_HI(net153));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[76]$_DFFE_PP_  (.RESET_B(net154),
    .D(_08106_),
    .Q(_01812_),
    .CLK(clknet_leaf_50__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[76]$_DFFE_PP__155  (.L_HI(net154));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[77]$_DFFE_PP_  (.RESET_B(net155),
    .D(_08105_),
    .Q(_01813_),
    .CLK(clknet_leaf_48__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[77]$_DFFE_PP__156  (.L_HI(net155));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[78]$_DFFE_PP_  (.RESET_B(net156),
    .D(_08104_),
    .Q(_01814_),
    .CLK(clknet_leaf_49__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[78]$_DFFE_PP__157  (.L_HI(net156));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[79]$_DFFE_PP_  (.RESET_B(net157),
    .D(_08103_),
    .Q(_01815_),
    .CLK(clknet_leaf_50__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[79]$_DFFE_PP__158  (.L_HI(net157));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[7]$_DFFE_PP_  (.RESET_B(net158),
    .D(_08101_),
    .Q(_01816_),
    .CLK(clknet_leaf_0__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[7]$_DFFE_PP__159  (.L_HI(net158));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[80]$_DFFE_PP_  (.RESET_B(net159),
    .D(_08099_),
    .Q(_01817_),
    .CLK(clknet_leaf_48__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[80]$_DFFE_PP__160  (.L_HI(net159));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[81]$_DFFE_PP_  (.RESET_B(net160),
    .D(_08098_),
    .Q(_01818_),
    .CLK(clknet_leaf_48__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[81]$_DFFE_PP__161  (.L_HI(net160));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[82]$_DFFE_PP_  (.RESET_B(net161),
    .D(_08097_),
    .Q(_01819_),
    .CLK(clknet_leaf_51__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[82]$_DFFE_PP__162  (.L_HI(net161));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[83]$_DFFE_PP_  (.RESET_B(net162),
    .D(_08096_),
    .Q(_01820_),
    .CLK(clknet_leaf_50__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[83]$_DFFE_PP__163  (.L_HI(net162));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[84]$_DFFE_PP_  (.RESET_B(net163),
    .D(_08095_),
    .Q(_01821_),
    .CLK(clknet_leaf_51__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[84]$_DFFE_PP__164  (.L_HI(net163));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[85]$_DFFE_PP_  (.RESET_B(net164),
    .D(_08094_),
    .Q(_01822_),
    .CLK(clknet_leaf_51__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[85]$_DFFE_PP__165  (.L_HI(net164));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[86]$_DFFE_PP_  (.RESET_B(net165),
    .D(_08093_),
    .Q(_01823_),
    .CLK(clknet_leaf_51__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[86]$_DFFE_PP__166  (.L_HI(net165));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[87]$_DFFE_PP_  (.RESET_B(net166),
    .D(_08092_),
    .Q(_01824_),
    .CLK(clknet_leaf_0__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[87]$_DFFE_PP__167  (.L_HI(net166));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[88]$_DFFE_PP_  (.RESET_B(net167),
    .D(_08091_),
    .Q(_01825_),
    .CLK(clknet_leaf_51__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[88]$_DFFE_PP__168  (.L_HI(net167));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[89]$_DFFE_PP_  (.RESET_B(net168),
    .D(_08089_),
    .Q(_01826_),
    .CLK(clknet_leaf_48__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[89]$_DFFE_PP__169  (.L_HI(net168));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[8]$_DFFE_PP_  (.RESET_B(net169),
    .D(_08088_),
    .Q(_01827_),
    .CLK(clknet_leaf_0__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[8]$_DFFE_PP__170  (.L_HI(net169));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[90]$_DFFE_PP_  (.RESET_B(net170),
    .D(_08087_),
    .Q(_01828_),
    .CLK(clknet_leaf_51__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[90]$_DFFE_PP__171  (.L_HI(net170));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[91]$_DFFE_PP_  (.RESET_B(net171),
    .D(_08086_),
    .Q(_01829_),
    .CLK(clknet_leaf_50__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[91]$_DFFE_PP__172  (.L_HI(net171));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[92]$_DFFE_PP_  (.RESET_B(net172),
    .D(_08085_),
    .Q(_01830_),
    .CLK(clknet_leaf_49__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[92]$_DFFE_PP__173  (.L_HI(net172));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[93]$_DFFE_PP_  (.RESET_B(net173),
    .D(_08084_),
    .Q(_01831_),
    .CLK(clknet_leaf_48__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[93]$_DFFE_PP__174  (.L_HI(net173));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[94]$_DFFE_PP_  (.RESET_B(net174),
    .D(_08083_),
    .Q(_01832_),
    .CLK(clknet_leaf_49__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[94]$_DFFE_PP__175  (.L_HI(net174));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[95]$_DFFE_PP_  (.RESET_B(net175),
    .D(_08082_),
    .Q(_01833_),
    .CLK(clknet_leaf_50__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[95]$_DFFE_PP__176  (.L_HI(net175));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[9]$_DFFE_PP_  (.RESET_B(net176),
    .D(_08080_),
    .Q(_01834_),
    .CLK(clknet_leaf_48__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[9]$_DFFE_PP__177  (.L_HI(net176));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0]$_DFF_PN0_  (.RESET_B(net8239),
    .D(_08075_),
    .Q(_01835_),
    .CLK(clknet_leaf_44__06563_));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[1]$_DFF_PN0_  (.RESET_B(net8239),
    .D(_08073_),
    .Q(_01836_),
    .CLK(clknet_leaf_44__06563_));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[2]$_DFF_PN0_  (.RESET_B(net8239),
    .D(_08070_),
    .Q(_01837_),
    .CLK(clknet_leaf_44__06563_));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[0]$_DFF_PN0_  (.RESET_B(net8239),
    .D(_08060_),
    .Q(_01838_),
    .CLK(clknet_leaf_44__06563_));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[1]$_DFF_PN0_  (.RESET_B(net8240),
    .D(_08057_),
    .Q(_01839_),
    .CLK(clknet_leaf_44__06563_));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[10]$_DFFE_PP_  (.RESET_B(net177),
    .D(_08054_),
    .Q(_01840_),
    .CLK(clknet_leaf_46__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[10]$_DFFE_PP__178  (.L_HI(net177));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[11]$_DFFE_PP_  (.RESET_B(net178),
    .D(_08045_),
    .Q(_01841_),
    .CLK(clknet_leaf_37__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[11]$_DFFE_PP__179  (.L_HI(net178));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[12]$_DFFE_PP_  (.RESET_B(net179),
    .D(_08035_),
    .Q(_01842_),
    .CLK(clknet_leaf_47__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[12]$_DFFE_PP__180  (.L_HI(net179));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[13]$_DFFE_PP_  (.RESET_B(net180),
    .D(_08024_),
    .Q(_01843_),
    .CLK(clknet_leaf_47__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[13]$_DFFE_PP__181  (.L_HI(net180));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[14]$_DFFE_PP_  (.RESET_B(net181),
    .D(_08009_),
    .Q(_01844_),
    .CLK(clknet_leaf_47__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[14]$_DFFE_PP__182  (.L_HI(net181));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[15]$_DFFE_PP_  (.RESET_B(net182),
    .D(_07998_),
    .Q(_01845_),
    .CLK(clknet_leaf_47__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[15]$_DFFE_PP__183  (.L_HI(net182));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[16]$_DFFE_PP_  (.RESET_B(net183),
    .D(_07989_),
    .Q(_01846_),
    .CLK(clknet_leaf_47__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[16]$_DFFE_PP__184  (.L_HI(net183));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[17]$_DFFE_PP_  (.RESET_B(net184),
    .D(_07976_),
    .Q(_01847_),
    .CLK(clknet_leaf_47__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[17]$_DFFE_PP__185  (.L_HI(net184));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[18]$_DFFE_PP_  (.RESET_B(net185),
    .D(_07965_),
    .Q(_01848_),
    .CLK(clknet_leaf_47__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[18]$_DFFE_PP__186  (.L_HI(net185));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[19]$_DFFE_PP_  (.RESET_B(net186),
    .D(_07955_),
    .Q(_01849_),
    .CLK(clknet_leaf_47__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[19]$_DFFE_PP__187  (.L_HI(net186));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[20]$_DFFE_PP_  (.RESET_B(net187),
    .D(_07943_),
    .Q(_01850_),
    .CLK(clknet_leaf_46__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[20]$_DFFE_PP__188  (.L_HI(net187));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[21]$_DFFE_PP_  (.RESET_B(net188),
    .D(_07933_),
    .Q(_01851_),
    .CLK(clknet_leaf_46__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[21]$_DFFE_PP__189  (.L_HI(net188));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[22]$_DFFE_PP_  (.RESET_B(net189),
    .D(_07923_),
    .Q(_01852_),
    .CLK(clknet_leaf_46__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[22]$_DFFE_PP__190  (.L_HI(net189));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[23]$_DFFE_PP_  (.RESET_B(net190),
    .D(_07914_),
    .Q(_01853_),
    .CLK(clknet_leaf_46__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[23]$_DFFE_PP__191  (.L_HI(net190));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[24]$_DFFE_PP_  (.RESET_B(net191),
    .D(_07905_),
    .Q(_01854_),
    .CLK(clknet_leaf_46__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[24]$_DFFE_PP__192  (.L_HI(net191));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[25]$_DFFE_PP_  (.RESET_B(net192),
    .D(_07894_),
    .Q(_01855_),
    .CLK(clknet_leaf_46__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[25]$_DFFE_PP__193  (.L_HI(net192));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[26]$_DFFE_PP_  (.RESET_B(net193),
    .D(_07885_),
    .Q(_01856_),
    .CLK(clknet_leaf_46__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[26]$_DFFE_PP__194  (.L_HI(net193));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[27]$_DFFE_PP_  (.RESET_B(net194),
    .D(_07875_),
    .Q(_01857_),
    .CLK(clknet_leaf_37__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[27]$_DFFE_PP__195  (.L_HI(net194));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[28]$_DFFE_PP_  (.RESET_B(net195),
    .D(_07865_),
    .Q(_01858_),
    .CLK(clknet_leaf_37__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[28]$_DFFE_PP__196  (.L_HI(net195));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[29]$_DFFE_PP_  (.RESET_B(net196),
    .D(_07855_),
    .Q(_01859_),
    .CLK(clknet_leaf_37__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[29]$_DFFE_PP__197  (.L_HI(net196));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[2]$_DFFE_PP_  (.RESET_B(net197),
    .D(_07846_),
    .Q(_01860_),
    .CLK(clknet_leaf_47__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[2]$_DFFE_PP__198  (.L_HI(net197));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[30]$_DFFE_PP_  (.RESET_B(net198),
    .D(_07819_),
    .Q(_01861_),
    .CLK(clknet_leaf_37__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[30]$_DFFE_PP__199  (.L_HI(net198));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[31]$_DFFE_PP_  (.RESET_B(net199),
    .D(_07809_),
    .Q(_01862_),
    .CLK(clknet_leaf_47__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[31]$_DFFE_PP__200  (.L_HI(net199));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[3]$_DFFE_PP_  (.RESET_B(net200),
    .D(_07796_),
    .Q(_01863_),
    .CLK(clknet_leaf_45__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[3]$_DFFE_PP__201  (.L_HI(net200));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[4]$_DFFE_PP_  (.RESET_B(net201),
    .D(_07769_),
    .Q(_01864_),
    .CLK(clknet_leaf_46__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[4]$_DFFE_PP__202  (.L_HI(net201));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[5]$_DFFE_PP_  (.RESET_B(net202),
    .D(_07758_),
    .Q(_01865_),
    .CLK(clknet_leaf_46__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[5]$_DFFE_PP__203  (.L_HI(net202));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[6]$_DFFE_PP_  (.RESET_B(net203),
    .D(_07743_),
    .Q(_01866_),
    .CLK(clknet_leaf_45__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[6]$_DFFE_PP__204  (.L_HI(net203));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[7]$_DFFE_PP_  (.RESET_B(net204),
    .D(_07731_),
    .Q(_01867_),
    .CLK(clknet_leaf_47__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[7]$_DFFE_PP__205  (.L_HI(net204));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[8]$_DFFE_PP_  (.RESET_B(net205),
    .D(_07725_),
    .Q(_01868_),
    .CLK(clknet_leaf_46__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[8]$_DFFE_PP__206  (.L_HI(net205));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[9]$_DFFE_PP_  (.RESET_B(net206),
    .D(_07713_),
    .Q(_01869_),
    .CLK(clknet_leaf_46__06563_));
 sg13g2_tiehi \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[9]$_DFFE_PP__207  (.L_HI(net206));
 sg13g2_dfrbpq_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q$_DFF_PN0_  (.RESET_B(net8239),
    .D(_07670_),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .CLK(clknet_leaf_45__06563_));
 sg13g2_dfrbpq_1 \if_stage_i.illegal_c_insn_id_o$_DFFE_PP_  (.RESET_B(net207),
    .D(_07656_),
    .Q(\id_stage_i.decoder_i.illegal_c_insn_i ),
    .CLK(clknet_leaf_2__06563_));
 sg13g2_tiehi \if_stage_i.illegal_c_insn_id_o$_DFFE_PP__208  (.L_HI(net207));
 sg13g2_dfrbpq_1 \if_stage_i.instr_fetch_err_o$_DFFE_PP_  (.RESET_B(net208),
    .D(_07641_),
    .Q(\id_stage_i.controller_i.instr_fetch_err_i ),
    .CLK(clknet_leaf_41__06563_));
 sg13g2_tiehi \if_stage_i.instr_fetch_err_o$_DFFE_PP__209  (.L_HI(net208));
 sg13g2_dfrbpq_1 \if_stage_i.instr_fetch_err_plus2_o$_SDFFCE_PN0P_  (.RESET_B(net209),
    .D(_07631_),
    .Q(\id_stage_i.controller_i.instr_fetch_err_plus2_i ),
    .CLK(clknet_leaf_44__06563_));
 sg13g2_tiehi \if_stage_i.instr_fetch_err_plus2_o$_SDFFCE_PN0P__210  (.L_HI(net209));
 sg13g2_dfrbpq_1 \if_stage_i.instr_is_compressed_id_o$_DFFE_PP_  (.RESET_B(net210),
    .D(_07626_),
    .Q(\id_stage_i.controller_i.instr_is_compressed_i ),
    .CLK(clknet_leaf_43__06563_));
 sg13g2_tiehi \if_stage_i.instr_is_compressed_id_o$_DFFE_PP__211  (.L_HI(net210));
 sg13g2_dfrbpq_1 \if_stage_i.instr_rdata_c_id_o[0]$_DFFE_PP_  (.RESET_B(net211),
    .D(_07625_),
    .Q(_01870_),
    .CLK(clknet_leaf_44__06563_));
 sg13g2_tiehi \if_stage_i.instr_rdata_c_id_o[0]$_DFFE_PP__212  (.L_HI(net211));
 sg13g2_dfrbpq_1 \if_stage_i.instr_rdata_c_id_o[10]$_DFFE_PP_  (.RESET_B(net212),
    .D(_07624_),
    .Q(_01871_),
    .CLK(clknet_leaf_44__06563_));
 sg13g2_tiehi \if_stage_i.instr_rdata_c_id_o[10]$_DFFE_PP__213  (.L_HI(net212));
 sg13g2_dfrbpq_1 \if_stage_i.instr_rdata_c_id_o[11]$_DFFE_PP_  (.RESET_B(net213),
    .D(_07623_),
    .Q(_01872_),
    .CLK(clknet_leaf_43__06563_));
 sg13g2_tiehi \if_stage_i.instr_rdata_c_id_o[11]$_DFFE_PP__214  (.L_HI(net213));
 sg13g2_dfrbpq_1 \if_stage_i.instr_rdata_c_id_o[12]$_DFFE_PP_  (.RESET_B(net214),
    .D(_07621_),
    .Q(_01873_),
    .CLK(clknet_leaf_43__06563_));
 sg13g2_tiehi \if_stage_i.instr_rdata_c_id_o[12]$_DFFE_PP__215  (.L_HI(net214));
 sg13g2_dfrbpq_1 \if_stage_i.instr_rdata_c_id_o[13]$_DFFE_PP_  (.RESET_B(net215),
    .D(_07620_),
    .Q(_01874_),
    .CLK(clknet_leaf_43__06563_));
 sg13g2_tiehi \if_stage_i.instr_rdata_c_id_o[13]$_DFFE_PP__216  (.L_HI(net215));
 sg13g2_dfrbpq_1 \if_stage_i.instr_rdata_c_id_o[14]$_DFFE_PP_  (.RESET_B(net216),
    .D(_07618_),
    .Q(_01875_),
    .CLK(clknet_leaf_44__06563_));
 sg13g2_tiehi \if_stage_i.instr_rdata_c_id_o[14]$_DFFE_PP__217  (.L_HI(net216));
 sg13g2_dfrbpq_1 \if_stage_i.instr_rdata_c_id_o[15]$_DFFE_PP_  (.RESET_B(net217),
    .D(_07617_),
    .Q(_01876_),
    .CLK(clknet_leaf_44__06563_));
 sg13g2_tiehi \if_stage_i.instr_rdata_c_id_o[15]$_DFFE_PP__218  (.L_HI(net217));
 sg13g2_dfrbpq_1 \if_stage_i.instr_rdata_c_id_o[1]$_DFFE_PP_  (.RESET_B(net218),
    .D(_07615_),
    .Q(_01877_),
    .CLK(clknet_leaf_42__06563_));
 sg13g2_tiehi \if_stage_i.instr_rdata_c_id_o[1]$_DFFE_PP__219  (.L_HI(net218));
 sg13g2_dfrbpq_1 \if_stage_i.instr_rdata_c_id_o[2]$_DFFE_PP_  (.RESET_B(net219),
    .D(_07613_),
    .Q(_01878_),
    .CLK(clknet_leaf_43__06563_));
 sg13g2_tiehi \if_stage_i.instr_rdata_c_id_o[2]$_DFFE_PP__220  (.L_HI(net219));
 sg13g2_dfrbpq_1 \if_stage_i.instr_rdata_c_id_o[3]$_DFFE_PP_  (.RESET_B(net220),
    .D(_07612_),
    .Q(_01879_),
    .CLK(clknet_leaf_43__06563_));
 sg13g2_tiehi \if_stage_i.instr_rdata_c_id_o[3]$_DFFE_PP__221  (.L_HI(net220));
 sg13g2_dfrbpq_1 \if_stage_i.instr_rdata_c_id_o[4]$_DFFE_PP_  (.RESET_B(net221),
    .D(_07611_),
    .Q(_01880_),
    .CLK(clknet_leaf_43__06563_));
 sg13g2_tiehi \if_stage_i.instr_rdata_c_id_o[4]$_DFFE_PP__222  (.L_HI(net221));
 sg13g2_dfrbpq_1 \if_stage_i.instr_rdata_c_id_o[5]$_DFFE_PP_  (.RESET_B(net222),
    .D(_07610_),
    .Q(_01881_),
    .CLK(clknet_leaf_43__06563_));
 sg13g2_tiehi \if_stage_i.instr_rdata_c_id_o[5]$_DFFE_PP__223  (.L_HI(net222));
 sg13g2_dfrbpq_1 \if_stage_i.instr_rdata_c_id_o[6]$_DFFE_PP_  (.RESET_B(net223),
    .D(_07609_),
    .Q(_01882_),
    .CLK(clknet_leaf_43__06563_));
 sg13g2_tiehi \if_stage_i.instr_rdata_c_id_o[6]$_DFFE_PP__224  (.L_HI(net223));
 sg13g2_dfrbpq_1 \if_stage_i.instr_rdata_c_id_o[7]$_DFFE_PP_  (.RESET_B(net224),
    .D(_07607_),
    .Q(_01883_),
    .CLK(clknet_leaf_43__06563_));
 sg13g2_tiehi \if_stage_i.instr_rdata_c_id_o[7]$_DFFE_PP__225  (.L_HI(net224));
 sg13g2_dfrbpq_1 \if_stage_i.instr_rdata_c_id_o[8]$_DFFE_PP_  (.RESET_B(net225),
    .D(_07606_),
    .Q(_01884_),
    .CLK(clknet_leaf_43__06563_));
 sg13g2_tiehi \if_stage_i.instr_rdata_c_id_o[8]$_DFFE_PP__226  (.L_HI(net225));
 sg13g2_dfrbpq_1 \if_stage_i.instr_rdata_c_id_o[9]$_DFFE_PP_  (.RESET_B(net226),
    .D(_07604_),
    .Q(_01885_),
    .CLK(clknet_leaf_43__06563_));
 sg13g2_tiehi \if_stage_i.instr_rdata_c_id_o[9]$_DFFE_PP__227  (.L_HI(net226));
 sg13g2_dfrbpq_1 \if_stage_i.instr_rdata_id_o[0]$_DFFE_PP_  (.RESET_B(net227),
    .D(_07603_),
    .Q(_01886_),
    .CLK(clknet_leaf_43__06563_));
 sg13g2_tiehi \if_stage_i.instr_rdata_id_o[0]$_DFFE_PP__228  (.L_HI(net227));
 sg13g2_dfrbpq_1 \if_stage_i.instr_rdata_id_o[10]$_DFFE_PP_  (.RESET_B(net228),
    .D(_07600_),
    .Q(_01887_),
    .CLK(clknet_leaf_43__06563_));
 sg13g2_tiehi \if_stage_i.instr_rdata_id_o[10]$_DFFE_PP__229  (.L_HI(net228));
 sg13g2_dfrbpq_1 \if_stage_i.instr_rdata_id_o[11]$_DFFE_PP_  (.RESET_B(net229),
    .D(_07588_),
    .Q(_01888_),
    .CLK(clknet_leaf_1__06563_));
 sg13g2_tiehi \if_stage_i.instr_rdata_id_o[11]$_DFFE_PP__230  (.L_HI(net229));
 sg13g2_dfrbpq_1 \if_stage_i.instr_rdata_id_o[12]$_DFFE_PP_  (.RESET_B(net230),
    .D(_07580_),
    .Q(_01889_),
    .CLK(clknet_leaf_43__06563_));
 sg13g2_tiehi \if_stage_i.instr_rdata_id_o[12]$_DFFE_PP__231  (.L_HI(net230));
 sg13g2_dfrbpq_1 \if_stage_i.instr_rdata_id_o[13]$_DFFE_PP_  (.RESET_B(net231),
    .D(_07565_),
    .Q(_01890_),
    .CLK(clknet_leaf_2__06563_));
 sg13g2_tiehi \if_stage_i.instr_rdata_id_o[13]$_DFFE_PP__232  (.L_HI(net231));
 sg13g2_dfrbpq_1 \if_stage_i.instr_rdata_id_o[14]$_DFFE_PP_  (.RESET_B(net232),
    .D(_07554_),
    .Q(_01891_),
    .CLK(clknet_leaf_42__06563_));
 sg13g2_tiehi \if_stage_i.instr_rdata_id_o[14]$_DFFE_PP__233  (.L_HI(net232));
 sg13g2_dfrbpq_1 \if_stage_i.instr_rdata_id_o[15]$_DFFE_PP_  (.RESET_B(net233),
    .D(_07547_),
    .Q(_01892_),
    .CLK(clknet_leaf_1__06563_));
 sg13g2_tiehi \if_stage_i.instr_rdata_id_o[15]$_DFFE_PP__234  (.L_HI(net233));
 sg13g2_dfrbpq_1 \if_stage_i.instr_rdata_id_o[16]$_DFFE_PP_  (.RESET_B(net234),
    .D(_07534_),
    .Q(_01893_),
    .CLK(clknet_leaf_1__06563_));
 sg13g2_tiehi \if_stage_i.instr_rdata_id_o[16]$_DFFE_PP__235  (.L_HI(net234));
 sg13g2_dfrbpq_1 \if_stage_i.instr_rdata_id_o[17]$_DFFE_PP_  (.RESET_B(net235),
    .D(_07511_),
    .Q(_01894_),
    .CLK(clknet_leaf_1__06563_));
 sg13g2_tiehi \if_stage_i.instr_rdata_id_o[17]$_DFFE_PP__236  (.L_HI(net235));
 sg13g2_dfrbpq_1 \if_stage_i.instr_rdata_id_o[18]$_DFFE_PP_  (.RESET_B(net236),
    .D(_07496_),
    .Q(_01895_),
    .CLK(clknet_leaf_1__06563_));
 sg13g2_tiehi \if_stage_i.instr_rdata_id_o[18]$_DFFE_PP__237  (.L_HI(net236));
 sg13g2_dfrbpq_1 \if_stage_i.instr_rdata_id_o[19]$_DFFE_PP_  (.RESET_B(net237),
    .D(_07474_),
    .Q(_01896_),
    .CLK(clknet_leaf_43__06563_));
 sg13g2_tiehi \if_stage_i.instr_rdata_id_o[19]$_DFFE_PP__238  (.L_HI(net237));
 sg13g2_dfrbpq_1 \if_stage_i.instr_rdata_id_o[1]$_DFFE_PP_  (.RESET_B(net238),
    .D(_07461_),
    .Q(_01897_),
    .CLK(clknet_leaf_43__06563_));
 sg13g2_tiehi \if_stage_i.instr_rdata_id_o[1]$_DFFE_PP__239  (.L_HI(net238));
 sg13g2_dfrbpq_1 \if_stage_i.instr_rdata_id_o[20]$_DFFE_PP_  (.RESET_B(net239),
    .D(_07459_),
    .Q(_01898_),
    .CLK(clknet_leaf_2__06563_));
 sg13g2_tiehi \if_stage_i.instr_rdata_id_o[20]$_DFFE_PP__240  (.L_HI(net239));
 sg13g2_dfrbpq_1 \if_stage_i.instr_rdata_id_o[21]$_DFFE_PP_  (.RESET_B(net240),
    .D(_07437_),
    .Q(_01899_),
    .CLK(clknet_leaf_1__06563_));
 sg13g2_tiehi \if_stage_i.instr_rdata_id_o[21]$_DFFE_PP__241  (.L_HI(net240));
 sg13g2_dfrbpq_1 \if_stage_i.instr_rdata_id_o[22]$_DFFE_PP_  (.RESET_B(net241),
    .D(_07421_),
    .Q(_01900_),
    .CLK(clknet_leaf_1__06563_));
 sg13g2_tiehi \if_stage_i.instr_rdata_id_o[22]$_DFFE_PP__242  (.L_HI(net241));
 sg13g2_dfrbpq_1 \if_stage_i.instr_rdata_id_o[23]$_DFFE_PP_  (.RESET_B(net242),
    .D(_07401_),
    .Q(_01901_),
    .CLK(clknet_leaf_1__06563_));
 sg13g2_tiehi \if_stage_i.instr_rdata_id_o[23]$_DFFE_PP__243  (.L_HI(net242));
 sg13g2_dfrbpq_1 \if_stage_i.instr_rdata_id_o[24]$_DFFE_PP_  (.RESET_B(net243),
    .D(_07383_),
    .Q(_01902_),
    .CLK(clknet_leaf_1__06563_));
 sg13g2_tiehi \if_stage_i.instr_rdata_id_o[24]$_DFFE_PP__244  (.L_HI(net243));
 sg13g2_dfrbpq_1 \if_stage_i.instr_rdata_id_o[25]$_DFFE_PP_  (.RESET_B(net244),
    .D(_07369_),
    .Q(_01903_),
    .CLK(clknet_leaf_2__06563_));
 sg13g2_tiehi \if_stage_i.instr_rdata_id_o[25]$_DFFE_PP__245  (.L_HI(net244));
 sg13g2_dfrbpq_1 \if_stage_i.instr_rdata_id_o[26]$_DFFE_PP_  (.RESET_B(net245),
    .D(_07356_),
    .Q(_01904_),
    .CLK(clknet_leaf_42__06563_));
 sg13g2_tiehi \if_stage_i.instr_rdata_id_o[26]$_DFFE_PP__246  (.L_HI(net245));
 sg13g2_dfrbpq_1 \if_stage_i.instr_rdata_id_o[27]$_DFFE_PP_  (.RESET_B(net246),
    .D(_07334_),
    .Q(_01905_),
    .CLK(clknet_leaf_43__06563_));
 sg13g2_tiehi \if_stage_i.instr_rdata_id_o[27]$_DFFE_PP__247  (.L_HI(net246));
 sg13g2_dfrbpq_1 \if_stage_i.instr_rdata_id_o[28]$_DFFE_PP_  (.RESET_B(net247),
    .D(_07314_),
    .Q(_01906_),
    .CLK(clknet_leaf_43__06563_));
 sg13g2_tiehi \if_stage_i.instr_rdata_id_o[28]$_DFFE_PP__248  (.L_HI(net247));
 sg13g2_dfrbpq_1 \if_stage_i.instr_rdata_id_o[29]$_DFFE_PP_  (.RESET_B(net248),
    .D(_07298_),
    .Q(_01907_),
    .CLK(clknet_leaf_43__06563_));
 sg13g2_tiehi \if_stage_i.instr_rdata_id_o[29]$_DFFE_PP__249  (.L_HI(net248));
 sg13g2_dfrbpq_1 \if_stage_i.instr_rdata_id_o[2]$_DFFE_PP_  (.RESET_B(net249),
    .D(_07283_),
    .Q(_01908_),
    .CLK(clknet_leaf_42__06563_));
 sg13g2_tiehi \if_stage_i.instr_rdata_id_o[2]$_DFFE_PP__250  (.L_HI(net249));
 sg13g2_dfrbpq_1 \if_stage_i.instr_rdata_id_o[30]$_DFFE_PP_  (.RESET_B(net250),
    .D(_07277_),
    .Q(_01909_),
    .CLK(clknet_leaf_42__06563_));
 sg13g2_tiehi \if_stage_i.instr_rdata_id_o[30]$_DFFE_PP__251  (.L_HI(net250));
 sg13g2_dfrbpq_1 \if_stage_i.instr_rdata_id_o[31]$_DFFE_PP_  (.RESET_B(net251),
    .D(_07262_),
    .Q(_01910_),
    .CLK(clknet_leaf_42__06563_));
 sg13g2_tiehi \if_stage_i.instr_rdata_id_o[31]$_DFFE_PP__252  (.L_HI(net251));
 sg13g2_dfrbpq_1 \if_stage_i.instr_rdata_id_o[3]$_DFFE_PP_  (.RESET_B(net252),
    .D(_07251_),
    .Q(_01911_),
    .CLK(clknet_leaf_42__06563_));
 sg13g2_tiehi \if_stage_i.instr_rdata_id_o[3]$_DFFE_PP__253  (.L_HI(net252));
 sg13g2_dfrbpq_1 \if_stage_i.instr_rdata_id_o[4]$_DFFE_PP_  (.RESET_B(net253),
    .D(_07248_),
    .Q(_01912_),
    .CLK(clknet_leaf_44__06563_));
 sg13g2_tiehi \if_stage_i.instr_rdata_id_o[4]$_DFFE_PP__254  (.L_HI(net253));
 sg13g2_dfrbpq_1 \if_stage_i.instr_rdata_id_o[5]$_DFFE_PP_  (.RESET_B(net254),
    .D(_07236_),
    .Q(_01913_),
    .CLK(clknet_leaf_44__06563_));
 sg13g2_tiehi \if_stage_i.instr_rdata_id_o[5]$_DFFE_PP__255  (.L_HI(net254));
 sg13g2_dfrbpq_1 \if_stage_i.instr_rdata_id_o[6]$_DFFE_PP_  (.RESET_B(net255),
    .D(_07222_),
    .Q(_01914_),
    .CLK(clknet_leaf_42__06563_));
 sg13g2_tiehi \if_stage_i.instr_rdata_id_o[6]$_DFFE_PP__256  (.L_HI(net255));
 sg13g2_dfrbpq_1 \if_stage_i.instr_rdata_id_o[7]$_DFFE_PP_  (.RESET_B(net256),
    .D(_07212_),
    .Q(_01915_),
    .CLK(clknet_leaf_1__06563_));
 sg13g2_tiehi \if_stage_i.instr_rdata_id_o[7]$_DFFE_PP__257  (.L_HI(net256));
 sg13g2_dfrbpq_1 \if_stage_i.instr_rdata_id_o[8]$_DFFE_PP_  (.RESET_B(net257),
    .D(_07187_),
    .Q(_01916_),
    .CLK(clknet_leaf_43__06563_));
 sg13g2_tiehi \if_stage_i.instr_rdata_id_o[8]$_DFFE_PP__258  (.L_HI(net257));
 sg13g2_dfrbpq_1 \if_stage_i.instr_rdata_id_o[9]$_DFFE_PP_  (.RESET_B(net258),
    .D(_07166_),
    .Q(_01917_),
    .CLK(clknet_leaf_1__06563_));
 sg13g2_tiehi \if_stage_i.instr_rdata_id_o[9]$_DFFE_PP__259  (.L_HI(net258));
 sg13g2_dfrbpq_1 \if_stage_i.instr_valid_id_o$_DFF_PN0_  (.RESET_B(net8241),
    .D(_07096_),
    .Q(\id_stage_i.controller_i.instr_valid_i ),
    .CLK(clknet_leaf_40__06563_));
 sg13g2_dfrbpq_1 \if_stage_i.pc_id_o[10]$_DFFE_PP_  (.RESET_B(net259),
    .D(_07080_),
    .Q(_01918_),
    .CLK(clknet_leaf_38__06563_));
 sg13g2_tiehi \if_stage_i.pc_id_o[10]$_DFFE_PP__260  (.L_HI(net259));
 sg13g2_dfrbpq_1 \if_stage_i.pc_id_o[11]$_DFFE_PP_  (.RESET_B(net260),
    .D(_07078_),
    .Q(_01919_),
    .CLK(clknet_leaf_38__06563_));
 sg13g2_tiehi \if_stage_i.pc_id_o[11]$_DFFE_PP__261  (.L_HI(net260));
 sg13g2_dfrbpq_1 \if_stage_i.pc_id_o[12]$_DFFE_PP_  (.RESET_B(net261),
    .D(_07077_),
    .Q(_01920_),
    .CLK(clknet_leaf_38__06563_));
 sg13g2_tiehi \if_stage_i.pc_id_o[12]$_DFFE_PP__262  (.L_HI(net261));
 sg13g2_dfrbpq_1 \if_stage_i.pc_id_o[13]$_DFFE_PP_  (.RESET_B(net262),
    .D(_07076_),
    .Q(_01921_),
    .CLK(clknet_leaf_38__06563_));
 sg13g2_tiehi \if_stage_i.pc_id_o[13]$_DFFE_PP__263  (.L_HI(net262));
 sg13g2_dfrbpq_1 \if_stage_i.pc_id_o[14]$_DFFE_PP_  (.RESET_B(net263),
    .D(_07075_),
    .Q(_01922_),
    .CLK(clknet_leaf_39__06563_));
 sg13g2_tiehi \if_stage_i.pc_id_o[14]$_DFFE_PP__264  (.L_HI(net263));
 sg13g2_dfrbpq_1 \if_stage_i.pc_id_o[15]$_DFFE_PP_  (.RESET_B(net264),
    .D(_07074_),
    .Q(_01923_),
    .CLK(clknet_leaf_38__06563_));
 sg13g2_tiehi \if_stage_i.pc_id_o[15]$_DFFE_PP__265  (.L_HI(net264));
 sg13g2_dfrbpq_1 \if_stage_i.pc_id_o[16]$_DFFE_PP_  (.RESET_B(net265),
    .D(_07073_),
    .Q(_01924_),
    .CLK(clknet_leaf_39__06563_));
 sg13g2_tiehi \if_stage_i.pc_id_o[16]$_DFFE_PP__266  (.L_HI(net265));
 sg13g2_dfrbpq_1 \if_stage_i.pc_id_o[17]$_DFFE_PP_  (.RESET_B(net266),
    .D(_07072_),
    .Q(_01925_),
    .CLK(clknet_leaf_38__06563_));
 sg13g2_tiehi \if_stage_i.pc_id_o[17]$_DFFE_PP__267  (.L_HI(net266));
 sg13g2_dfrbpq_1 \if_stage_i.pc_id_o[18]$_DFFE_PP_  (.RESET_B(net267),
    .D(_07071_),
    .Q(_01926_),
    .CLK(clknet_leaf_39__06563_));
 sg13g2_tiehi \if_stage_i.pc_id_o[18]$_DFFE_PP__268  (.L_HI(net267));
 sg13g2_dfrbpq_1 \if_stage_i.pc_id_o[19]$_DFFE_PP_  (.RESET_B(net268),
    .D(_07069_),
    .Q(_01927_),
    .CLK(clknet_leaf_36__06563_));
 sg13g2_tiehi \if_stage_i.pc_id_o[19]$_DFFE_PP__269  (.L_HI(net268));
 sg13g2_dfrbpq_1 \if_stage_i.pc_id_o[1]$_DFFE_PP_  (.RESET_B(net269),
    .D(_07068_),
    .Q(_01928_),
    .CLK(clknet_leaf_42__06563_));
 sg13g2_tiehi \if_stage_i.pc_id_o[1]$_DFFE_PP__270  (.L_HI(net269));
 sg13g2_dfrbpq_1 \if_stage_i.pc_id_o[20]$_DFFE_PP_  (.RESET_B(net270),
    .D(_07067_),
    .Q(_01929_),
    .CLK(clknet_leaf_39__06563_));
 sg13g2_tiehi \if_stage_i.pc_id_o[20]$_DFFE_PP__271  (.L_HI(net270));
 sg13g2_dfrbpq_1 \if_stage_i.pc_id_o[21]$_DFFE_PP_  (.RESET_B(net271),
    .D(_07066_),
    .Q(_01930_),
    .CLK(clknet_leaf_39__06563_));
 sg13g2_tiehi \if_stage_i.pc_id_o[21]$_DFFE_PP__272  (.L_HI(net271));
 sg13g2_dfrbpq_1 \if_stage_i.pc_id_o[22]$_DFFE_PP_  (.RESET_B(net272),
    .D(_07065_),
    .Q(_01931_),
    .CLK(clknet_leaf_39__06563_));
 sg13g2_tiehi \if_stage_i.pc_id_o[22]$_DFFE_PP__273  (.L_HI(net272));
 sg13g2_dfrbpq_1 \if_stage_i.pc_id_o[23]$_DFFE_PP_  (.RESET_B(net273),
    .D(_07064_),
    .Q(_01932_),
    .CLK(clknet_leaf_39__06563_));
 sg13g2_tiehi \if_stage_i.pc_id_o[23]$_DFFE_PP__274  (.L_HI(net273));
 sg13g2_dfrbpq_1 \if_stage_i.pc_id_o[24]$_DFFE_PP_  (.RESET_B(net274),
    .D(_07063_),
    .Q(_01933_),
    .CLK(clknet_leaf_39__06563_));
 sg13g2_tiehi \if_stage_i.pc_id_o[24]$_DFFE_PP__275  (.L_HI(net274));
 sg13g2_dfrbpq_1 \if_stage_i.pc_id_o[25]$_DFFE_PP_  (.RESET_B(net275),
    .D(_07062_),
    .Q(_01934_),
    .CLK(clknet_leaf_36__06563_));
 sg13g2_tiehi \if_stage_i.pc_id_o[25]$_DFFE_PP__276  (.L_HI(net275));
 sg13g2_dfrbpq_1 \if_stage_i.pc_id_o[26]$_DFFE_PP_  (.RESET_B(net276),
    .D(_07061_),
    .Q(_01935_),
    .CLK(clknet_leaf_36__06563_));
 sg13g2_tiehi \if_stage_i.pc_id_o[26]$_DFFE_PP__277  (.L_HI(net276));
 sg13g2_dfrbpq_1 \if_stage_i.pc_id_o[27]$_DFFE_PP_  (.RESET_B(net277),
    .D(_07060_),
    .Q(_01936_),
    .CLK(clknet_leaf_39__06563_));
 sg13g2_tiehi \if_stage_i.pc_id_o[27]$_DFFE_PP__278  (.L_HI(net277));
 sg13g2_dfrbpq_1 \if_stage_i.pc_id_o[28]$_DFFE_PP_  (.RESET_B(net278),
    .D(_07059_),
    .Q(_01937_),
    .CLK(clknet_leaf_36__06563_));
 sg13g2_tiehi \if_stage_i.pc_id_o[28]$_DFFE_PP__279  (.L_HI(net278));
 sg13g2_dfrbpq_1 \if_stage_i.pc_id_o[29]$_DFFE_PP_  (.RESET_B(net279),
    .D(_07058_),
    .Q(_01938_),
    .CLK(clknet_leaf_36__06563_));
 sg13g2_tiehi \if_stage_i.pc_id_o[29]$_DFFE_PP__280  (.L_HI(net279));
 sg13g2_dfrbpq_1 \if_stage_i.pc_id_o[2]$_DFFE_PP_  (.RESET_B(net280),
    .D(_07057_),
    .Q(_01939_),
    .CLK(clknet_leaf_42__06563_));
 sg13g2_tiehi \if_stage_i.pc_id_o[2]$_DFFE_PP__281  (.L_HI(net280));
 sg13g2_dfrbpq_1 \if_stage_i.pc_id_o[30]$_DFFE_PP_  (.RESET_B(net281),
    .D(_07056_),
    .Q(_01940_),
    .CLK(clknet_leaf_36__06563_));
 sg13g2_tiehi \if_stage_i.pc_id_o[30]$_DFFE_PP__282  (.L_HI(net281));
 sg13g2_dfrbpq_1 \if_stage_i.pc_id_o[31]$_DFFE_PP_  (.RESET_B(net282),
    .D(_07055_),
    .Q(_01941_),
    .CLK(clknet_leaf_36__06563_));
 sg13g2_tiehi \if_stage_i.pc_id_o[31]$_DFFE_PP__283  (.L_HI(net282));
 sg13g2_dfrbpq_1 \if_stage_i.pc_id_o[3]$_DFFE_PP_  (.RESET_B(net283),
    .D(_07054_),
    .Q(_01942_),
    .CLK(clknet_leaf_42__06563_));
 sg13g2_tiehi \if_stage_i.pc_id_o[3]$_DFFE_PP__284  (.L_HI(net283));
 sg13g2_dfrbpq_1 \if_stage_i.pc_id_o[4]$_DFFE_PP_  (.RESET_B(net284),
    .D(_07052_),
    .Q(_01943_),
    .CLK(clknet_leaf_41__06563_));
 sg13g2_tiehi \if_stage_i.pc_id_o[4]$_DFFE_PP__285  (.L_HI(net284));
 sg13g2_dfrbpq_1 \if_stage_i.pc_id_o[5]$_DFFE_PP_  (.RESET_B(net285),
    .D(_07051_),
    .Q(_01944_),
    .CLK(clknet_leaf_38__06563_));
 sg13g2_tiehi \if_stage_i.pc_id_o[5]$_DFFE_PP__286  (.L_HI(net285));
 sg13g2_dfrbpq_1 \if_stage_i.pc_id_o[6]$_DFFE_PP_  (.RESET_B(net286),
    .D(_07050_),
    .Q(_01945_),
    .CLK(clknet_leaf_38__06563_));
 sg13g2_tiehi \if_stage_i.pc_id_o[6]$_DFFE_PP__287  (.L_HI(net286));
 sg13g2_dfrbpq_1 \if_stage_i.pc_id_o[7]$_DFFE_PP_  (.RESET_B(net287),
    .D(_07049_),
    .Q(_01946_),
    .CLK(clknet_leaf_41__06563_));
 sg13g2_tiehi \if_stage_i.pc_id_o[7]$_DFFE_PP__288  (.L_HI(net287));
 sg13g2_dfrbpq_1 \if_stage_i.pc_id_o[8]$_DFFE_PP_  (.RESET_B(net288),
    .D(_07047_),
    .Q(_01947_),
    .CLK(clknet_leaf_38__06563_));
 sg13g2_tiehi \if_stage_i.pc_id_o[8]$_DFFE_PP__289  (.L_HI(net288));
 sg13g2_dfrbpq_1 \if_stage_i.pc_id_o[9]$_DFFE_PP_  (.RESET_B(net289),
    .D(_07046_),
    .Q(_01948_),
    .CLK(clknet_leaf_38__06563_));
 sg13g2_tiehi \if_stage_i.pc_id_o[9]$_DFFE_PP__290  (.L_HI(net289));
 sg13g2_buf_1 input291 (.A(boot_addr_i[10]),
    .X(net290));
 sg13g2_buf_1 input292 (.A(boot_addr_i[11]),
    .X(net291));
 sg13g2_buf_1 input293 (.A(boot_addr_i[12]),
    .X(net292));
 sg13g2_buf_1 input294 (.A(boot_addr_i[13]),
    .X(net293));
 sg13g2_buf_1 input295 (.A(boot_addr_i[14]),
    .X(net294));
 sg13g2_buf_1 input296 (.A(boot_addr_i[15]),
    .X(net295));
 sg13g2_buf_1 input297 (.A(boot_addr_i[16]),
    .X(net296));
 sg13g2_buf_1 input298 (.A(boot_addr_i[17]),
    .X(net297));
 sg13g2_buf_1 input299 (.A(boot_addr_i[18]),
    .X(net298));
 sg13g2_buf_1 input300 (.A(boot_addr_i[19]),
    .X(net299));
 sg13g2_buf_1 input301 (.A(boot_addr_i[20]),
    .X(net300));
 sg13g2_buf_1 input302 (.A(boot_addr_i[21]),
    .X(net301));
 sg13g2_buf_1 input303 (.A(boot_addr_i[22]),
    .X(net302));
 sg13g2_buf_1 input304 (.A(boot_addr_i[23]),
    .X(net303));
 sg13g2_buf_1 input305 (.A(boot_addr_i[24]),
    .X(net304));
 sg13g2_buf_1 input306 (.A(boot_addr_i[25]),
    .X(net305));
 sg13g2_buf_1 input307 (.A(boot_addr_i[26]),
    .X(net306));
 sg13g2_buf_1 input308 (.A(boot_addr_i[27]),
    .X(net307));
 sg13g2_buf_1 input309 (.A(boot_addr_i[28]),
    .X(net308));
 sg13g2_buf_1 input310 (.A(boot_addr_i[29]),
    .X(net309));
 sg13g2_buf_1 input311 (.A(boot_addr_i[30]),
    .X(net310));
 sg13g2_buf_1 input312 (.A(boot_addr_i[31]),
    .X(net311));
 sg13g2_buf_1 input313 (.A(boot_addr_i[8]),
    .X(net312));
 sg13g2_buf_1 input314 (.A(boot_addr_i[9]),
    .X(net313));
 sg13g2_buf_1 input315 (.A(data_err_i),
    .X(net314));
 sg13g2_buf_1 input316 (.A(data_gnt_i),
    .X(net315));
 sg13g2_buf_1 input317 (.A(data_rdata_i[0]),
    .X(net316));
 sg13g2_buf_1 input318 (.A(data_rdata_i[10]),
    .X(net317));
 sg13g2_buf_1 input319 (.A(data_rdata_i[11]),
    .X(net318));
 sg13g2_buf_1 input320 (.A(data_rdata_i[12]),
    .X(net319));
 sg13g2_buf_1 input321 (.A(data_rdata_i[13]),
    .X(net320));
 sg13g2_buf_1 input322 (.A(data_rdata_i[14]),
    .X(net321));
 sg13g2_buf_1 input323 (.A(data_rdata_i[15]),
    .X(net322));
 sg13g2_buf_1 input324 (.A(data_rdata_i[16]),
    .X(net323));
 sg13g2_buf_1 input325 (.A(data_rdata_i[17]),
    .X(net324));
 sg13g2_buf_1 input326 (.A(data_rdata_i[18]),
    .X(net325));
 sg13g2_buf_1 input327 (.A(data_rdata_i[19]),
    .X(net326));
 sg13g2_buf_1 input328 (.A(data_rdata_i[1]),
    .X(net327));
 sg13g2_buf_1 input329 (.A(data_rdata_i[20]),
    .X(net328));
 sg13g2_buf_1 input330 (.A(data_rdata_i[21]),
    .X(net329));
 sg13g2_buf_1 input331 (.A(data_rdata_i[22]),
    .X(net330));
 sg13g2_buf_1 input332 (.A(data_rdata_i[23]),
    .X(net331));
 sg13g2_buf_1 input333 (.A(data_rdata_i[24]),
    .X(net332));
 sg13g2_buf_1 input334 (.A(data_rdata_i[25]),
    .X(net333));
 sg13g2_buf_1 input335 (.A(data_rdata_i[26]),
    .X(net334));
 sg13g2_buf_1 input336 (.A(data_rdata_i[27]),
    .X(net335));
 sg13g2_buf_1 input337 (.A(data_rdata_i[28]),
    .X(net336));
 sg13g2_buf_1 input338 (.A(data_rdata_i[29]),
    .X(net337));
 sg13g2_buf_1 input339 (.A(data_rdata_i[2]),
    .X(net338));
 sg13g2_buf_1 input340 (.A(data_rdata_i[30]),
    .X(net339));
 sg13g2_buf_1 input341 (.A(data_rdata_i[31]),
    .X(net340));
 sg13g2_buf_1 input342 (.A(data_rdata_i[3]),
    .X(net341));
 sg13g2_buf_1 input343 (.A(data_rdata_i[4]),
    .X(net342));
 sg13g2_buf_1 input344 (.A(data_rdata_i[5]),
    .X(net343));
 sg13g2_buf_1 input345 (.A(data_rdata_i[6]),
    .X(net344));
 sg13g2_buf_1 input346 (.A(data_rdata_i[7]),
    .X(net345));
 sg13g2_buf_1 input347 (.A(data_rdata_i[8]),
    .X(net346));
 sg13g2_buf_1 input348 (.A(data_rdata_i[9]),
    .X(net347));
 sg13g2_buf_1 input349 (.A(data_rvalid_i),
    .X(net348));
 sg13g2_buf_1 input350 (.A(debug_req_i),
    .X(net349));
 sg13g2_buf_1 input351 (.A(fetch_enable_i),
    .X(net350));
 sg13g2_buf_1 input352 (.A(hart_id_i[0]),
    .X(net351));
 sg13g2_buf_1 input353 (.A(hart_id_i[10]),
    .X(net352));
 sg13g2_buf_1 input354 (.A(hart_id_i[11]),
    .X(net353));
 sg13g2_buf_1 input355 (.A(hart_id_i[12]),
    .X(net354));
 sg13g2_buf_1 input356 (.A(hart_id_i[13]),
    .X(net355));
 sg13g2_buf_1 input357 (.A(hart_id_i[14]),
    .X(net356));
 sg13g2_buf_1 input358 (.A(hart_id_i[15]),
    .X(net357));
 sg13g2_buf_1 input359 (.A(hart_id_i[16]),
    .X(net358));
 sg13g2_buf_1 input360 (.A(hart_id_i[17]),
    .X(net359));
 sg13g2_buf_1 input361 (.A(hart_id_i[18]),
    .X(net360));
 sg13g2_buf_1 input362 (.A(hart_id_i[19]),
    .X(net361));
 sg13g2_buf_1 input363 (.A(hart_id_i[1]),
    .X(net362));
 sg13g2_buf_1 input364 (.A(hart_id_i[20]),
    .X(net363));
 sg13g2_buf_1 input365 (.A(hart_id_i[21]),
    .X(net364));
 sg13g2_buf_1 input366 (.A(hart_id_i[22]),
    .X(net365));
 sg13g2_buf_1 input367 (.A(hart_id_i[23]),
    .X(net366));
 sg13g2_buf_1 input368 (.A(hart_id_i[24]),
    .X(net367));
 sg13g2_buf_1 input369 (.A(hart_id_i[25]),
    .X(net368));
 sg13g2_buf_1 input370 (.A(hart_id_i[26]),
    .X(net369));
 sg13g2_buf_1 input371 (.A(hart_id_i[27]),
    .X(net370));
 sg13g2_buf_1 input372 (.A(hart_id_i[28]),
    .X(net371));
 sg13g2_buf_1 input373 (.A(hart_id_i[29]),
    .X(net372));
 sg13g2_buf_1 input374 (.A(hart_id_i[2]),
    .X(net373));
 sg13g2_buf_1 input375 (.A(hart_id_i[30]),
    .X(net374));
 sg13g2_buf_1 input376 (.A(hart_id_i[31]),
    .X(net375));
 sg13g2_buf_1 input377 (.A(hart_id_i[3]),
    .X(net376));
 sg13g2_buf_1 input378 (.A(hart_id_i[4]),
    .X(net377));
 sg13g2_buf_1 input379 (.A(hart_id_i[5]),
    .X(net378));
 sg13g2_buf_1 input380 (.A(hart_id_i[6]),
    .X(net379));
 sg13g2_buf_1 input381 (.A(hart_id_i[7]),
    .X(net380));
 sg13g2_buf_1 input382 (.A(hart_id_i[8]),
    .X(net381));
 sg13g2_buf_1 input383 (.A(hart_id_i[9]),
    .X(net382));
 sg13g2_buf_1 input384 (.A(instr_err_i),
    .X(net383));
 sg13g2_buf_1 input385 (.A(instr_gnt_i),
    .X(net384));
 sg13g2_buf_1 input386 (.A(instr_rdata_i[0]),
    .X(net385));
 sg13g2_buf_1 input387 (.A(instr_rdata_i[10]),
    .X(net386));
 sg13g2_buf_1 input388 (.A(instr_rdata_i[11]),
    .X(net387));
 sg13g2_buf_1 input389 (.A(instr_rdata_i[12]),
    .X(net388));
 sg13g2_buf_1 input390 (.A(instr_rdata_i[13]),
    .X(net389));
 sg13g2_buf_1 input391 (.A(instr_rdata_i[14]),
    .X(net390));
 sg13g2_buf_1 input392 (.A(instr_rdata_i[15]),
    .X(net391));
 sg13g2_buf_1 input393 (.A(instr_rdata_i[16]),
    .X(net392));
 sg13g2_buf_1 input394 (.A(instr_rdata_i[17]),
    .X(net393));
 sg13g2_buf_1 input395 (.A(instr_rdata_i[18]),
    .X(net394));
 sg13g2_buf_1 input396 (.A(instr_rdata_i[19]),
    .X(net395));
 sg13g2_buf_1 input397 (.A(instr_rdata_i[1]),
    .X(net396));
 sg13g2_buf_1 input398 (.A(instr_rdata_i[20]),
    .X(net397));
 sg13g2_buf_1 input399 (.A(instr_rdata_i[21]),
    .X(net398));
 sg13g2_buf_1 input400 (.A(instr_rdata_i[22]),
    .X(net399));
 sg13g2_buf_1 input401 (.A(instr_rdata_i[23]),
    .X(net400));
 sg13g2_buf_1 input402 (.A(instr_rdata_i[24]),
    .X(net401));
 sg13g2_buf_1 input403 (.A(instr_rdata_i[25]),
    .X(net402));
 sg13g2_buf_1 input404 (.A(instr_rdata_i[26]),
    .X(net403));
 sg13g2_buf_1 input405 (.A(instr_rdata_i[27]),
    .X(net404));
 sg13g2_buf_1 input406 (.A(instr_rdata_i[28]),
    .X(net405));
 sg13g2_buf_1 input407 (.A(instr_rdata_i[29]),
    .X(net406));
 sg13g2_buf_1 input408 (.A(instr_rdata_i[2]),
    .X(net407));
 sg13g2_buf_1 input409 (.A(instr_rdata_i[30]),
    .X(net408));
 sg13g2_buf_1 input410 (.A(instr_rdata_i[31]),
    .X(net409));
 sg13g2_buf_1 input411 (.A(instr_rdata_i[3]),
    .X(net410));
 sg13g2_buf_1 input412 (.A(instr_rdata_i[4]),
    .X(net411));
 sg13g2_buf_1 input413 (.A(instr_rdata_i[5]),
    .X(net412));
 sg13g2_buf_1 input414 (.A(instr_rdata_i[6]),
    .X(net413));
 sg13g2_buf_1 input415 (.A(instr_rdata_i[7]),
    .X(net414));
 sg13g2_buf_1 input416 (.A(instr_rdata_i[8]),
    .X(net415));
 sg13g2_buf_1 input417 (.A(instr_rdata_i[9]),
    .X(net416));
 sg13g2_buf_1 input418 (.A(instr_rvalid_i),
    .X(net417));
 sg13g2_buf_1 input419 (.A(irq_external_i),
    .X(net418));
 sg13g2_buf_1 input420 (.A(irq_fast_i[0]),
    .X(net419));
 sg13g2_buf_1 input421 (.A(irq_fast_i[10]),
    .X(net420));
 sg13g2_buf_1 input422 (.A(irq_fast_i[11]),
    .X(net421));
 sg13g2_buf_1 input423 (.A(irq_fast_i[12]),
    .X(net422));
 sg13g2_buf_1 input424 (.A(irq_fast_i[13]),
    .X(net423));
 sg13g2_buf_1 input425 (.A(irq_fast_i[14]),
    .X(net424));
 sg13g2_buf_1 input426 (.A(irq_fast_i[1]),
    .X(net425));
 sg13g2_buf_1 input427 (.A(irq_fast_i[2]),
    .X(net426));
 sg13g2_buf_1 input428 (.A(irq_fast_i[3]),
    .X(net427));
 sg13g2_buf_1 input429 (.A(irq_fast_i[4]),
    .X(net428));
 sg13g2_buf_1 input430 (.A(irq_fast_i[5]),
    .X(net429));
 sg13g2_buf_1 input431 (.A(irq_fast_i[6]),
    .X(net430));
 sg13g2_buf_1 input432 (.A(irq_fast_i[7]),
    .X(net431));
 sg13g2_buf_1 input433 (.A(irq_fast_i[8]),
    .X(net432));
 sg13g2_buf_1 input434 (.A(irq_fast_i[9]),
    .X(net433));
 sg13g2_buf_1 input435 (.A(irq_nm_i),
    .X(net434));
 sg13g2_buf_1 input436 (.A(irq_software_i),
    .X(net435));
 sg13g2_buf_1 input437 (.A(irq_timer_i),
    .X(net436));
 sg13g2_buf_1 input438 (.A(rst_ni),
    .X(net437));
 sg13g2_buf_1 input439 (.A(test_en_i),
    .X(net438));
 sg13g2_dfrbpq_1 \load_store_unit_i.addr_last_o[0]$_DFFE_PN0P_  (.RESET_B(net8238),
    .D(_06728_),
    .Q(_01949_),
    .CLK(clknet_leaf_42__06563_));
 sg13g2_dfrbpq_1 \load_store_unit_i.addr_last_o[10]$_DFFE_PN0P_  (.RESET_B(net8238),
    .D(_06727_),
    .Q(_01950_),
    .CLK(clknet_leaf_41__06563_));
 sg13g2_dfrbpq_1 \load_store_unit_i.addr_last_o[11]$_DFFE_PN0P_  (.RESET_B(net8238),
    .D(_06726_),
    .Q(_01951_),
    .CLK(clknet_leaf_41__06563_));
 sg13g2_dfrbpq_1 \load_store_unit_i.addr_last_o[12]$_DFFE_PN0P_  (.RESET_B(net8283),
    .D(_06725_),
    .Q(_01952_),
    .CLK(clknet_leaf_40__06563_));
 sg13g2_dfrbpq_1 \load_store_unit_i.addr_last_o[13]$_DFFE_PN0P_  (.RESET_B(net8283),
    .D(_06724_),
    .Q(_01953_),
    .CLK(clknet_leaf_41__06563_));
 sg13g2_dfrbpq_1 \load_store_unit_i.addr_last_o[14]$_DFFE_PN0P_  (.RESET_B(net8283),
    .D(_06723_),
    .Q(_01954_),
    .CLK(clknet_leaf_41__06563_));
 sg13g2_dfrbpq_1 \load_store_unit_i.addr_last_o[15]$_DFFE_PN0P_  (.RESET_B(net8283),
    .D(_06722_),
    .Q(_01955_),
    .CLK(clknet_leaf_41__06563_));
 sg13g2_dfrbpq_1 \load_store_unit_i.addr_last_o[16]$_DFFE_PN0P_  (.RESET_B(net8243),
    .D(_06721_),
    .Q(_01956_),
    .CLK(clknet_leaf_20__06563_));
 sg13g2_dfrbpq_1 \load_store_unit_i.addr_last_o[17]$_DFFE_PN0P_  (.RESET_B(net8243),
    .D(_06720_),
    .Q(_01957_),
    .CLK(clknet_leaf_20__06563_));
 sg13g2_dfrbpq_1 \load_store_unit_i.addr_last_o[18]$_DFFE_PN0P_  (.RESET_B(net8244),
    .D(_06719_),
    .Q(_01958_),
    .CLK(clknet_leaf_20__06563_));
 sg13g2_dfrbpq_1 \load_store_unit_i.addr_last_o[19]$_DFFE_PN0P_  (.RESET_B(net8245),
    .D(_06718_),
    .Q(_01959_),
    .CLK(clknet_leaf_20__06563_));
 sg13g2_dfrbpq_1 \load_store_unit_i.addr_last_o[1]$_DFFE_PN0P_  (.RESET_B(net8238),
    .D(_06717_),
    .Q(_01960_),
    .CLK(clknet_leaf_42__06563_));
 sg13g2_dfrbpq_1 \load_store_unit_i.addr_last_o[20]$_DFFE_PN0P_  (.RESET_B(net8244),
    .D(_06716_),
    .Q(_01961_),
    .CLK(clknet_leaf_20__06563_));
 sg13g2_dfrbpq_1 \load_store_unit_i.addr_last_o[21]$_DFFE_PN0P_  (.RESET_B(net8244),
    .D(_06715_),
    .Q(_01962_),
    .CLK(clknet_leaf_20__06563_));
 sg13g2_dfrbpq_1 \load_store_unit_i.addr_last_o[22]$_DFFE_PN0P_  (.RESET_B(net8244),
    .D(_06714_),
    .Q(_01963_),
    .CLK(clknet_leaf_20__06563_));
 sg13g2_dfrbpq_1 \load_store_unit_i.addr_last_o[23]$_DFFE_PN0P_  (.RESET_B(net8244),
    .D(_06713_),
    .Q(_01964_),
    .CLK(clknet_leaf_20__06563_));
 sg13g2_dfrbpq_1 \load_store_unit_i.addr_last_o[24]$_DFFE_PN0P_  (.RESET_B(net8244),
    .D(_06712_),
    .Q(_01965_),
    .CLK(clknet_leaf_20__06563_));
 sg13g2_dfrbpq_1 \load_store_unit_i.addr_last_o[25]$_DFFE_PN0P_  (.RESET_B(net8243),
    .D(_06711_),
    .Q(_01966_),
    .CLK(clknet_leaf_20__06563_));
 sg13g2_dfrbpq_1 \load_store_unit_i.addr_last_o[26]$_DFFE_PN0P_  (.RESET_B(net8244),
    .D(_06710_),
    .Q(_01967_),
    .CLK(clknet_leaf_20__06563_));
 sg13g2_dfrbpq_1 \load_store_unit_i.addr_last_o[27]$_DFFE_PN0P_  (.RESET_B(net8245),
    .D(_06709_),
    .Q(_01968_),
    .CLK(clknet_leaf_20__06563_));
 sg13g2_dfrbpq_1 \load_store_unit_i.addr_last_o[28]$_DFFE_PN0P_  (.RESET_B(net8245),
    .D(_06708_),
    .Q(_01969_),
    .CLK(clknet_leaf_20__06563_));
 sg13g2_dfrbpq_1 \load_store_unit_i.addr_last_o[29]$_DFFE_PN0P_  (.RESET_B(net8244),
    .D(_06707_),
    .Q(_01970_),
    .CLK(clknet_leaf_20__06563_));
 sg13g2_dfrbpq_1 \load_store_unit_i.addr_last_o[2]$_DFFE_PN0P_  (.RESET_B(net8238),
    .D(_06706_),
    .Q(_01971_),
    .CLK(clknet_leaf_42__06563_));
 sg13g2_dfrbpq_1 \load_store_unit_i.addr_last_o[30]$_DFFE_PN0P_  (.RESET_B(net8243),
    .D(_06705_),
    .Q(_01972_),
    .CLK(clknet_leaf_20__06563_));
 sg13g2_dfrbpq_1 \load_store_unit_i.addr_last_o[31]$_DFFE_PN0P_  (.RESET_B(net8243),
    .D(_06704_),
    .Q(_01973_),
    .CLK(clknet_leaf_41__06563_));
 sg13g2_dfrbpq_1 \load_store_unit_i.addr_last_o[3]$_DFFE_PN0P_  (.RESET_B(net8238),
    .D(_06703_),
    .Q(_01974_),
    .CLK(clknet_leaf_42__06563_));
 sg13g2_dfrbpq_1 \load_store_unit_i.addr_last_o[4]$_DFFE_PN0P_  (.RESET_B(net8283),
    .D(_06702_),
    .Q(_01975_),
    .CLK(clknet_leaf_41__06563_));
 sg13g2_dfrbpq_1 \load_store_unit_i.addr_last_o[5]$_DFFE_PN0P_  (.RESET_B(net8243),
    .D(_06701_),
    .Q(_01976_),
    .CLK(clknet_leaf_41__06563_));
 sg13g2_dfrbpq_1 \load_store_unit_i.addr_last_o[6]$_DFFE_PN0P_  (.RESET_B(net8252),
    .D(_06700_),
    .Q(_01977_),
    .CLK(clknet_leaf_41__06563_));
 sg13g2_dfrbpq_1 \load_store_unit_i.addr_last_o[7]$_DFFE_PN0P_  (.RESET_B(net8243),
    .D(_06699_),
    .Q(_01978_),
    .CLK(clknet_leaf_41__06563_));
 sg13g2_dfrbpq_1 \load_store_unit_i.addr_last_o[8]$_DFFE_PN0P_  (.RESET_B(net8243),
    .D(_06698_),
    .Q(_01979_),
    .CLK(clknet_leaf_41__06563_));
 sg13g2_dfrbpq_1 \load_store_unit_i.addr_last_o[9]$_DFFE_PN0P_  (.RESET_B(net8257),
    .D(_06697_),
    .Q(_01980_),
    .CLK(clknet_leaf_40__06563_));
 sg13g2_dfrbpq_1 \load_store_unit_i.data_sign_ext_q$_DFFE_PN0P_  (.RESET_B(net8230),
    .D(_06689_),
    .Q(\load_store_unit_i.data_sign_ext_q ),
    .CLK(clknet_leaf_2__06563_));
 sg13g2_dfrbpq_1 \load_store_unit_i.data_type_q[0]$_DFF_PN1_  (.RESET_B(net8230),
    .D(_06687_),
    .Q(_00007_),
    .CLK(clknet_leaf_2__06563_));
 sg13g2_dfrbpq_1 \load_store_unit_i.data_type_q[1]$_DFF_PN0_  (.RESET_B(net8230),
    .D(_06685_),
    .Q(_01981_),
    .CLK(clknet_leaf_2__06563_));
 sg13g2_dfrbpq_1 \load_store_unit_i.data_type_q[2]$_DFF_PN0_  (.RESET_B(net8231),
    .D(_06682_),
    .Q(_01982_),
    .CLK(clknet_leaf_2__06563_));
 sg13g2_dfrbpq_1 \load_store_unit_i.data_we_q$_DFFE_PN0P_  (.RESET_B(net8240),
    .D(_06680_),
    .Q(\load_store_unit_i.data_we_q ),
    .CLK(clknet_leaf_42__06563_));
 sg13g2_dfrbpq_1 \load_store_unit_i.handle_misaligned_q$_DFFE_PN0P_  (.RESET_B(net8240),
    .D(_06679_),
    .Q(\load_store_unit_i.handle_misaligned_q ),
    .CLK(clknet_leaf_42__06563_));
 sg13g2_dfrbpq_1 \load_store_unit_i.ls_fsm_cs[0]$_DFFE_PN0P_  (.RESET_B(net8240),
    .D(_06671_),
    .Q(_01983_),
    .CLK(clknet_leaf_44__06563_));
 sg13g2_dfrbpq_1 \load_store_unit_i.ls_fsm_cs[1]$_DFFE_PN0P_  (.RESET_B(net8240),
    .D(_06668_),
    .Q(_01984_),
    .CLK(clknet_leaf_42__06563_));
 sg13g2_dfrbpq_1 \load_store_unit_i.ls_fsm_cs[2]$_DFFE_PN0P_  (.RESET_B(net8240),
    .D(_06656_),
    .Q(_01985_),
    .CLK(clknet_leaf_42__06563_));
 sg13g2_dfrbpq_1 \load_store_unit_i.lsu_err_q$_DFFE_PN0P_  (.RESET_B(net8240),
    .D(_06654_),
    .Q(\load_store_unit_i.lsu_err_q ),
    .CLK(clknet_leaf_45__06563_));
 sg13g2_dfrbpq_1 \load_store_unit_i.rdata_offset_q[0]$_DFFE_PN0P_  (.RESET_B(net8230),
    .D(_06650_),
    .Q(_01986_),
    .CLK(clknet_leaf_2__06563_));
 sg13g2_dfrbpq_1 \load_store_unit_i.rdata_offset_q[1]$_DFFE_PN0P_  (.RESET_B(net8230),
    .D(_06649_),
    .Q(_01987_),
    .CLK(clknet_leaf_2__06563_));
 sg13g2_dfrbpq_1 \load_store_unit_i.rdata_q[10]$_DFFE_PN0P_  (.RESET_B(net8037),
    .D(_06596_),
    .Q(_01988_),
    .CLK(clknet_leaf_3__06563_));
 sg13g2_dfrbpq_1 \load_store_unit_i.rdata_q[11]$_DFFE_PN0P_  (.RESET_B(net8036),
    .D(_06595_),
    .Q(_01989_),
    .CLK(clknet_leaf_4__06563_));
 sg13g2_dfrbpq_1 \load_store_unit_i.rdata_q[12]$_DFFE_PN0P_  (.RESET_B(net8036),
    .D(_06594_),
    .Q(_01990_),
    .CLK(clknet_leaf_4__06563_));
 sg13g2_dfrbpq_1 \load_store_unit_i.rdata_q[13]$_DFFE_PN0P_  (.RESET_B(net8231),
    .D(_06593_),
    .Q(_01991_),
    .CLK(clknet_leaf_3__06563_));
 sg13g2_dfrbpq_1 \load_store_unit_i.rdata_q[14]$_DFFE_PN0P_  (.RESET_B(net8036),
    .D(_06591_),
    .Q(_01992_),
    .CLK(clknet_leaf_3__06563_));
 sg13g2_dfrbpq_1 \load_store_unit_i.rdata_q[15]$_DFFE_PN0P_  (.RESET_B(net8037),
    .D(_06590_),
    .Q(_01993_),
    .CLK(clknet_leaf_3__06563_));
 sg13g2_dfrbpq_1 \load_store_unit_i.rdata_q[16]$_DFFE_PN0P_  (.RESET_B(net8284),
    .D(_06589_),
    .Q(_01994_),
    .CLK(clknet_leaf_2__06563_));
 sg13g2_dfrbpq_1 \load_store_unit_i.rdata_q[17]$_DFFE_PN0P_  (.RESET_B(net8037),
    .D(_06588_),
    .Q(_01995_),
    .CLK(clknet_leaf_3__06563_));
 sg13g2_dfrbpq_1 \load_store_unit_i.rdata_q[18]$_DFFE_PN0P_  (.RESET_B(net8037),
    .D(_06587_),
    .Q(_01996_),
    .CLK(clknet_leaf_3__06563_));
 sg13g2_dfrbpq_1 \load_store_unit_i.rdata_q[19]$_DFFE_PN0P_  (.RESET_B(net8036),
    .D(_06586_),
    .Q(_01997_),
    .CLK(clknet_leaf_4__06563_));
 sg13g2_dfrbpq_1 \load_store_unit_i.rdata_q[20]$_DFFE_PN0P_  (.RESET_B(net8053),
    .D(_06584_),
    .Q(_01998_),
    .CLK(clknet_leaf_4__06563_));
 sg13g2_dfrbpq_1 \load_store_unit_i.rdata_q[21]$_DFFE_PN0P_  (.RESET_B(net8230),
    .D(_06583_),
    .Q(_01999_),
    .CLK(clknet_leaf_2__06563_));
 sg13g2_dfrbpq_1 \load_store_unit_i.rdata_q[22]$_DFFE_PN0P_  (.RESET_B(net8036),
    .D(_06582_),
    .Q(_02000_),
    .CLK(clknet_leaf_3__06563_));
 sg13g2_dfrbpq_1 \load_store_unit_i.rdata_q[23]$_DFFE_PN0P_  (.RESET_B(net8037),
    .D(_06581_),
    .Q(_02001_),
    .CLK(clknet_leaf_3__06563_));
 sg13g2_dfrbpq_1 \load_store_unit_i.rdata_q[24]$_DFFE_PN0P_  (.RESET_B(net8284),
    .D(_06580_),
    .Q(_02002_),
    .CLK(clknet_leaf_2__06563_));
 sg13g2_dfrbpq_1 \load_store_unit_i.rdata_q[25]$_DFFE_PN0P_  (.RESET_B(net8037),
    .D(_06579_),
    .Q(_02003_),
    .CLK(clknet_leaf_3__06563_));
 sg13g2_dfrbpq_1 \load_store_unit_i.rdata_q[26]$_DFFE_PN0P_  (.RESET_B(net8037),
    .D(_06578_),
    .Q(_02004_),
    .CLK(clknet_leaf_3__06563_));
 sg13g2_dfrbpq_1 \load_store_unit_i.rdata_q[27]$_DFFE_PN0P_  (.RESET_B(net8053),
    .D(_06577_),
    .Q(_02005_),
    .CLK(clknet_leaf_4__06563_));
 sg13g2_dfrbpq_1 \load_store_unit_i.rdata_q[28]$_DFFE_PN0P_  (.RESET_B(net8053),
    .D(_06576_),
    .Q(_02006_),
    .CLK(clknet_leaf_4__06563_));
 sg13g2_dfrbpq_1 \load_store_unit_i.rdata_q[29]$_DFFE_PN0P_  (.RESET_B(net8230),
    .D(_06575_),
    .Q(_02007_),
    .CLK(clknet_leaf_2__06563_));
 sg13g2_dfrbpq_1 \load_store_unit_i.rdata_q[30]$_DFFE_PN0P_  (.RESET_B(net8036),
    .D(_06573_),
    .Q(_02008_),
    .CLK(clknet_leaf_3__06563_));
 sg13g2_dfrbpq_1 \load_store_unit_i.rdata_q[31]$_DFFE_PN0P_  (.RESET_B(net8037),
    .D(_06572_),
    .Q(_02009_),
    .CLK(clknet_leaf_3__06563_));
 sg13g2_dfrbpq_1 \load_store_unit_i.rdata_q[8]$_DFFE_PN0P_  (.RESET_B(net8230),
    .D(_06571_),
    .Q(_02010_),
    .CLK(clknet_leaf_2__06563_));
 sg13g2_dfrbpq_1 \load_store_unit_i.rdata_q[9]$_DFFE_PN0P_  (.RESET_B(net8036),
    .D(_06570_),
    .Q(_02011_),
    .CLK(clknet_leaf_3__06563_));
 sg13g2_buf_1 output440 (.A(net439),
    .X(core_sleep_o));
 sg13g2_buf_1 output441 (.A(net6622),
    .X(data_addr_o[10]));
 sg13g2_buf_1 output442 (.A(net6621),
    .X(data_addr_o[11]));
 sg13g2_buf_1 output443 (.A(net6601),
    .X(data_addr_o[12]));
 sg13g2_buf_1 output444 (.A(net443),
    .X(data_addr_o[13]));
 sg13g2_buf_1 output445 (.A(net6615),
    .X(data_addr_o[14]));
 sg13g2_buf_1 output446 (.A(net6613),
    .X(data_addr_o[15]));
 sg13g2_buf_1 output447 (.A(net6610),
    .X(data_addr_o[16]));
 sg13g2_buf_1 output448 (.A(net6609),
    .X(data_addr_o[17]));
 sg13g2_buf_1 output449 (.A(net6608),
    .X(data_addr_o[18]));
 sg13g2_buf_1 output450 (.A(net6607),
    .X(data_addr_o[19]));
 sg13g2_buf_1 output451 (.A(net6586),
    .X(data_addr_o[20]));
 sg13g2_buf_1 output452 (.A(net6584),
    .X(data_addr_o[21]));
 sg13g2_buf_1 output453 (.A(net6605),
    .X(data_addr_o[22]));
 sg13g2_buf_1 output454 (.A(net6603),
    .X(data_addr_o[23]));
 sg13g2_buf_1 output455 (.A(net6582),
    .X(data_addr_o[24]));
 sg13g2_buf_1 output456 (.A(net6579),
    .X(data_addr_o[25]));
 sg13g2_buf_1 output457 (.A(net6576),
    .X(data_addr_o[26]));
 sg13g2_buf_1 output458 (.A(net6575),
    .X(data_addr_o[27]));
 sg13g2_buf_1 output459 (.A(net6573),
    .X(data_addr_o[28]));
 sg13g2_buf_1 output460 (.A(net6571),
    .X(data_addr_o[29]));
 sg13g2_buf_1 output461 (.A(net6640),
    .X(data_addr_o[2]));
 sg13g2_buf_1 output462 (.A(net6570),
    .X(data_addr_o[30]));
 sg13g2_buf_1 output463 (.A(net6567),
    .X(data_addr_o[31]));
 sg13g2_buf_1 output464 (.A(net6639),
    .X(data_addr_o[3]));
 sg13g2_buf_1 output465 (.A(net464),
    .X(data_addr_o[4]));
 sg13g2_buf_1 output466 (.A(net6637),
    .X(data_addr_o[5]));
 sg13g2_buf_1 output467 (.A(net6628),
    .X(data_addr_o[6]));
 sg13g2_buf_1 output468 (.A(net467),
    .X(data_addr_o[7]));
 sg13g2_buf_1 output469 (.A(net6626),
    .X(data_addr_o[8]));
 sg13g2_buf_1 output470 (.A(net6624),
    .X(data_addr_o[9]));
 sg13g2_buf_1 output471 (.A(net470),
    .X(data_be_o[0]));
 sg13g2_buf_1 output472 (.A(net471),
    .X(data_be_o[1]));
 sg13g2_buf_1 output473 (.A(net472),
    .X(data_be_o[2]));
 sg13g2_buf_1 output474 (.A(net473),
    .X(data_be_o[3]));
 sg13g2_buf_1 output475 (.A(net474),
    .X(data_req_o));
 sg13g2_buf_1 output476 (.A(net475),
    .X(data_wdata_o[0]));
 sg13g2_buf_1 output477 (.A(net476),
    .X(data_wdata_o[10]));
 sg13g2_buf_1 output478 (.A(net477),
    .X(data_wdata_o[11]));
 sg13g2_buf_1 output479 (.A(net478),
    .X(data_wdata_o[12]));
 sg13g2_buf_1 output480 (.A(net479),
    .X(data_wdata_o[13]));
 sg13g2_buf_1 output481 (.A(net480),
    .X(data_wdata_o[14]));
 sg13g2_buf_1 output482 (.A(net481),
    .X(data_wdata_o[15]));
 sg13g2_buf_1 output483 (.A(net482),
    .X(data_wdata_o[16]));
 sg13g2_buf_1 output484 (.A(net483),
    .X(data_wdata_o[17]));
 sg13g2_buf_1 output485 (.A(net484),
    .X(data_wdata_o[18]));
 sg13g2_buf_1 output486 (.A(net485),
    .X(data_wdata_o[19]));
 sg13g2_buf_1 output487 (.A(net486),
    .X(data_wdata_o[1]));
 sg13g2_buf_1 output488 (.A(net487),
    .X(data_wdata_o[20]));
 sg13g2_buf_1 output489 (.A(net488),
    .X(data_wdata_o[21]));
 sg13g2_buf_1 output490 (.A(net489),
    .X(data_wdata_o[22]));
 sg13g2_buf_1 output491 (.A(net490),
    .X(data_wdata_o[23]));
 sg13g2_buf_1 output492 (.A(net491),
    .X(data_wdata_o[24]));
 sg13g2_buf_1 output493 (.A(net492),
    .X(data_wdata_o[25]));
 sg13g2_buf_1 output494 (.A(net493),
    .X(data_wdata_o[26]));
 sg13g2_buf_1 output495 (.A(net494),
    .X(data_wdata_o[27]));
 sg13g2_buf_1 output496 (.A(net495),
    .X(data_wdata_o[28]));
 sg13g2_buf_1 output497 (.A(net496),
    .X(data_wdata_o[29]));
 sg13g2_buf_1 output498 (.A(net497),
    .X(data_wdata_o[2]));
 sg13g2_buf_1 output499 (.A(net498),
    .X(data_wdata_o[30]));
 sg13g2_buf_1 output500 (.A(net499),
    .X(data_wdata_o[31]));
 sg13g2_buf_1 output501 (.A(net500),
    .X(data_wdata_o[3]));
 sg13g2_buf_1 output502 (.A(net501),
    .X(data_wdata_o[4]));
 sg13g2_buf_1 output503 (.A(net502),
    .X(data_wdata_o[5]));
 sg13g2_buf_1 output504 (.A(net503),
    .X(data_wdata_o[6]));
 sg13g2_buf_1 output505 (.A(net504),
    .X(data_wdata_o[7]));
 sg13g2_buf_1 output506 (.A(net505),
    .X(data_wdata_o[8]));
 sg13g2_buf_1 output507 (.A(net506),
    .X(data_wdata_o[9]));
 sg13g2_buf_1 output508 (.A(net507),
    .X(data_we_o));
 sg13g2_buf_1 output509 (.A(net508),
    .X(instr_addr_o[10]));
 sg13g2_buf_1 output510 (.A(net509),
    .X(instr_addr_o[11]));
 sg13g2_buf_1 output511 (.A(net510),
    .X(instr_addr_o[12]));
 sg13g2_buf_1 output512 (.A(net511),
    .X(instr_addr_o[13]));
 sg13g2_buf_1 output513 (.A(net512),
    .X(instr_addr_o[14]));
 sg13g2_buf_1 output514 (.A(net513),
    .X(instr_addr_o[15]));
 sg13g2_buf_1 output515 (.A(net514),
    .X(instr_addr_o[16]));
 sg13g2_buf_1 output516 (.A(net515),
    .X(instr_addr_o[17]));
 sg13g2_buf_1 output517 (.A(net516),
    .X(instr_addr_o[18]));
 sg13g2_buf_1 output518 (.A(net517),
    .X(instr_addr_o[19]));
 sg13g2_buf_1 output519 (.A(net518),
    .X(instr_addr_o[20]));
 sg13g2_buf_1 output520 (.A(net519),
    .X(instr_addr_o[21]));
 sg13g2_buf_1 output521 (.A(net520),
    .X(instr_addr_o[22]));
 sg13g2_buf_1 output522 (.A(net521),
    .X(instr_addr_o[23]));
 sg13g2_buf_1 output523 (.A(net522),
    .X(instr_addr_o[24]));
 sg13g2_buf_1 output524 (.A(net523),
    .X(instr_addr_o[25]));
 sg13g2_buf_1 output525 (.A(net524),
    .X(instr_addr_o[26]));
 sg13g2_buf_1 output526 (.A(net525),
    .X(instr_addr_o[27]));
 sg13g2_buf_1 output527 (.A(net526),
    .X(instr_addr_o[28]));
 sg13g2_buf_1 output528 (.A(net527),
    .X(instr_addr_o[29]));
 sg13g2_buf_1 output529 (.A(net528),
    .X(instr_addr_o[2]));
 sg13g2_buf_1 output530 (.A(net529),
    .X(instr_addr_o[30]));
 sg13g2_buf_1 output531 (.A(net530),
    .X(instr_addr_o[31]));
 sg13g2_buf_1 output532 (.A(net531),
    .X(instr_addr_o[3]));
 sg13g2_buf_1 output533 (.A(net532),
    .X(instr_addr_o[4]));
 sg13g2_buf_1 output534 (.A(net533),
    .X(instr_addr_o[5]));
 sg13g2_buf_1 output535 (.A(net534),
    .X(instr_addr_o[6]));
 sg13g2_buf_1 output536 (.A(net535),
    .X(instr_addr_o[7]));
 sg13g2_buf_1 output537 (.A(net536),
    .X(instr_addr_o[8]));
 sg13g2_buf_1 output538 (.A(net537),
    .X(instr_addr_o[9]));
 sg13g2_buf_1 output539 (.A(net538),
    .X(instr_req_o));
 sg13g2_buf_1 place5762 (.A(net5764),
    .X(net5761));
 sg13g2_buf_1 place5763 (.A(net5764),
    .X(net5762));
 sg13g2_buf_1 place5764 (.A(net5764),
    .X(net5763));
 sg13g2_buf_1 place5765 (.A(_14609_),
    .X(net5764));
 sg13g2_buf_1 place5766 (.A(net5771),
    .X(net5765));
 sg13g2_buf_1 place5767 (.A(net5771),
    .X(net5766));
 sg13g2_buf_2 place5768 (.A(net5771),
    .X(net5767));
 sg13g2_buf_1 place5769 (.A(net5771),
    .X(net5768));
 sg13g2_buf_1 place5770 (.A(net5771),
    .X(net5769));
 sg13g2_buf_2 place5771 (.A(net5771),
    .X(net5770));
 sg13g2_buf_8 place5772 (.A(_14609_),
    .X(net5771));
 sg13g2_buf_1 place5773 (.A(net5777),
    .X(net5772));
 sg13g2_buf_4 place5774 (.X(net5773),
    .A(net5777));
 sg13g2_buf_4 place5775 (.X(net5774),
    .A(net5777));
 sg13g2_buf_4 place5776 (.X(net5775),
    .A(net5777));
 sg13g2_buf_1 place5777 (.A(net5777),
    .X(net5776));
 sg13g2_buf_4 place5778 (.X(net5777),
    .A(_10724_));
 sg13g2_buf_4 place5779 (.X(net5778),
    .A(net5784));
 sg13g2_buf_1 place5780 (.A(net5784),
    .X(net5779));
 sg13g2_buf_1 place5781 (.A(net5784),
    .X(net5780));
 sg13g2_buf_8 place5782 (.A(net5784),
    .X(net5781));
 sg13g2_buf_1 place5783 (.A(net5784),
    .X(net5782));
 sg13g2_buf_8 place5784 (.A(net5784),
    .X(net5783));
 sg13g2_buf_4 place5785 (.X(net5784),
    .A(_10456_));
 sg13g2_buf_1 place5786 (.A(net5791),
    .X(net5785));
 sg13g2_buf_8 place5787 (.A(net5791),
    .X(net5786));
 sg13g2_buf_2 place5788 (.A(net5791),
    .X(net5787));
 sg13g2_buf_2 place5789 (.A(net5791),
    .X(net5788));
 sg13g2_buf_4 place5790 (.X(net5789),
    .A(net5791));
 sg13g2_buf_16 place5791 (.X(net5790),
    .A(net5791));
 sg13g2_buf_8 place5792 (.A(_10373_),
    .X(net5791));
 sg13g2_buf_1 place5793 (.A(_10308_),
    .X(net5792));
 sg13g2_buf_1 place5794 (.A(net5797),
    .X(net5793));
 sg13g2_buf_4 place5795 (.X(net5794),
    .A(net5797));
 sg13g2_buf_4 place5796 (.X(net5795),
    .A(net5797));
 sg13g2_buf_8 place5797 (.A(net5797),
    .X(net5796));
 sg13g2_buf_4 place5798 (.X(net5797),
    .A(_10308_));
 sg13g2_buf_1 place5799 (.A(net5803),
    .X(net5798));
 sg13g2_buf_1 place5800 (.A(net5803),
    .X(net5799));
 sg13g2_buf_1 place5801 (.A(net5802),
    .X(net5800));
 sg13g2_buf_4 place5802 (.X(net5801),
    .A(net5802));
 sg13g2_buf_8 place5803 (.A(net5803),
    .X(net5802));
 sg13g2_buf_8 place5804 (.A(_10269_),
    .X(net5803));
 sg13g2_buf_8 place5805 (.A(net5809),
    .X(net5804));
 sg13g2_buf_2 place5806 (.A(net5809),
    .X(net5805));
 sg13g2_buf_2 place5807 (.A(net5809),
    .X(net5806));
 sg13g2_buf_8 place5808 (.A(net5809),
    .X(net5807));
 sg13g2_buf_8 place5809 (.A(net5809),
    .X(net5808));
 sg13g2_buf_8 place5810 (.A(_10204_),
    .X(net5809));
 sg13g2_buf_1 place5811 (.A(net5819),
    .X(net5810));
 sg13g2_buf_1 place5812 (.A(net5812),
    .X(net5811));
 sg13g2_buf_1 place5813 (.A(net5819),
    .X(net5812));
 sg13g2_buf_1 place5814 (.A(net5819),
    .X(net5813));
 sg13g2_buf_1 place5815 (.A(net5819),
    .X(net5814));
 sg13g2_buf_1 place5816 (.A(net5819),
    .X(net5815));
 sg13g2_buf_1 place5817 (.A(net5819),
    .X(net5816));
 sg13g2_buf_1 place5818 (.A(net5818),
    .X(net5817));
 sg13g2_buf_1 place5819 (.A(net5819),
    .X(net5818));
 sg13g2_buf_2 place5820 (.A(_08077_),
    .X(net5819));
 sg13g2_buf_1 place5821 (.A(net5822),
    .X(net5820));
 sg13g2_buf_1 place5822 (.A(net5822),
    .X(net5821));
 sg13g2_buf_1 place5823 (.A(net5827),
    .X(net5822));
 sg13g2_buf_1 place5824 (.A(net5827),
    .X(net5823));
 sg13g2_buf_2 place5825 (.A(net5827),
    .X(net5824));
 sg13g2_buf_2 place5826 (.A(net5826),
    .X(net5825));
 sg13g2_buf_1 place5827 (.A(net5827),
    .X(net5826));
 sg13g2_buf_2 place5828 (.A(_14572_),
    .X(net5827));
 sg13g2_buf_1 place5829 (.A(net5829),
    .X(net5828));
 sg13g2_buf_1 place5830 (.A(net5832),
    .X(net5829));
 sg13g2_buf_1 place5831 (.A(net5832),
    .X(net5830));
 sg13g2_buf_1 place5832 (.A(net5832),
    .X(net5831));
 sg13g2_buf_1 place5833 (.A(_14572_),
    .X(net5832));
 sg13g2_buf_2 place5834 (.A(net5837),
    .X(net5833));
 sg13g2_buf_2 place5835 (.A(net5837),
    .X(net5834));
 sg13g2_buf_4 place5836 (.X(net5835),
    .A(net5837));
 sg13g2_buf_2 place5837 (.A(net5837),
    .X(net5836));
 sg13g2_buf_4 place5838 (.X(net5837),
    .A(_10572_));
 sg13g2_buf_8 place5839 (.A(net5843),
    .X(net5838));
 sg13g2_buf_8 place5840 (.A(net5843),
    .X(net5839));
 sg13g2_buf_8 place5841 (.A(net5843),
    .X(net5840));
 sg13g2_buf_1 place5842 (.A(net5843),
    .X(net5841));
 sg13g2_buf_8 place5843 (.A(net5843),
    .X(net5842));
 sg13g2_buf_8 place5844 (.A(_10532_),
    .X(net5843));
 sg13g2_buf_8 place5845 (.A(_10450_),
    .X(net5844));
 sg13g2_buf_4 place5846 (.X(net5845),
    .A(_10369_));
 sg13g2_buf_4 place5847 (.X(net5846),
    .A(_10301_));
 sg13g2_buf_4 place5848 (.X(net5847),
    .A(net5851));
 sg13g2_buf_4 place5849 (.X(net5848),
    .A(net5851));
 sg13g2_buf_2 place5850 (.A(net5851),
    .X(net5849));
 sg13g2_buf_4 place5851 (.X(net5850),
    .A(net5851));
 sg13g2_buf_8 place5852 (.A(_10236_),
    .X(net5851));
 sg13g2_buf_8 place5853 (.A(_10201_),
    .X(net5852));
 sg13g2_buf_1 place5854 (.A(net5858),
    .X(net5853));
 sg13g2_buf_2 place5855 (.A(net5858),
    .X(net5854));
 sg13g2_buf_2 place5856 (.A(net5858),
    .X(net5855));
 sg13g2_buf_1 place5857 (.A(net5858),
    .X(net5856));
 sg13g2_buf_2 place5858 (.A(net5858),
    .X(net5857));
 sg13g2_buf_8 place5859 (.A(_10159_),
    .X(net5858));
 sg13g2_buf_4 place5860 (.X(net5859),
    .A(net5863));
 sg13g2_buf_1 place5861 (.A(net5863),
    .X(net5860));
 sg13g2_buf_1 place5862 (.A(net5863),
    .X(net5861));
 sg13g2_buf_1 place5863 (.A(net5863),
    .X(net5862));
 sg13g2_buf_8 place5864 (.A(_10132_),
    .X(net5863));
 sg13g2_buf_1 place5865 (.A(_10088_),
    .X(net5864));
 sg13g2_buf_1 place5866 (.A(_10088_),
    .X(net5865));
 sg13g2_buf_1 place5867 (.A(_10088_),
    .X(net5866));
 sg13g2_buf_1 place5868 (.A(_10088_),
    .X(net5867));
 sg13g2_buf_1 place5869 (.A(_08396_),
    .X(net5868));
 sg13g2_buf_1 place5870 (.A(_08122_),
    .X(net5869));
 sg13g2_buf_1 place5871 (.A(_08122_),
    .X(net5870));
 sg13g2_buf_1 place5872 (.A(_08122_),
    .X(net5871));
 sg13g2_buf_1 place5873 (.A(net5880),
    .X(net5872));
 sg13g2_buf_1 place5874 (.A(net5880),
    .X(net5873));
 sg13g2_buf_1 place5875 (.A(net5880),
    .X(net5874));
 sg13g2_buf_1 place5876 (.A(net5880),
    .X(net5875));
 sg13g2_buf_1 place5877 (.A(net5880),
    .X(net5876));
 sg13g2_buf_1 place5878 (.A(net5880),
    .X(net5877));
 sg13g2_buf_1 place5879 (.A(net5880),
    .X(net5878));
 sg13g2_buf_1 place5880 (.A(net5880),
    .X(net5879));
 sg13g2_buf_4 place5881 (.X(net5880),
    .A(_08122_));
 sg13g2_buf_1 place5882 (.A(_14564_),
    .X(net5881));
 sg13g2_buf_2 place5883 (.A(net5886),
    .X(net5882));
 sg13g2_buf_2 place5884 (.A(net5886),
    .X(net5883));
 sg13g2_buf_1 place5885 (.A(net5886),
    .X(net5884));
 sg13g2_buf_2 place5886 (.A(net5886),
    .X(net5885));
 sg13g2_buf_4 place5887 (.X(net5886),
    .A(_10758_));
 sg13g2_buf_2 place5888 (.A(_10710_),
    .X(net5887));
 sg13g2_buf_2 place5889 (.A(net5894),
    .X(net5888));
 sg13g2_buf_2 place5890 (.A(net5894),
    .X(net5889));
 sg13g2_buf_1 place5891 (.A(net5894),
    .X(net5890));
 sg13g2_buf_4 place5892 (.X(net5891),
    .A(net5894));
 sg13g2_buf_1 place5893 (.A(net5894),
    .X(net5892));
 sg13g2_buf_16 place5894 (.X(net5893),
    .A(net5894));
 sg13g2_buf_8 place5895 (.A(_10693_),
    .X(net5894));
 sg13g2_buf_1 place5896 (.A(net5899),
    .X(net5895));
 sg13g2_buf_4 place5897 (.X(net5896),
    .A(net5899));
 sg13g2_buf_4 place5898 (.X(net5897),
    .A(net5899));
 sg13g2_buf_1 place5899 (.A(net5899),
    .X(net5898));
 sg13g2_buf_4 place5900 (.X(net5899),
    .A(_10652_));
 sg13g2_buf_4 place5901 (.X(net5900),
    .A(net5904));
 sg13g2_buf_16 place5902 (.X(net5901),
    .A(net5904));
 sg13g2_buf_4 place5903 (.X(net5902),
    .A(net5904));
 sg13g2_buf_1 place5904 (.A(net5904),
    .X(net5903));
 sg13g2_buf_8 place5905 (.A(_10615_),
    .X(net5904));
 sg13g2_buf_2 place5906 (.A(_10567_),
    .X(net5905));
 sg13g2_buf_4 place5907 (.X(net5906),
    .A(_10527_));
 sg13g2_buf_1 place5908 (.A(net5911),
    .X(net5907));
 sg13g2_buf_1 place5909 (.A(net5911),
    .X(net5908));
 sg13g2_buf_1 place5910 (.A(net5911),
    .X(net5909));
 sg13g2_buf_1 place5911 (.A(net5911),
    .X(net5910));
 sg13g2_buf_2 place5912 (.A(_10488_),
    .X(net5911));
 sg13g2_buf_1 place5913 (.A(net5916),
    .X(net5912));
 sg13g2_buf_1 place5914 (.A(net5916),
    .X(net5913));
 sg13g2_buf_1 place5915 (.A(net5916),
    .X(net5914));
 sg13g2_buf_1 place5916 (.A(net5916),
    .X(net5915));
 sg13g2_buf_8 place5917 (.A(_10411_),
    .X(net5916));
 sg13g2_buf_2 place5918 (.A(net5921),
    .X(net5917));
 sg13g2_buf_1 place5919 (.A(net5921),
    .X(net5918));
 sg13g2_buf_1 place5920 (.A(net5921),
    .X(net5919));
 sg13g2_buf_1 place5921 (.A(net5921),
    .X(net5920));
 sg13g2_buf_8 place5922 (.A(_10337_),
    .X(net5921));
 sg13g2_buf_1 place5923 (.A(_07045_),
    .X(net5922));
 sg13g2_buf_1 place5924 (.A(_00101_),
    .X(net5923));
 sg13g2_buf_2 place5925 (.A(_00096_),
    .X(net5924));
 sg13g2_buf_1 place5926 (.A(net5929),
    .X(net5925));
 sg13g2_buf_4 place5927 (.X(net5926),
    .A(net5929));
 sg13g2_buf_1 place5928 (.A(net5929),
    .X(net5927));
 sg13g2_buf_1 place5929 (.A(net5929),
    .X(net5928));
 sg13g2_buf_8 place5930 (.A(_10790_),
    .X(net5929));
 sg13g2_buf_4 place5931 (.X(net5930),
    .A(_10692_));
 sg13g2_buf_2 place5932 (.A(_10647_),
    .X(net5931));
 sg13g2_buf_4 place5933 (.X(net5932),
    .A(_10609_));
 sg13g2_buf_1 place5934 (.A(_08956_),
    .X(net5933));
 sg13g2_buf_1 place5935 (.A(net5935),
    .X(net5934));
 sg13g2_buf_1 place5936 (.A(net5939),
    .X(net5935));
 sg13g2_buf_1 place5937 (.A(net5937),
    .X(net5936));
 sg13g2_buf_2 place5938 (.A(net5939),
    .X(net5937));
 sg13g2_buf_1 place5939 (.A(net5939),
    .X(net5938));
 sg13g2_buf_2 place5940 (.A(net5940),
    .X(net5939));
 sg13g2_buf_1 place5941 (.A(_07044_),
    .X(net5940));
 sg13g2_buf_1 place5942 (.A(net5953),
    .X(net5941));
 sg13g2_buf_1 place5943 (.A(net5943),
    .X(net5942));
 sg13g2_buf_1 place5944 (.A(net5953),
    .X(net5943));
 sg13g2_buf_1 place5945 (.A(net5945),
    .X(net5944));
 sg13g2_buf_1 place5946 (.A(net5953),
    .X(net5945));
 sg13g2_buf_1 place5947 (.A(net5949),
    .X(net5946));
 sg13g2_buf_1 place5948 (.A(net5949),
    .X(net5947));
 sg13g2_buf_1 place5949 (.A(net5949),
    .X(net5948));
 sg13g2_buf_1 place5950 (.A(net5953),
    .X(net5949));
 sg13g2_buf_1 place5951 (.A(net5951),
    .X(net5950));
 sg13g2_buf_1 place5952 (.A(net5953),
    .X(net5951));
 sg13g2_buf_1 place5953 (.A(net5953),
    .X(net5952));
 sg13g2_buf_1 place5954 (.A(_07044_),
    .X(net5953));
 sg13g2_buf_1 place5955 (.A(_00090_),
    .X(net5954));
 sg13g2_buf_1 place5956 (.A(_00088_),
    .X(net5955));
 sg13g2_buf_1 place5958 (.A(net5961),
    .X(net5957));
 sg13g2_buf_1 place5959 (.A(net5961),
    .X(net5958));
 sg13g2_buf_1 place5960 (.A(net5961),
    .X(net5959));
 sg13g2_buf_1 place5961 (.A(net5961),
    .X(net5960));
 sg13g2_buf_8 place5962 (.A(_10893_),
    .X(net5961));
 sg13g2_buf_1 place5963 (.A(_10822_),
    .X(net5962));
 sg13g2_buf_1 place5964 (.A(_10822_),
    .X(net5963));
 sg13g2_buf_1 place5965 (.A(_10822_),
    .X(net5964));
 sg13g2_buf_1 place5966 (.A(_10822_),
    .X(net5965));
 sg13g2_buf_1 place5967 (.A(_10822_),
    .X(net5966));
 sg13g2_buf_2 place5968 (.A(_10691_),
    .X(net5967));
 sg13g2_buf_1 place5969 (.A(_07042_),
    .X(net5968));
 sg13g2_buf_2 place5970 (.A(_00087_),
    .X(net5969));
 sg13g2_buf_1 place5971 (.A(_00084_),
    .X(net5970));
 sg13g2_buf_1 place5972 (.A(_12816_),
    .X(net5971));
 sg13g2_buf_1 place5973 (.A(net5979),
    .X(net5972));
 sg13g2_buf_1 place5974 (.A(net5979),
    .X(net5973));
 sg13g2_buf_1 place5975 (.A(net5979),
    .X(net5974));
 sg13g2_buf_1 place5976 (.A(net5979),
    .X(net5975));
 sg13g2_buf_1 place5977 (.A(net5979),
    .X(net5976));
 sg13g2_buf_1 place5978 (.A(net5979),
    .X(net5977));
 sg13g2_buf_1 place5979 (.A(net5979),
    .X(net5978));
 sg13g2_buf_2 place5980 (.A(_12743_),
    .X(net5979));
 sg13g2_buf_1 place5981 (.A(_12743_),
    .X(net5980));
 sg13g2_buf_1 place5982 (.A(_12517_),
    .X(net5981));
 sg13g2_buf_1 place5983 (.A(_12441_),
    .X(net5982));
 sg13g2_buf_1 place5984 (.A(_12441_),
    .X(net5983));
 sg13g2_buf_1 place5985 (.A(net5991),
    .X(net5984));
 sg13g2_buf_2 place5986 (.A(net5991),
    .X(net5985));
 sg13g2_buf_1 place5987 (.A(net5991),
    .X(net5986));
 sg13g2_buf_1 place5988 (.A(net5991),
    .X(net5987));
 sg13g2_buf_1 place5989 (.A(net5991),
    .X(net5988));
 sg13g2_buf_1 place5990 (.A(net5991),
    .X(net5989));
 sg13g2_buf_1 place5991 (.A(net5991),
    .X(net5990));
 sg13g2_buf_4 place5992 (.X(net5991),
    .A(_12441_));
 sg13g2_buf_1 place5993 (.A(_12201_),
    .X(net5992));
 sg13g2_buf_1 place5994 (.A(_12119_),
    .X(net5993));
 sg13g2_buf_1 place5995 (.A(_11886_),
    .X(net5994));
 sg13g2_buf_1 place5996 (.A(_11804_),
    .X(net5995));
 sg13g2_buf_1 place5997 (.A(_11559_),
    .X(net5996));
 sg13g2_buf_1 place5998 (.A(_11481_),
    .X(net5997));
 sg13g2_buf_1 place5999 (.A(_11243_),
    .X(net5998));
 sg13g2_buf_1 place6000 (.A(_11161_),
    .X(net5999));
 sg13g2_buf_1 place6001 (.A(_10986_),
    .X(net6000));
 sg13g2_buf_1 place6002 (.A(net6007),
    .X(net6001));
 sg13g2_buf_1 place6003 (.A(net6007),
    .X(net6002));
 sg13g2_buf_1 place6004 (.A(net6007),
    .X(net6003));
 sg13g2_buf_1 place6005 (.A(net6007),
    .X(net6004));
 sg13g2_buf_1 place6006 (.A(net6007),
    .X(net6005));
 sg13g2_buf_1 place6007 (.A(net6007),
    .X(net6006));
 sg13g2_buf_2 place6008 (.A(_10962_),
    .X(net6007));
 sg13g2_buf_1 place6009 (.A(_10929_),
    .X(net6008));
 sg13g2_buf_1 place6010 (.A(_10929_),
    .X(net6009));
 sg13g2_buf_1 place6011 (.A(_10929_),
    .X(net6010));
 sg13g2_buf_1 place6012 (.A(_10929_),
    .X(net6011));
 sg13g2_buf_1 place6013 (.A(_10857_),
    .X(net6012));
 sg13g2_buf_1 place6014 (.A(_10857_),
    .X(net6013));
 sg13g2_buf_1 place6015 (.A(_10857_),
    .X(net6014));
 sg13g2_buf_1 place6016 (.A(_10857_),
    .X(net6015));
 sg13g2_buf_1 place6017 (.A(_10820_),
    .X(net6016));
 sg13g2_buf_1 place6018 (.A(_10127_),
    .X(net6017));
 sg13g2_buf_1 place6019 (.A(_10095_),
    .X(net6018));
 sg13g2_buf_1 place6020 (.A(_09961_),
    .X(net6019));
 sg13g2_buf_1 place6021 (.A(_09961_),
    .X(net6020));
 sg13g2_buf_1 place6022 (.A(_09961_),
    .X(net6021));
 sg13g2_buf_1 place6023 (.A(_09961_),
    .X(net6022));
 sg13g2_buf_2 place6024 (.A(net6028),
    .X(net6023));
 sg13g2_buf_1 place6025 (.A(net6028),
    .X(net6024));
 sg13g2_buf_2 place6026 (.A(net6028),
    .X(net6025));
 sg13g2_buf_1 place6027 (.A(net6028),
    .X(net6026));
 sg13g2_buf_1 place6028 (.A(net6028),
    .X(net6027));
 sg13g2_buf_8 place6029 (.A(_09902_),
    .X(net6028));
 sg13g2_buf_1 place6030 (.A(_09774_),
    .X(net6029));
 sg13g2_buf_1 place6031 (.A(_09774_),
    .X(net6030));
 sg13g2_buf_1 place6032 (.A(_09774_),
    .X(net6031));
 sg13g2_buf_2 place6033 (.A(_09774_),
    .X(net6032));
 sg13g2_buf_2 place6034 (.A(_09774_),
    .X(net6033));
 sg13g2_buf_1 place6035 (.A(net6035),
    .X(net6034));
 sg13g2_buf_1 place6036 (.A(net6036),
    .X(net6035));
 sg13g2_buf_2 place6037 (.A(_09686_),
    .X(net6036));
 sg13g2_buf_1 place6038 (.A(net6039),
    .X(net6037));
 sg13g2_buf_1 place6039 (.A(net6039),
    .X(net6038));
 sg13g2_buf_1 place6040 (.A(net6042),
    .X(net6039));
 sg13g2_buf_1 place6041 (.A(net6042),
    .X(net6040));
 sg13g2_buf_1 place6042 (.A(net6042),
    .X(net6041));
 sg13g2_buf_2 place6043 (.A(_09686_),
    .X(net6042));
 sg13g2_buf_1 place6044 (.A(_09611_),
    .X(net6043));
 sg13g2_buf_1 place6045 (.A(net6047),
    .X(net6044));
 sg13g2_buf_1 place6046 (.A(net6047),
    .X(net6045));
 sg13g2_buf_1 place6047 (.A(net6047),
    .X(net6046));
 sg13g2_buf_1 place6048 (.A(_09611_),
    .X(net6047));
 sg13g2_buf_1 place6049 (.A(net6050),
    .X(net6048));
 sg13g2_buf_1 place6050 (.A(net6050),
    .X(net6049));
 sg13g2_buf_2 place6051 (.A(_09611_),
    .X(net6050));
 sg13g2_buf_1 place6052 (.A(_09601_),
    .X(net6051));
 sg13g2_buf_1 place6053 (.A(net6053),
    .X(net6052));
 sg13g2_buf_1 place6054 (.A(_09601_),
    .X(net6053));
 sg13g2_buf_1 place6055 (.A(_09601_),
    .X(net6054));
 sg13g2_buf_1 place6056 (.A(_09601_),
    .X(net6055));
 sg13g2_buf_1 place6057 (.A(_06766_),
    .X(net6056));
 sg13g2_buf_1 place6058 (.A(_00083_),
    .X(net6057));
 sg13g2_buf_2 place6059 (.A(_00082_),
    .X(net6058));
 sg13g2_buf_1 place6060 (.A(_15205_),
    .X(net6059));
 sg13g2_buf_1 place6061 (.A(_15011_),
    .X(net6060));
 sg13g2_buf_1 place6062 (.A(net6063),
    .X(net6061));
 sg13g2_buf_1 place6063 (.A(net6063),
    .X(net6062));
 sg13g2_buf_1 place6064 (.A(_15011_),
    .X(net6063));
 sg13g2_buf_1 place6065 (.A(net6065),
    .X(net6064));
 sg13g2_buf_1 place6066 (.A(_15011_),
    .X(net6065));
 sg13g2_buf_1 place6067 (.A(net6067),
    .X(net6066));
 sg13g2_buf_1 place6068 (.A(_15011_),
    .X(net6067));
 sg13g2_buf_1 place6069 (.A(_12967_),
    .X(net6068));
 sg13g2_buf_1 place6070 (.A(_12891_),
    .X(net6069));
 sg13g2_buf_1 place6071 (.A(_12672_),
    .X(net6070));
 sg13g2_buf_1 place6072 (.A(_12597_),
    .X(net6071));
 sg13g2_buf_1 place6073 (.A(_12358_),
    .X(net6072));
 sg13g2_buf_1 place6074 (.A(net6074),
    .X(net6073));
 sg13g2_buf_1 place6075 (.A(_12282_),
    .X(net6074));
 sg13g2_buf_1 place6076 (.A(net6082),
    .X(net6075));
 sg13g2_buf_1 place6077 (.A(net6082),
    .X(net6076));
 sg13g2_buf_1 place6078 (.A(net6078),
    .X(net6077));
 sg13g2_buf_1 place6079 (.A(net6082),
    .X(net6078));
 sg13g2_buf_1 place6080 (.A(net6082),
    .X(net6079));
 sg13g2_buf_1 place6081 (.A(net6081),
    .X(net6080));
 sg13g2_buf_1 place6082 (.A(net6082),
    .X(net6081));
 sg13g2_buf_2 place6083 (.A(_12282_),
    .X(net6082));
 sg13g2_buf_1 place6084 (.A(_12042_),
    .X(net6083));
 sg13g2_buf_1 place6085 (.A(net6085),
    .X(net6084));
 sg13g2_buf_1 place6086 (.A(_12042_),
    .X(net6085));
 sg13g2_buf_1 place6087 (.A(_12042_),
    .X(net6086));
 sg13g2_buf_1 place6088 (.A(net6092),
    .X(net6087));
 sg13g2_buf_1 place6089 (.A(net6092),
    .X(net6088));
 sg13g2_buf_1 place6090 (.A(net6092),
    .X(net6089));
 sg13g2_buf_1 place6091 (.A(net6092),
    .X(net6090));
 sg13g2_buf_1 place6092 (.A(net6092),
    .X(net6091));
 sg13g2_buf_4 place6093 (.X(net6092),
    .A(_12042_));
 sg13g2_buf_1 place6094 (.A(_11966_),
    .X(net6093));
 sg13g2_buf_1 place6095 (.A(_11966_),
    .X(net6094));
 sg13g2_buf_1 place6096 (.A(_11800_),
    .X(net6095));
 sg13g2_buf_1 place6097 (.A(_11719_),
    .X(net6096));
 sg13g2_buf_2 place6098 (.A(_11639_),
    .X(net6097));
 sg13g2_buf_1 place6099 (.A(_11399_),
    .X(net6098));
 sg13g2_buf_1 place6100 (.A(_11322_),
    .X(net6099));
 sg13g2_buf_1 place6101 (.A(_11076_),
    .X(net6100));
 sg13g2_buf_2 place6102 (.A(_10992_),
    .X(net6101));
 sg13g2_buf_1 place6103 (.A(_10921_),
    .X(net6102));
 sg13g2_buf_1 place6104 (.A(_10852_),
    .X(net6103));
 sg13g2_buf_1 place6105 (.A(_10022_),
    .X(net6104));
 sg13g2_buf_1 place6106 (.A(_10022_),
    .X(net6105));
 sg13g2_buf_1 place6107 (.A(_10022_),
    .X(net6106));
 sg13g2_buf_1 place6108 (.A(_10022_),
    .X(net6107));
 sg13g2_buf_1 place6109 (.A(_10022_),
    .X(net6108));
 sg13g2_buf_1 place6110 (.A(net6114),
    .X(net6109));
 sg13g2_buf_1 place6111 (.A(net6114),
    .X(net6110));
 sg13g2_buf_1 place6112 (.A(net6114),
    .X(net6111));
 sg13g2_buf_1 place6113 (.A(net6114),
    .X(net6112));
 sg13g2_buf_1 place6114 (.A(net6114),
    .X(net6113));
 sg13g2_buf_1 place6115 (.A(_09841_),
    .X(net6114));
 sg13g2_buf_1 place6116 (.A(_09773_),
    .X(net6115));
 sg13g2_buf_1 place6117 (.A(_09685_),
    .X(net6116));
 sg13g2_buf_1 place6118 (.A(_09678_),
    .X(net6117));
 sg13g2_buf_1 place6119 (.A(_09678_),
    .X(net6118));
 sg13g2_buf_1 place6120 (.A(_09678_),
    .X(net6119));
 sg13g2_buf_1 place6121 (.A(_09678_),
    .X(net6120));
 sg13g2_buf_1 place6122 (.A(_09600_),
    .X(net6121));
 sg13g2_buf_1 place6126 (.A(net6126),
    .X(net6125));
 sg13g2_buf_1 place6127 (.A(_15021_),
    .X(net6126));
 sg13g2_buf_1 place6128 (.A(net6128),
    .X(net6127));
 sg13g2_buf_1 place6129 (.A(net6129),
    .X(net6128));
 sg13g2_buf_1 place6130 (.A(net6130),
    .X(net6129));
 sg13g2_buf_1 place6131 (.A(_15021_),
    .X(net6130));
 sg13g2_buf_1 place6132 (.A(_13703_),
    .X(net6131));
 sg13g2_buf_4 place6133 (.X(net6132),
    .A(_13610_));
 sg13g2_buf_1 place6134 (.A(net6134),
    .X(net6133));
 sg13g2_buf_1 place6135 (.A(_13553_),
    .X(net6134));
 sg13g2_buf_1 place6136 (.A(net6136),
    .X(net6135));
 sg13g2_buf_1 place6137 (.A(_13542_),
    .X(net6136));
 sg13g2_buf_1 place6138 (.A(_13527_),
    .X(net6137));
 sg13g2_buf_2 place6139 (.A(_13522_),
    .X(net6138));
 sg13g2_buf_1 place6140 (.A(net6140),
    .X(net6139));
 sg13g2_buf_1 place6141 (.A(_13516_),
    .X(net6140));
 sg13g2_buf_1 place6142 (.A(_13511_),
    .X(net6141));
 sg13g2_buf_1 place6143 (.A(_13506_),
    .X(net6142));
 sg13g2_buf_2 place6144 (.A(_13501_),
    .X(net6143));
 sg13g2_buf_2 place6145 (.A(_13495_),
    .X(net6144));
 sg13g2_buf_1 place6146 (.A(_13490_),
    .X(net6145));
 sg13g2_buf_1 place6147 (.A(_13490_),
    .X(net6146));
 sg13g2_buf_2 place6148 (.A(_13484_),
    .X(net6147));
 sg13g2_buf_1 place6149 (.A(_13484_),
    .X(net6148));
 sg13g2_buf_1 place6150 (.A(_13477_),
    .X(net6149));
 sg13g2_buf_2 place6151 (.A(_13471_),
    .X(net6150));
 sg13g2_buf_1 place6152 (.A(_13471_),
    .X(net6151));
 sg13g2_buf_1 place6153 (.A(_13465_),
    .X(net6152));
 sg13g2_buf_1 place6154 (.A(_13465_),
    .X(net6153));
 sg13g2_buf_1 place6155 (.A(net6155),
    .X(net6154));
 sg13g2_buf_1 place6156 (.A(_13451_),
    .X(net6155));
 sg13g2_buf_1 place6157 (.A(_13446_),
    .X(net6156));
 sg13g2_buf_1 place6158 (.A(_13446_),
    .X(net6157));
 sg13g2_buf_2 place6159 (.A(_13441_),
    .X(net6158));
 sg13g2_buf_2 place6160 (.A(_13436_),
    .X(net6159));
 sg13g2_buf_1 place6161 (.A(net6165),
    .X(net6160));
 sg13g2_buf_1 place6162 (.A(net6165),
    .X(net6161));
 sg13g2_buf_1 place6163 (.A(net6165),
    .X(net6162));
 sg13g2_buf_1 place6164 (.A(net6165),
    .X(net6163));
 sg13g2_buf_1 place6165 (.A(net6165),
    .X(net6164));
 sg13g2_buf_1 place6166 (.A(_12966_),
    .X(net6165));
 sg13g2_buf_1 place6167 (.A(net6168),
    .X(net6166));
 sg13g2_buf_1 place6168 (.A(net6168),
    .X(net6167));
 sg13g2_buf_1 place6169 (.A(_12966_),
    .X(net6168));
 sg13g2_buf_1 place6170 (.A(_12890_),
    .X(net6169));
 sg13g2_buf_1 place6171 (.A(net6171),
    .X(net6170));
 sg13g2_buf_1 place6172 (.A(_12890_),
    .X(net6171));
 sg13g2_buf_1 place6173 (.A(net6173),
    .X(net6172));
 sg13g2_buf_1 place6174 (.A(_12890_),
    .X(net6173));
 sg13g2_buf_1 place6175 (.A(net6175),
    .X(net6174));
 sg13g2_buf_1 place6176 (.A(_12890_),
    .X(net6175));
 sg13g2_buf_1 place6177 (.A(_12890_),
    .X(net6176));
 sg13g2_buf_1 place6178 (.A(_12815_),
    .X(net6177));
 sg13g2_buf_1 place6179 (.A(net6185),
    .X(net6178));
 sg13g2_buf_1 place6180 (.A(net6181),
    .X(net6179));
 sg13g2_buf_1 place6181 (.A(net6181),
    .X(net6180));
 sg13g2_buf_2 place6182 (.A(net6185),
    .X(net6181));
 sg13g2_buf_1 place6183 (.A(net6184),
    .X(net6182));
 sg13g2_buf_1 place6184 (.A(net6184),
    .X(net6183));
 sg13g2_buf_2 place6185 (.A(net6185),
    .X(net6184));
 sg13g2_buf_1 place6186 (.A(_12815_),
    .X(net6185));
 sg13g2_buf_1 place6187 (.A(_12671_),
    .X(net6186));
 sg13g2_buf_1 place6188 (.A(net6189),
    .X(net6187));
 sg13g2_buf_1 place6189 (.A(net6189),
    .X(net6188));
 sg13g2_buf_1 place6190 (.A(_12671_),
    .X(net6189));
 sg13g2_buf_1 place6191 (.A(net6193),
    .X(net6190));
 sg13g2_buf_1 place6192 (.A(net6193),
    .X(net6191));
 sg13g2_buf_1 place6193 (.A(net6193),
    .X(net6192));
 sg13g2_buf_1 place6194 (.A(_12671_),
    .X(net6193));
 sg13g2_buf_1 place6195 (.A(net6197),
    .X(net6194));
 sg13g2_buf_1 place6196 (.A(net6197),
    .X(net6195));
 sg13g2_buf_1 place6197 (.A(net6197),
    .X(net6196));
 sg13g2_buf_1 place6198 (.A(_12596_),
    .X(net6197));
 sg13g2_buf_1 place6199 (.A(net6200),
    .X(net6198));
 sg13g2_buf_1 place6200 (.A(net6200),
    .X(net6199));
 sg13g2_buf_1 place6201 (.A(_12596_),
    .X(net6200));
 sg13g2_buf_1 place6202 (.A(net6202),
    .X(net6201));
 sg13g2_buf_1 place6203 (.A(net6203),
    .X(net6202));
 sg13g2_buf_1 place6204 (.A(_12516_),
    .X(net6203));
 sg13g2_buf_1 place6205 (.A(net6206),
    .X(net6204));
 sg13g2_buf_1 place6206 (.A(net6206),
    .X(net6205));
 sg13g2_buf_2 place6207 (.A(net6208),
    .X(net6206));
 sg13g2_buf_1 place6208 (.A(net6208),
    .X(net6207));
 sg13g2_buf_1 place6209 (.A(_12516_),
    .X(net6208));
 sg13g2_buf_1 place6210 (.A(net6210),
    .X(net6209));
 sg13g2_buf_1 place6211 (.A(_12357_),
    .X(net6210));
 sg13g2_buf_1 place6212 (.A(net6215),
    .X(net6211));
 sg13g2_buf_1 place6213 (.A(net6215),
    .X(net6212));
 sg13g2_buf_1 place6214 (.A(net6215),
    .X(net6213));
 sg13g2_buf_1 place6215 (.A(net6215),
    .X(net6214));
 sg13g2_buf_1 place6216 (.A(_12357_),
    .X(net6215));
 sg13g2_buf_1 place6217 (.A(_12357_),
    .X(net6216));
 sg13g2_buf_1 place6218 (.A(net6218),
    .X(net6217));
 sg13g2_buf_2 place6219 (.A(_12200_),
    .X(net6218));
 sg13g2_buf_1 place6220 (.A(net6221),
    .X(net6219));
 sg13g2_buf_1 place6221 (.A(net6221),
    .X(net6220));
 sg13g2_buf_4 place6222 (.X(net6221),
    .A(_12200_));
 sg13g2_buf_1 place6223 (.A(net6224),
    .X(net6222));
 sg13g2_buf_2 place6224 (.A(net6224),
    .X(net6223));
 sg13g2_buf_1 place6225 (.A(_12200_),
    .X(net6224));
 sg13g2_buf_1 place6226 (.A(net6228),
    .X(net6225));
 sg13g2_buf_1 place6227 (.A(net6227),
    .X(net6226));
 sg13g2_buf_1 place6228 (.A(net6228),
    .X(net6227));
 sg13g2_buf_1 place6229 (.A(_12118_),
    .X(net6228));
 sg13g2_buf_1 place6230 (.A(net6231),
    .X(net6229));
 sg13g2_buf_1 place6231 (.A(net6231),
    .X(net6230));
 sg13g2_buf_1 place6232 (.A(net6232),
    .X(net6231));
 sg13g2_buf_1 place6233 (.A(_12118_),
    .X(net6232));
 sg13g2_buf_1 place6234 (.A(net6234),
    .X(net6233));
 sg13g2_buf_1 place6235 (.A(_11965_),
    .X(net6234));
 sg13g2_buf_1 place6236 (.A(_11965_),
    .X(net6235));
 sg13g2_buf_1 place6237 (.A(net6238),
    .X(net6236));
 sg13g2_buf_1 place6238 (.A(net6238),
    .X(net6237));
 sg13g2_buf_1 place6239 (.A(_11965_),
    .X(net6238));
 sg13g2_buf_1 place6240 (.A(net6240),
    .X(net6239));
 sg13g2_buf_1 place6241 (.A(_11965_),
    .X(net6240));
 sg13g2_buf_1 place6242 (.A(_11885_),
    .X(net6241));
 sg13g2_buf_1 place6243 (.A(net6244),
    .X(net6242));
 sg13g2_buf_1 place6244 (.A(net6244),
    .X(net6243));
 sg13g2_buf_1 place6245 (.A(_11885_),
    .X(net6244));
 sg13g2_buf_1 place6246 (.A(net6247),
    .X(net6245));
 sg13g2_buf_1 place6247 (.A(net6247),
    .X(net6246));
 sg13g2_buf_1 place6248 (.A(_11885_),
    .X(net6247));
 sg13g2_buf_1 place6249 (.A(net6249),
    .X(net6248));
 sg13g2_buf_1 place6250 (.A(_11885_),
    .X(net6249));
 sg13g2_buf_1 place6251 (.A(net6251),
    .X(net6250));
 sg13g2_buf_1 place6252 (.A(_11803_),
    .X(net6251));
 sg13g2_buf_1 place6253 (.A(net6253),
    .X(net6252));
 sg13g2_buf_1 place6254 (.A(net6254),
    .X(net6253));
 sg13g2_buf_1 place6255 (.A(net6258),
    .X(net6254));
 sg13g2_buf_1 place6256 (.A(net6256),
    .X(net6255));
 sg13g2_buf_1 place6257 (.A(net6258),
    .X(net6256));
 sg13g2_buf_1 place6258 (.A(net6258),
    .X(net6257));
 sg13g2_buf_1 place6259 (.A(_11803_),
    .X(net6258));
 sg13g2_buf_1 place6260 (.A(_11799_),
    .X(net6259));
 sg13g2_buf_1 place6261 (.A(net6261),
    .X(net6260));
 sg13g2_buf_1 place6262 (.A(net6262),
    .X(net6261));
 sg13g2_buf_1 place6263 (.A(_11798_),
    .X(net6262));
 sg13g2_buf_1 place6264 (.A(net6264),
    .X(net6263));
 sg13g2_buf_1 place6265 (.A(_11798_),
    .X(net6264));
 sg13g2_buf_1 place6266 (.A(net6267),
    .X(net6265));
 sg13g2_buf_1 place6267 (.A(net6267),
    .X(net6266));
 sg13g2_buf_1 place6268 (.A(_11798_),
    .X(net6267));
 sg13g2_buf_1 place6269 (.A(_11718_),
    .X(net6268));
 sg13g2_buf_1 place6270 (.A(net6270),
    .X(net6269));
 sg13g2_buf_1 place6271 (.A(_11718_),
    .X(net6270));
 sg13g2_buf_1 place6272 (.A(net6272),
    .X(net6271));
 sg13g2_buf_1 place6273 (.A(_11718_),
    .X(net6272));
 sg13g2_buf_1 place6274 (.A(net6274),
    .X(net6273));
 sg13g2_buf_1 place6275 (.A(_11718_),
    .X(net6274));
 sg13g2_buf_1 place6276 (.A(_11718_),
    .X(net6275));
 sg13g2_buf_1 place6277 (.A(_11718_),
    .X(net6276));
 sg13g2_buf_1 place6278 (.A(_11638_),
    .X(net6277));
 sg13g2_buf_2 place6279 (.A(net6285),
    .X(net6278));
 sg13g2_buf_1 place6280 (.A(net6285),
    .X(net6279));
 sg13g2_buf_1 place6281 (.A(net6285),
    .X(net6280));
 sg13g2_buf_1 place6282 (.A(net6285),
    .X(net6281));
 sg13g2_buf_1 place6283 (.A(net6285),
    .X(net6282));
 sg13g2_buf_2 place6284 (.A(net6284),
    .X(net6283));
 sg13g2_buf_4 place6285 (.X(net6284),
    .A(net6285));
 sg13g2_buf_8 place6286 (.A(_11638_),
    .X(net6285));
 sg13g2_buf_1 place6287 (.A(net6287),
    .X(net6286));
 sg13g2_buf_2 place6288 (.A(_11558_),
    .X(net6287));
 sg13g2_buf_1 place6289 (.A(net6290),
    .X(net6288));
 sg13g2_buf_1 place6290 (.A(net6290),
    .X(net6289));
 sg13g2_buf_1 place6291 (.A(_11558_),
    .X(net6290));
 sg13g2_buf_1 place6292 (.A(net6293),
    .X(net6291));
 sg13g2_buf_1 place6293 (.A(net6293),
    .X(net6292));
 sg13g2_buf_2 place6294 (.A(_11558_),
    .X(net6293));
 sg13g2_buf_1 place6295 (.A(_11558_),
    .X(net6294));
 sg13g2_buf_1 place6296 (.A(net6296),
    .X(net6295));
 sg13g2_buf_2 place6297 (.A(_11479_),
    .X(net6296));
 sg13g2_buf_1 place6298 (.A(net6299),
    .X(net6297));
 sg13g2_buf_1 place6299 (.A(net6299),
    .X(net6298));
 sg13g2_buf_1 place6300 (.A(_11479_),
    .X(net6299));
 sg13g2_buf_1 place6301 (.A(net6302),
    .X(net6300));
 sg13g2_buf_2 place6302 (.A(net6302),
    .X(net6301));
 sg13g2_buf_1 place6303 (.A(_11479_),
    .X(net6302));
 sg13g2_buf_1 place6304 (.A(_11479_),
    .X(net6303));
 sg13g2_buf_1 place6305 (.A(net6307),
    .X(net6304));
 sg13g2_buf_1 place6306 (.A(net6307),
    .X(net6305));
 sg13g2_buf_1 place6307 (.A(net6307),
    .X(net6306));
 sg13g2_buf_2 place6308 (.A(_11398_),
    .X(net6307));
 sg13g2_buf_1 place6309 (.A(_11398_),
    .X(net6308));
 sg13g2_buf_1 place6310 (.A(net6310),
    .X(net6309));
 sg13g2_buf_1 place6311 (.A(_11398_),
    .X(net6310));
 sg13g2_buf_1 place6312 (.A(net6315),
    .X(net6311));
 sg13g2_buf_1 place6313 (.A(net6315),
    .X(net6312));
 sg13g2_buf_1 place6314 (.A(net6315),
    .X(net6313));
 sg13g2_buf_1 place6315 (.A(net6315),
    .X(net6314));
 sg13g2_buf_1 place6316 (.A(_11321_),
    .X(net6315));
 sg13g2_buf_1 place6317 (.A(_11321_),
    .X(net6316));
 sg13g2_buf_1 place6318 (.A(net6318),
    .X(net6317));
 sg13g2_buf_1 place6319 (.A(_11321_),
    .X(net6318));
 sg13g2_buf_1 place6320 (.A(net6321),
    .X(net6319));
 sg13g2_buf_1 place6321 (.A(net6321),
    .X(net6320));
 sg13g2_buf_1 place6322 (.A(_11242_),
    .X(net6321));
 sg13g2_buf_1 place6323 (.A(_11242_),
    .X(net6322));
 sg13g2_buf_1 place6324 (.A(net6326),
    .X(net6323));
 sg13g2_buf_1 place6325 (.A(net6326),
    .X(net6324));
 sg13g2_buf_1 place6326 (.A(net6326),
    .X(net6325));
 sg13g2_buf_2 place6327 (.A(_11242_),
    .X(net6326));
 sg13g2_buf_1 place6328 (.A(_11160_),
    .X(net6327));
 sg13g2_buf_1 place6329 (.A(net6330),
    .X(net6328));
 sg13g2_buf_1 place6330 (.A(net6330),
    .X(net6329));
 sg13g2_buf_1 place6331 (.A(_11160_),
    .X(net6330));
 sg13g2_buf_1 place6332 (.A(net6334),
    .X(net6331));
 sg13g2_buf_1 place6333 (.A(net6334),
    .X(net6332));
 sg13g2_buf_1 place6334 (.A(net6334),
    .X(net6333));
 sg13g2_buf_1 place6335 (.A(_11160_),
    .X(net6334));
 sg13g2_buf_1 place6336 (.A(_11075_),
    .X(net6335));
 sg13g2_buf_1 place6337 (.A(_11075_),
    .X(net6336));
 sg13g2_buf_1 place6338 (.A(net6340),
    .X(net6337));
 sg13g2_buf_1 place6339 (.A(net6340),
    .X(net6338));
 sg13g2_buf_1 place6340 (.A(net6340),
    .X(net6339));
 sg13g2_buf_1 place6341 (.A(_11074_),
    .X(net6340));
 sg13g2_buf_1 place6342 (.A(_11074_),
    .X(net6341));
 sg13g2_buf_1 place6343 (.A(net6345),
    .X(net6342));
 sg13g2_buf_1 place6344 (.A(net6345),
    .X(net6343));
 sg13g2_buf_1 place6345 (.A(net6345),
    .X(net6344));
 sg13g2_buf_1 place6346 (.A(_11074_),
    .X(net6345));
 sg13g2_buf_1 place6347 (.A(_10991_),
    .X(net6346));
 sg13g2_buf_1 place6348 (.A(_10989_),
    .X(net6347));
 sg13g2_buf_1 place6349 (.A(net6351),
    .X(net6348));
 sg13g2_buf_1 place6350 (.A(net6351),
    .X(net6349));
 sg13g2_buf_1 place6351 (.A(net6351),
    .X(net6350));
 sg13g2_buf_1 place6352 (.A(_10989_),
    .X(net6351));
 sg13g2_buf_1 place6353 (.A(net6355),
    .X(net6352));
 sg13g2_buf_1 place6354 (.A(net6355),
    .X(net6353));
 sg13g2_buf_1 place6355 (.A(net6355),
    .X(net6354));
 sg13g2_buf_1 place6356 (.A(_10989_),
    .X(net6355));
 sg13g2_buf_1 place6357 (.A(net6357),
    .X(net6356));
 sg13g2_buf_1 place6358 (.A(_10984_),
    .X(net6357));
 sg13g2_buf_1 place6359 (.A(net6360),
    .X(net6358));
 sg13g2_buf_1 place6360 (.A(net6360),
    .X(net6359));
 sg13g2_buf_1 place6361 (.A(_10984_),
    .X(net6360));
 sg13g2_buf_1 place6362 (.A(net6362),
    .X(net6361));
 sg13g2_buf_1 place6363 (.A(_10984_),
    .X(net6362));
 sg13g2_buf_1 place6364 (.A(_10984_),
    .X(net6363));
 sg13g2_buf_1 place6365 (.A(net6365),
    .X(net6364));
 sg13g2_buf_1 place6366 (.A(_10493_),
    .X(net6365));
 sg13g2_buf_1 place6367 (.A(net6368),
    .X(net6366));
 sg13g2_buf_1 place6368 (.A(net6368),
    .X(net6367));
 sg13g2_buf_1 place6369 (.A(_10493_),
    .X(net6368));
 sg13g2_buf_1 place6370 (.A(net6376),
    .X(net6369));
 sg13g2_buf_1 place6371 (.A(net6376),
    .X(net6370));
 sg13g2_buf_1 place6372 (.A(net6376),
    .X(net6371));
 sg13g2_buf_1 place6373 (.A(net6376),
    .X(net6372));
 sg13g2_buf_1 place6374 (.A(net6376),
    .X(net6373));
 sg13g2_buf_1 place6375 (.A(net6376),
    .X(net6374));
 sg13g2_buf_1 place6376 (.A(net6376),
    .X(net6375));
 sg13g2_buf_1 place6377 (.A(_10415_),
    .X(net6376));
 sg13g2_buf_1 place6378 (.A(_10341_),
    .X(net6377));
 sg13g2_buf_1 place6379 (.A(_10341_),
    .X(net6378));
 sg13g2_buf_1 place6380 (.A(_10341_),
    .X(net6379));
 sg13g2_buf_1 place6381 (.A(_10341_),
    .X(net6380));
 sg13g2_buf_1 place6382 (.A(net6382),
    .X(net6381));
 sg13g2_buf_1 place6383 (.A(_10162_),
    .X(net6382));
 sg13g2_buf_1 place6384 (.A(net6384),
    .X(net6383));
 sg13g2_buf_1 place6385 (.A(_10162_),
    .X(net6384));
 sg13g2_buf_1 place6386 (.A(_10104_),
    .X(net6385));
 sg13g2_buf_1 place6387 (.A(_10093_),
    .X(net6386));
 sg13g2_buf_1 place6388 (.A(net6393),
    .X(net6387));
 sg13g2_buf_1 place6389 (.A(net6393),
    .X(net6388));
 sg13g2_buf_2 place6390 (.A(net6393),
    .X(net6389));
 sg13g2_buf_1 place6391 (.A(net6392),
    .X(net6390));
 sg13g2_buf_1 place6392 (.A(net6392),
    .X(net6391));
 sg13g2_buf_4 place6393 (.X(net6392),
    .A(net6393));
 sg13g2_buf_4 place6394 (.X(net6393),
    .A(_10093_));
 sg13g2_buf_1 place6395 (.A(_10009_),
    .X(net6394));
 sg13g2_buf_1 place6396 (.A(_06741_),
    .X(net6395));
 sg13g2_buf_1 place6398 (.A(_00081_),
    .X(net6397));
 sg13g2_buf_1 place6399 (.A(_00080_),
    .X(net6398));
 sg13g2_buf_1 place6400 (.A(_00079_),
    .X(net6399));
 sg13g2_buf_1 place6401 (.A(_00111_),
    .X(net6400));
 sg13g2_buf_1 place6406 (.A(net6409),
    .X(net6405));
 sg13g2_buf_1 place6407 (.A(net6407),
    .X(net6406));
 sg13g2_buf_1 place6408 (.A(net6408),
    .X(net6407));
 sg13g2_buf_1 place6409 (.A(net6409),
    .X(net6408));
 sg13g2_buf_1 place6410 (.A(_15048_),
    .X(net6409));
 sg13g2_buf_1 place6411 (.A(net6414),
    .X(net6410));
 sg13g2_buf_1 place6412 (.A(net6412),
    .X(net6411));
 sg13g2_buf_1 place6413 (.A(net6413),
    .X(net6412));
 sg13g2_buf_1 place6414 (.A(net6414),
    .X(net6413));
 sg13g2_buf_1 place6415 (.A(_15048_),
    .X(net6414));
 sg13g2_buf_1 place6416 (.A(net6416),
    .X(net6415));
 sg13g2_buf_1 place6417 (.A(_15022_),
    .X(net6416));
 sg13g2_buf_1 place6418 (.A(_15022_),
    .X(net6417));
 sg13g2_buf_1 place6419 (.A(net6419),
    .X(net6418));
 sg13g2_buf_1 place6420 (.A(_15020_),
    .X(net6419));
 sg13g2_buf_1 place6421 (.A(_15020_),
    .X(net6420));
 sg13g2_buf_1 place6422 (.A(net6422),
    .X(net6421));
 sg13g2_buf_1 place6423 (.A(net6423),
    .X(net6422));
 sg13g2_buf_1 place6424 (.A(_15020_),
    .X(net6423));
 sg13g2_buf_1 place6425 (.A(net6425),
    .X(net6424));
 sg13g2_buf_1 place6426 (.A(net6426),
    .X(net6425));
 sg13g2_buf_1 place6427 (.A(_15020_),
    .X(net6426));
 sg13g2_buf_1 place6428 (.A(net6428),
    .X(net6427));
 sg13g2_buf_1 place6429 (.A(net6430),
    .X(net6428));
 sg13g2_buf_1 place6430 (.A(net6430),
    .X(net6429));
 sg13g2_buf_2 place6431 (.A(_15020_),
    .X(net6430));
 sg13g2_buf_1 place6432 (.A(net6433),
    .X(net6431));
 sg13g2_buf_1 place6433 (.A(net6433),
    .X(net6432));
 sg13g2_buf_1 place6434 (.A(net6434),
    .X(net6433));
 sg13g2_buf_1 place6435 (.A(_14582_),
    .X(net6434));
 sg13g2_buf_1 place6436 (.A(_14571_),
    .X(net6435));
 sg13g2_buf_1 place6437 (.A(_14571_),
    .X(net6436));
 sg13g2_buf_1 place6438 (.A(net6440),
    .X(net6437));
 sg13g2_buf_1 place6439 (.A(net6439),
    .X(net6438));
 sg13g2_buf_1 place6440 (.A(net6440),
    .X(net6439));
 sg13g2_buf_1 place6441 (.A(_14571_),
    .X(net6440));
 sg13g2_buf_1 place6442 (.A(net6453),
    .X(net6441));
 sg13g2_buf_1 place6443 (.A(net6444),
    .X(net6442));
 sg13g2_buf_1 place6444 (.A(net6444),
    .X(net6443));
 sg13g2_buf_1 place6445 (.A(net6453),
    .X(net6444));
 sg13g2_buf_1 place6446 (.A(net6446),
    .X(net6445));
 sg13g2_buf_1 place6447 (.A(net6453),
    .X(net6446));
 sg13g2_buf_1 place6448 (.A(net6453),
    .X(net6447));
 sg13g2_buf_1 place6449 (.A(net6452),
    .X(net6448));
 sg13g2_buf_1 place6450 (.A(net6452),
    .X(net6449));
 sg13g2_buf_1 place6451 (.A(net6452),
    .X(net6450));
 sg13g2_buf_1 place6452 (.A(net6452),
    .X(net6451));
 sg13g2_buf_1 place6453 (.A(net6453),
    .X(net6452));
 sg13g2_buf_1 place6454 (.A(_14570_),
    .X(net6453));
 sg13g2_buf_1 place6455 (.A(_13779_),
    .X(net6454));
 sg13g2_buf_2 place6456 (.A(_13559_),
    .X(net6455));
 sg13g2_buf_1 place6457 (.A(_13547_),
    .X(net6456));
 sg13g2_buf_1 place6458 (.A(_13547_),
    .X(net6457));
 sg13g2_buf_1 place6459 (.A(_13458_),
    .X(net6458));
 sg13g2_buf_1 place6460 (.A(_13431_),
    .X(net6459));
 sg13g2_buf_1 place6461 (.A(net6461),
    .X(net6460));
 sg13g2_buf_1 place6462 (.A(_13427_),
    .X(net6461));
 sg13g2_buf_1 place6463 (.A(_13427_),
    .X(net6462));
 sg13g2_buf_1 place6464 (.A(net6464),
    .X(net6463));
 sg13g2_buf_1 place6465 (.A(_10101_),
    .X(net6464));
 sg13g2_buf_1 place6466 (.A(_10101_),
    .X(net6465));
 sg13g2_buf_1 place6467 (.A(_09604_),
    .X(net6466));
 sg13g2_buf_1 place6468 (.A(net6468),
    .X(net6467));
 sg13g2_buf_1 place6469 (.A(_09603_),
    .X(net6468));
 sg13g2_buf_1 place6470 (.A(net6472),
    .X(net6469));
 sg13g2_buf_1 place6471 (.A(net6471),
    .X(net6470));
 sg13g2_buf_1 place6472 (.A(net6472),
    .X(net6471));
 sg13g2_buf_1 place6473 (.A(_08728_),
    .X(net6472));
 sg13g2_buf_1 place6474 (.A(net6474),
    .X(net6473));
 sg13g2_buf_1 place6475 (.A(_08728_),
    .X(net6474));
 sg13g2_buf_1 place6479 (.A(_00110_),
    .X(net6478));
 sg13g2_buf_1 place6480 (.A(_00108_),
    .X(net6479));
 sg13g2_buf_1 place6488 (.A(_14531_),
    .X(net6487));
 sg13g2_buf_1 place6489 (.A(net6490),
    .X(net6488));
 sg13g2_buf_1 place6490 (.A(net6490),
    .X(net6489));
 sg13g2_buf_1 place6491 (.A(net6491),
    .X(net6490));
 sg13g2_buf_1 place6492 (.A(_14426_),
    .X(net6491));
 sg13g2_buf_1 place6493 (.A(_14426_),
    .X(net6492));
 sg13g2_buf_1 place6494 (.A(net6494),
    .X(net6493));
 sg13g2_buf_1 place6495 (.A(_14353_),
    .X(net6494));
 sg13g2_buf_1 place6496 (.A(net6500),
    .X(net6495));
 sg13g2_buf_1 place6497 (.A(net6497),
    .X(net6496));
 sg13g2_buf_1 place6498 (.A(net6500),
    .X(net6497));
 sg13g2_buf_1 place6499 (.A(net6499),
    .X(net6498));
 sg13g2_buf_1 place6500 (.A(net6500),
    .X(net6499));
 sg13g2_buf_1 place6501 (.A(_14353_),
    .X(net6500));
 sg13g2_buf_1 place6502 (.A(_14353_),
    .X(net6501));
 sg13g2_buf_1 place6503 (.A(net6504),
    .X(net6502));
 sg13g2_buf_1 place6504 (.A(net6504),
    .X(net6503));
 sg13g2_buf_1 place6505 (.A(_14282_),
    .X(net6504));
 sg13g2_buf_1 place6506 (.A(net6506),
    .X(net6505));
 sg13g2_buf_1 place6507 (.A(net6507),
    .X(net6506));
 sg13g2_buf_1 place6508 (.A(net6511),
    .X(net6507));
 sg13g2_buf_1 place6509 (.A(net6509),
    .X(net6508));
 sg13g2_buf_1 place6510 (.A(net6511),
    .X(net6509));
 sg13g2_buf_1 place6511 (.A(net6511),
    .X(net6510));
 sg13g2_buf_1 place6512 (.A(_14282_),
    .X(net6511));
 sg13g2_buf_1 place6513 (.A(_14246_),
    .X(net6512));
 sg13g2_buf_1 place6514 (.A(_14075_),
    .X(net6513));
 sg13g2_buf_1 place6515 (.A(net6515),
    .X(net6514));
 sg13g2_buf_1 place6516 (.A(_14075_),
    .X(net6515));
 sg13g2_buf_1 place6517 (.A(net6517),
    .X(net6516));
 sg13g2_buf_1 place6518 (.A(_14075_),
    .X(net6517));
 sg13g2_buf_1 place6519 (.A(_14033_),
    .X(net6518));
 sg13g2_buf_1 place6520 (.A(net6522),
    .X(net6519));
 sg13g2_buf_1 place6521 (.A(net6521),
    .X(net6520));
 sg13g2_buf_1 place6522 (.A(net6522),
    .X(net6521));
 sg13g2_buf_1 place6523 (.A(_14033_),
    .X(net6522));
 sg13g2_buf_1 place6524 (.A(net6524),
    .X(net6523));
 sg13g2_buf_1 place6525 (.A(_13959_),
    .X(net6524));
 sg13g2_buf_1 place6526 (.A(net6526),
    .X(net6525));
 sg13g2_buf_1 place6527 (.A(_13959_),
    .X(net6526));
 sg13g2_buf_1 place6528 (.A(net6531),
    .X(net6527));
 sg13g2_buf_1 place6529 (.A(net6529),
    .X(net6528));
 sg13g2_buf_1 place6530 (.A(net6531),
    .X(net6529));
 sg13g2_buf_1 place6531 (.A(net6531),
    .X(net6530));
 sg13g2_buf_1 place6532 (.A(_13959_),
    .X(net6531));
 sg13g2_buf_1 place6533 (.A(_13880_),
    .X(net6532));
 sg13g2_buf_1 place6534 (.A(_13634_),
    .X(net6533));
 sg13g2_buf_1 place6535 (.A(net6535),
    .X(net6534));
 sg13g2_buf_1 place6536 (.A(_13576_),
    .X(net6535));
 sg13g2_buf_1 place6537 (.A(_13576_),
    .X(net6536));
 sg13g2_buf_1 place6538 (.A(net6538),
    .X(net6537));
 sg13g2_buf_1 place6539 (.A(_13574_),
    .X(net6538));
 sg13g2_buf_1 place6540 (.A(net6540),
    .X(net6539));
 sg13g2_buf_1 place6541 (.A(_13574_),
    .X(net6540));
 sg13g2_buf_1 place6542 (.A(_13574_),
    .X(net6541));
 sg13g2_buf_1 place6543 (.A(_13537_),
    .X(net6542));
 sg13g2_buf_1 place6544 (.A(_13532_),
    .X(net6543));
 sg13g2_buf_1 place6545 (.A(_13424_),
    .X(net6544));
 sg13g2_buf_1 place6546 (.A(net6546),
    .X(net6545));
 sg13g2_buf_1 place6547 (.A(_13424_),
    .X(net6546));
 sg13g2_buf_1 place6548 (.A(_09365_),
    .X(net6547));
 sg13g2_buf_1 place6549 (.A(net6550),
    .X(net6548));
 sg13g2_buf_1 place6550 (.A(net6550),
    .X(net6549));
 sg13g2_buf_1 place6551 (.A(net6551),
    .X(net6550));
 sg13g2_buf_1 place6552 (.A(_09364_),
    .X(net6551));
 sg13g2_buf_2 place6553 (.A(_09364_),
    .X(net6552));
 sg13g2_buf_1 place6554 (.A(_08033_),
    .X(net6553));
 sg13g2_buf_1 place6555 (.A(_08022_),
    .X(net6554));
 sg13g2_buf_1 place6558 (.A(_00109_),
    .X(net6557));
 sg13g2_buf_2 place6568 (.A(net462),
    .X(net6567));
 sg13g2_buf_1 place6569 (.A(net462),
    .X(net6568));
 sg13g2_buf_1 place6570 (.A(net461),
    .X(net6569));
 sg13g2_buf_2 place6571 (.A(net461),
    .X(net6570));
 sg13g2_buf_8 place6572 (.A(net459),
    .X(net6571));
 sg13g2_buf_1 place6573 (.A(net458),
    .X(net6572));
 sg13g2_buf_2 place6574 (.A(net458),
    .X(net6573));
 sg13g2_buf_1 place6575 (.A(net457),
    .X(net6574));
 sg13g2_buf_4 place6576 (.X(net6575),
    .A(net457));
 sg13g2_buf_1 place6577 (.A(net6577),
    .X(net6576));
 sg13g2_buf_2 place6578 (.A(net456),
    .X(net6577));
 sg13g2_buf_1 place6579 (.A(net455),
    .X(net6578));
 sg13g2_buf_1 place6580 (.A(net6580),
    .X(net6579));
 sg13g2_buf_1 place6581 (.A(net455),
    .X(net6580));
 sg13g2_buf_1 place6582 (.A(net454),
    .X(net6581));
 sg13g2_buf_1 place6583 (.A(net6583),
    .X(net6582));
 sg13g2_buf_1 place6584 (.A(net454),
    .X(net6583));
 sg13g2_buf_4 place6585 (.X(net6584),
    .A(net451));
 sg13g2_buf_1 place6586 (.A(net450),
    .X(net6585));
 sg13g2_buf_1 place6587 (.A(net450),
    .X(net6586));
 sg13g2_buf_1 place6588 (.A(net6589),
    .X(net6587));
 sg13g2_buf_1 place6589 (.A(net6589),
    .X(net6588));
 sg13g2_buf_1 place6590 (.A(net6591),
    .X(net6589));
 sg13g2_buf_1 place6591 (.A(net6591),
    .X(net6590));
 sg13g2_buf_1 place6592 (.A(_14425_),
    .X(net6591));
 sg13g2_buf_1 place6593 (.A(_13420_),
    .X(net6592));
 sg13g2_buf_1 place6600 (.A(net443),
    .X(net6599));
 sg13g2_buf_1 place6601 (.A(net443),
    .X(net6600));
 sg13g2_buf_1 place6602 (.A(net442),
    .X(net6601));
 sg13g2_buf_1 place6603 (.A(net442),
    .X(net6602));
 sg13g2_buf_1 place6604 (.A(net6604),
    .X(net6603));
 sg13g2_buf_2 place6605 (.A(net453),
    .X(net6604));
 sg13g2_buf_1 place6606 (.A(net6606),
    .X(net6605));
 sg13g2_buf_2 place6607 (.A(net452),
    .X(net6606));
 sg13g2_buf_4 place6608 (.X(net6607),
    .A(net449));
 sg13g2_buf_4 place6609 (.X(net6608),
    .A(net448));
 sg13g2_buf_4 place6610 (.X(net6609),
    .A(net447));
 sg13g2_buf_1 place6611 (.A(net446),
    .X(net6610));
 sg13g2_buf_1 place6612 (.A(net446),
    .X(net6611));
 sg13g2_buf_1 place6613 (.A(net445),
    .X(net6612));
 sg13g2_buf_1 place6614 (.A(net445),
    .X(net6613));
 sg13g2_buf_1 place6615 (.A(net444),
    .X(net6614));
 sg13g2_buf_1 place6616 (.A(net444),
    .X(net6615));
 sg13g2_buf_1 place6618 (.A(_06381_),
    .X(net6617));
 sg13g2_buf_1 place6621 (.A(_00106_),
    .X(net6620));
 sg13g2_buf_4 place6622 (.X(net6621),
    .A(net441));
 sg13g2_buf_1 place6623 (.A(net440),
    .X(net6622));
 sg13g2_buf_1 place6624 (.A(net440),
    .X(net6623));
 sg13g2_buf_1 place6625 (.A(net469),
    .X(net6624));
 sg13g2_buf_1 place6626 (.A(net469),
    .X(net6625));
 sg13g2_buf_1 place6627 (.A(net468),
    .X(net6626));
 sg13g2_buf_1 place6628 (.A(net467),
    .X(net6627));
 sg13g2_buf_1 place6629 (.A(net466),
    .X(net6628));
 sg13g2_buf_1 place6630 (.A(net6630),
    .X(net6629));
 sg13g2_buf_1 place6631 (.A(_14076_),
    .X(net6630));
 sg13g2_buf_1 place6632 (.A(net6632),
    .X(net6631));
 sg13g2_buf_1 place6633 (.A(_14076_),
    .X(net6632));
 sg13g2_buf_1 place6636 (.A(_00105_),
    .X(net6635));
 sg13g2_buf_1 place6637 (.A(net465),
    .X(net6636));
 sg13g2_buf_1 place6638 (.A(net465),
    .X(net6637));
 sg13g2_buf_1 place6639 (.A(net464),
    .X(net6638));
 sg13g2_buf_1 place6640 (.A(net463),
    .X(net6639));
 sg13g2_buf_1 place6641 (.A(net460),
    .X(net6640));
 sg13g2_buf_1 place6642 (.A(net6644),
    .X(net6641));
 sg13g2_buf_1 place6643 (.A(net6643),
    .X(net6642));
 sg13g2_buf_1 place6644 (.A(net6644),
    .X(net6643));
 sg13g2_buf_1 place6645 (.A(_13578_),
    .X(net6644));
 sg13g2_buf_1 place6646 (.A(_07712_),
    .X(net6645));
 sg13g2_buf_1 place6647 (.A(net6648),
    .X(net6646));
 sg13g2_buf_1 place6648 (.A(net6648),
    .X(net6647));
 sg13g2_buf_1 place6649 (.A(_07712_),
    .X(net6648));
 sg13g2_buf_1 place6650 (.A(net6650),
    .X(net6649));
 sg13g2_buf_1 place6651 (.A(_06865_),
    .X(net6650));
 sg13g2_buf_1 place6652 (.A(net6652),
    .X(net6651));
 sg13g2_buf_1 place6653 (.A(_06865_),
    .X(net6652));
 sg13g2_buf_1 place6654 (.A(net6656),
    .X(net6653));
 sg13g2_buf_1 place6655 (.A(net6655),
    .X(net6654));
 sg13g2_buf_1 place6656 (.A(net6656),
    .X(net6655));
 sg13g2_buf_1 place6657 (.A(net6657),
    .X(net6656));
 sg13g2_buf_1 place6658 (.A(_13573_),
    .X(net6657));
 sg13g2_buf_1 place6659 (.A(net6667),
    .X(net6658));
 sg13g2_buf_1 place6660 (.A(net6661),
    .X(net6659));
 sg13g2_buf_1 place6661 (.A(net6661),
    .X(net6660));
 sg13g2_buf_1 place6662 (.A(net6667),
    .X(net6661));
 sg13g2_buf_1 place6663 (.A(net6667),
    .X(net6662));
 sg13g2_buf_1 place6664 (.A(net6667),
    .X(net6663));
 sg13g2_buf_1 place6665 (.A(net6667),
    .X(net6664));
 sg13g2_buf_1 place6666 (.A(net6666),
    .X(net6665));
 sg13g2_buf_1 place6667 (.A(net6667),
    .X(net6666));
 sg13g2_buf_1 place6668 (.A(net6668),
    .X(net6667));
 sg13g2_buf_1 place6669 (.A(_13572_),
    .X(net6668));
 sg13g2_buf_1 place6670 (.A(_13572_),
    .X(net6669));
 sg13g2_buf_1 place6671 (.A(net6672),
    .X(net6670));
 sg13g2_buf_1 place6672 (.A(net6672),
    .X(net6671));
 sg13g2_buf_1 place6673 (.A(_10065_),
    .X(net6672));
 sg13g2_buf_1 place6674 (.A(_09661_),
    .X(net6673));
 sg13g2_buf_1 place6675 (.A(net6676),
    .X(net6674));
 sg13g2_buf_1 place6676 (.A(net6676),
    .X(net6675));
 sg13g2_buf_1 place6677 (.A(_09572_),
    .X(net6676));
 sg13g2_buf_1 place6678 (.A(_09572_),
    .X(net6677));
 sg13g2_buf_1 place6679 (.A(net6679),
    .X(net6678));
 sg13g2_buf_1 place6680 (.A(_09570_),
    .X(net6679));
 sg13g2_buf_1 place6681 (.A(_09570_),
    .X(net6680));
 sg13g2_buf_1 place6682 (.A(_09570_),
    .X(net6681));
 sg13g2_buf_1 place6683 (.A(net6684),
    .X(net6682));
 sg13g2_buf_1 place6684 (.A(net6684),
    .X(net6683));
 sg13g2_buf_1 place6685 (.A(_09569_),
    .X(net6684));
 sg13g2_buf_1 place6686 (.A(_09569_),
    .X(net6685));
 sg13g2_buf_1 place6687 (.A(net6687),
    .X(net6686));
 sg13g2_buf_1 place6688 (.A(net6688),
    .X(net6687));
 sg13g2_buf_1 place6689 (.A(_09568_),
    .X(net6688));
 sg13g2_buf_1 place6690 (.A(_09568_),
    .X(net6689));
 sg13g2_buf_1 place6691 (.A(net6691),
    .X(net6690));
 sg13g2_buf_1 place6692 (.A(_09567_),
    .X(net6691));
 sg13g2_buf_1 place6693 (.A(net6694),
    .X(net6692));
 sg13g2_buf_1 place6694 (.A(net6694),
    .X(net6693));
 sg13g2_buf_1 place6695 (.A(_09567_),
    .X(net6694));
 sg13g2_buf_1 place6696 (.A(_09566_),
    .X(net6695));
 sg13g2_buf_1 place6697 (.A(net6698),
    .X(net6696));
 sg13g2_buf_2 place6698 (.A(net6698),
    .X(net6697));
 sg13g2_buf_1 place6699 (.A(_09566_),
    .X(net6698));
 sg13g2_buf_1 place6700 (.A(net6700),
    .X(net6699));
 sg13g2_buf_1 place6701 (.A(net6701),
    .X(net6700));
 sg13g2_buf_1 place6702 (.A(_09563_),
    .X(net6701));
 sg13g2_buf_1 place6703 (.A(_09563_),
    .X(net6702));
 sg13g2_buf_1 place6704 (.A(_09560_),
    .X(net6703));
 sg13g2_buf_1 place6705 (.A(_09560_),
    .X(net6704));
 sg13g2_buf_1 place6706 (.A(net6706),
    .X(net6705));
 sg13g2_buf_1 place6707 (.A(_09558_),
    .X(net6706));
 sg13g2_buf_1 place6708 (.A(_06940_),
    .X(net6707));
 sg13g2_buf_1 place6709 (.A(net6709),
    .X(net6708));
 sg13g2_buf_1 place6710 (.A(net6711),
    .X(net6709));
 sg13g2_buf_1 place6711 (.A(net6711),
    .X(net6710));
 sg13g2_buf_1 place6712 (.A(_06919_),
    .X(net6711));
 sg13g2_buf_1 place6713 (.A(net6713),
    .X(net6712));
 sg13g2_buf_1 place6714 (.A(_06850_),
    .X(net6713));
 sg13g2_buf_1 place6715 (.A(_06134_),
    .X(net6714));
 sg13g2_buf_1 place6716 (.A(_05513_),
    .X(net6715));
 sg13g2_buf_1 place6717 (.A(_05264_),
    .X(net6716));
 sg13g2_buf_1 place6718 (.A(\alu_adder_result_ex[1] ),
    .X(net6717));
 sg13g2_buf_1 place6719 (.A(net6720),
    .X(net6718));
 sg13g2_buf_1 place6720 (.A(net6720),
    .X(net6719));
 sg13g2_buf_1 place6721 (.A(net6725),
    .X(net6720));
 sg13g2_buf_1 place6722 (.A(net6725),
    .X(net6721));
 sg13g2_buf_1 place6723 (.A(net6725),
    .X(net6722));
 sg13g2_buf_1 place6724 (.A(net6724),
    .X(net6723));
 sg13g2_buf_4 place6725 (.X(net6724),
    .A(net6725));
 sg13g2_buf_2 place6726 (.A(\alu_adder_result_ex[1] ),
    .X(net6725));
 sg13g2_buf_1 place6727 (.A(net6727),
    .X(net6726));
 sg13g2_buf_1 place6728 (.A(\alu_adder_result_ex[1] ),
    .X(net6727));
 sg13g2_buf_1 place6729 (.A(_13565_),
    .X(net6728));
 sg13g2_buf_1 place6730 (.A(_13418_),
    .X(net6729));
 sg13g2_buf_1 place6731 (.A(net6731),
    .X(net6730));
 sg13g2_buf_1 place6732 (.A(_13418_),
    .X(net6731));
 sg13g2_buf_1 place6733 (.A(net6733),
    .X(net6732));
 sg13g2_buf_1 place6734 (.A(_07026_),
    .X(net6733));
 sg13g2_buf_1 place6735 (.A(net6735),
    .X(net6734));
 sg13g2_buf_1 place6736 (.A(_07026_),
    .X(net6735));
 sg13g2_buf_1 place6737 (.A(_06696_),
    .X(net6736));
 sg13g2_buf_1 place6738 (.A(_06696_),
    .X(net6737));
 sg13g2_buf_1 place6739 (.A(net6739),
    .X(net6738));
 sg13g2_buf_1 place6740 (.A(_06696_),
    .X(net6739));
 sg13g2_buf_1 place6741 (.A(_05591_),
    .X(net6740));
 sg13g2_buf_1 place6742 (.A(_04817_),
    .X(net6741));
 sg13g2_buf_1 place6743 (.A(net6743),
    .X(net6742));
 sg13g2_buf_1 place6744 (.A(\alu_adder_result_ex[0] ),
    .X(net6743));
 sg13g2_buf_1 place6745 (.A(net6745),
    .X(net6744));
 sg13g2_buf_1 place6746 (.A(net6747),
    .X(net6745));
 sg13g2_buf_1 place6747 (.A(net6747),
    .X(net6746));
 sg13g2_buf_1 place6748 (.A(\alu_adder_result_ex[0] ),
    .X(net6747));
 sg13g2_buf_1 place6749 (.A(_15078_),
    .X(net6748));
 sg13g2_buf_1 place6750 (.A(net6752),
    .X(net6749));
 sg13g2_buf_1 place6751 (.A(net6751),
    .X(net6750));
 sg13g2_buf_1 place6752 (.A(net6752),
    .X(net6751));
 sg13g2_buf_1 place6753 (.A(_13162_),
    .X(net6752));
 sg13g2_buf_1 place6754 (.A(net6754),
    .X(net6753));
 sg13g2_buf_1 place6755 (.A(net6755),
    .X(net6754));
 sg13g2_buf_1 place6756 (.A(_09406_),
    .X(net6755));
 sg13g2_buf_1 place6757 (.A(_09405_),
    .X(net6756));
 sg13g2_buf_1 place6758 (.A(net6758),
    .X(net6757));
 sg13g2_buf_1 place6759 (.A(_09405_),
    .X(net6758));
 sg13g2_buf_1 place6760 (.A(_08969_),
    .X(net6759));
 sg13g2_buf_1 place6761 (.A(net6762),
    .X(net6760));
 sg13g2_buf_1 place6762 (.A(net6762),
    .X(net6761));
 sg13g2_buf_1 place6763 (.A(_07093_),
    .X(net6762));
 sg13g2_buf_1 place6764 (.A(net6767),
    .X(net6763));
 sg13g2_buf_1 place6765 (.A(net6766),
    .X(net6764));
 sg13g2_buf_1 place6766 (.A(net6766),
    .X(net6765));
 sg13g2_buf_1 place6767 (.A(net6767),
    .X(net6766));
 sg13g2_buf_1 place6768 (.A(_07093_),
    .X(net6767));
 sg13g2_buf_1 place6769 (.A(_07093_),
    .X(net6768));
 sg13g2_buf_1 place6770 (.A(net6770),
    .X(net6769));
 sg13g2_buf_1 place6771 (.A(_07092_),
    .X(net6770));
 sg13g2_buf_1 place6772 (.A(net6773),
    .X(net6771));
 sg13g2_buf_1 place6773 (.A(net6773),
    .X(net6772));
 sg13g2_buf_1 place6774 (.A(_07092_),
    .X(net6773));
 sg13g2_buf_1 place6775 (.A(net6775),
    .X(net6774));
 sg13g2_buf_1 place6776 (.A(net6776),
    .X(net6775));
 sg13g2_buf_2 place6777 (.A(_07092_),
    .X(net6776));
 sg13g2_buf_1 place6778 (.A(net6778),
    .X(net6777));
 sg13g2_buf_2 place6779 (.A(net6780),
    .X(net6778));
 sg13g2_buf_1 place6780 (.A(net6780),
    .X(net6779));
 sg13g2_buf_1 place6781 (.A(_06886_),
    .X(net6780));
 sg13g2_buf_1 place6782 (.A(_06886_),
    .X(net6781));
 sg13g2_buf_1 place6783 (.A(_05509_),
    .X(net6782));
 sg13g2_buf_1 place6784 (.A(net6784),
    .X(net6783));
 sg13g2_buf_1 place6785 (.A(net6793),
    .X(net6784));
 sg13g2_buf_1 place6786 (.A(net6787),
    .X(net6785));
 sg13g2_buf_1 place6787 (.A(net6787),
    .X(net6786));
 sg13g2_buf_1 place6788 (.A(net6788),
    .X(net6787));
 sg13g2_buf_1 place6789 (.A(net6793),
    .X(net6788));
 sg13g2_buf_1 place6790 (.A(net6793),
    .X(net6789));
 sg13g2_buf_1 place6791 (.A(net6792),
    .X(net6790));
 sg13g2_buf_1 place6792 (.A(net6792),
    .X(net6791));
 sg13g2_buf_1 place6793 (.A(net6793),
    .X(net6792));
 sg13g2_buf_1 place6794 (.A(_13161_),
    .X(net6793));
 sg13g2_buf_1 place6795 (.A(_09554_),
    .X(net6794));
 sg13g2_buf_1 place6796 (.A(_09539_),
    .X(net6795));
 sg13g2_buf_1 place6797 (.A(net6797),
    .X(net6796));
 sg13g2_buf_1 place6798 (.A(_09539_),
    .X(net6797));
 sg13g2_buf_1 place6799 (.A(_09403_),
    .X(net6798));
 sg13g2_buf_1 place6800 (.A(net6801),
    .X(net6799));
 sg13g2_buf_1 place6801 (.A(net6801),
    .X(net6800));
 sg13g2_buf_1 place6802 (.A(_09402_),
    .X(net6801));
 sg13g2_buf_1 place6803 (.A(_09402_),
    .X(net6802));
 sg13g2_buf_1 place6804 (.A(_09402_),
    .X(net6803));
 sg13g2_buf_1 place6805 (.A(net6806),
    .X(net6804));
 sg13g2_buf_1 place6806 (.A(net6806),
    .X(net6805));
 sg13g2_buf_1 place6807 (.A(_08701_),
    .X(net6806));
 sg13g2_buf_1 place6808 (.A(net6808),
    .X(net6807));
 sg13g2_buf_1 place6809 (.A(net6811),
    .X(net6808));
 sg13g2_buf_1 place6810 (.A(net6810),
    .X(net6809));
 sg13g2_buf_1 place6811 (.A(net6811),
    .X(net6810));
 sg13g2_buf_1 place6812 (.A(net6812),
    .X(net6811));
 sg13g2_buf_1 place6813 (.A(_08700_),
    .X(net6812));
 sg13g2_buf_1 place6814 (.A(net6823),
    .X(net6813));
 sg13g2_buf_1 place6815 (.A(net6823),
    .X(net6814));
 sg13g2_buf_1 place6816 (.A(net6816),
    .X(net6815));
 sg13g2_buf_1 place6817 (.A(net6819),
    .X(net6816));
 sg13g2_buf_1 place6818 (.A(net6819),
    .X(net6817));
 sg13g2_buf_1 place6819 (.A(net6819),
    .X(net6818));
 sg13g2_buf_1 place6820 (.A(net6823),
    .X(net6819));
 sg13g2_buf_1 place6821 (.A(net6822),
    .X(net6820));
 sg13g2_buf_1 place6822 (.A(net6822),
    .X(net6821));
 sg13g2_buf_1 place6823 (.A(net6823),
    .X(net6822));
 sg13g2_buf_1 place6824 (.A(_08660_),
    .X(net6823));
 sg13g2_buf_1 place6825 (.A(_06944_),
    .X(net6824));
 sg13g2_buf_1 place6826 (.A(net6826),
    .X(net6825));
 sg13g2_buf_1 place6827 (.A(_06802_),
    .X(net6826));
 sg13g2_buf_1 place6828 (.A(_06027_),
    .X(net6827));
 sg13g2_buf_1 place6829 (.A(_05995_),
    .X(net6828));
 sg13g2_buf_1 place6830 (.A(_05743_),
    .X(net6829));
 sg13g2_buf_1 place6831 (.A(_05507_),
    .X(net6830));
 sg13g2_buf_1 place6832 (.A(_04813_),
    .X(net6831));
 sg13g2_buf_1 place6833 (.A(net6837),
    .X(net6832));
 sg13g2_buf_1 place6834 (.A(net6837),
    .X(net6833));
 sg13g2_buf_1 place6835 (.A(net6835),
    .X(net6834));
 sg13g2_buf_1 place6836 (.A(net6837),
    .X(net6835));
 sg13g2_buf_1 place6837 (.A(net6837),
    .X(net6836));
 sg13g2_buf_1 place6838 (.A(_09540_),
    .X(net6837));
 sg13g2_buf_1 place6839 (.A(net6839),
    .X(net6838));
 sg13g2_buf_1 place6840 (.A(net6840),
    .X(net6839));
 sg13g2_buf_1 place6841 (.A(net6841),
    .X(net6840));
 sg13g2_buf_1 place6842 (.A(_09540_),
    .X(net6841));
 sg13g2_buf_1 place6843 (.A(net6843),
    .X(net6842));
 sg13g2_buf_1 place6844 (.A(_09416_),
    .X(net6843));
 sg13g2_buf_1 place6845 (.A(net6847),
    .X(net6844));
 sg13g2_buf_1 place6846 (.A(net6846),
    .X(net6845));
 sg13g2_buf_1 place6847 (.A(net6847),
    .X(net6846));
 sg13g2_buf_1 place6848 (.A(_09409_),
    .X(net6847));
 sg13g2_buf_1 place6849 (.A(net6851),
    .X(net6848));
 sg13g2_buf_1 place6850 (.A(net6850),
    .X(net6849));
 sg13g2_buf_1 place6851 (.A(net6851),
    .X(net6850));
 sg13g2_buf_1 place6852 (.A(_09408_),
    .X(net6851));
 sg13g2_buf_1 place6853 (.A(_08659_),
    .X(net6852));
 sg13g2_buf_1 place6854 (.A(net6854),
    .X(net6853));
 sg13g2_buf_1 place6855 (.A(net6855),
    .X(net6854));
 sg13g2_buf_1 place6856 (.A(_07089_),
    .X(net6855));
 sg13g2_buf_1 place6857 (.A(net6857),
    .X(net6856));
 sg13g2_buf_1 place6858 (.A(_07089_),
    .X(net6857));
 sg13g2_buf_1 place6859 (.A(_05956_),
    .X(net6858));
 sg13g2_buf_1 place6860 (.A(_05820_),
    .X(net6859));
 sg13g2_buf_1 place6861 (.A(_05724_),
    .X(net6860));
 sg13g2_buf_1 place6862 (.A(_05505_),
    .X(net6861));
 sg13g2_buf_1 place6863 (.A(net6868),
    .X(net6862));
 sg13g2_buf_1 place6864 (.A(net6868),
    .X(net6863));
 sg13g2_buf_1 place6865 (.A(net6865),
    .X(net6864));
 sg13g2_buf_1 place6866 (.A(net6868),
    .X(net6865));
 sg13g2_buf_1 place6867 (.A(net6868),
    .X(net6866));
 sg13g2_buf_1 place6868 (.A(net6868),
    .X(net6867));
 sg13g2_buf_1 place6869 (.A(_09541_),
    .X(net6868));
 sg13g2_buf_1 place6870 (.A(net6870),
    .X(net6869));
 sg13g2_buf_1 place6871 (.A(net6871),
    .X(net6870));
 sg13g2_buf_1 place6872 (.A(_09541_),
    .X(net6871));
 sg13g2_buf_1 place6873 (.A(net6873),
    .X(net6872));
 sg13g2_buf_1 place6874 (.A(net6874),
    .X(net6873));
 sg13g2_buf_1 place6875 (.A(net6877),
    .X(net6874));
 sg13g2_buf_1 place6876 (.A(net6876),
    .X(net6875));
 sg13g2_buf_1 place6877 (.A(net6877),
    .X(net6876));
 sg13g2_buf_1 place6878 (.A(_09417_),
    .X(net6877));
 sg13g2_buf_1 place6879 (.A(net6879),
    .X(net6878));
 sg13g2_buf_1 place6880 (.A(_09394_),
    .X(net6879));
 sg13g2_buf_1 place6881 (.A(_09394_),
    .X(net6880));
 sg13g2_buf_1 place6882 (.A(net6882),
    .X(net6881));
 sg13g2_buf_1 place6883 (.A(_07679_),
    .X(net6882));
 sg13g2_buf_1 place6884 (.A(_07671_),
    .X(net6883));
 sg13g2_buf_1 place6885 (.A(net6885),
    .X(net6884));
 sg13g2_buf_1 place6886 (.A(_07671_),
    .X(net6885));
 sg13g2_buf_1 place6887 (.A(_07671_),
    .X(net6886));
 sg13g2_buf_1 place6888 (.A(_06811_),
    .X(net6887));
 sg13g2_buf_1 place6889 (.A(_06787_),
    .X(net6888));
 sg13g2_buf_1 place6890 (.A(_06215_),
    .X(net6889));
 sg13g2_buf_1 place6891 (.A(_05938_),
    .X(net6890));
 sg13g2_buf_1 place6892 (.A(_05835_),
    .X(net6891));
 sg13g2_buf_1 place6893 (.A(net6893),
    .X(net6892));
 sg13g2_buf_1 place6894 (.A(_05726_),
    .X(net6893));
 sg13g2_buf_1 place6895 (.A(_05725_),
    .X(net6894));
 sg13g2_buf_1 place6896 (.A(_05578_),
    .X(net6895));
 sg13g2_buf_1 place6897 (.A(_05572_),
    .X(net6896));
 sg13g2_buf_1 place6898 (.A(_05418_),
    .X(net6897));
 sg13g2_buf_1 place6899 (.A(_04627_),
    .X(net6898));
 sg13g2_buf_1 place6900 (.A(_14748_),
    .X(net6899));
 sg13g2_buf_1 place6901 (.A(_10789_),
    .X(net6900));
 sg13g2_buf_1 place6902 (.A(_10788_),
    .X(net6901));
 sg13g2_buf_1 place6903 (.A(_09994_),
    .X(net6902));
 sg13g2_buf_1 place6904 (.A(_09945_),
    .X(net6903));
 sg13g2_buf_1 place6905 (.A(net6905),
    .X(net6904));
 sg13g2_buf_1 place6906 (.A(_09387_),
    .X(net6905));
 sg13g2_buf_1 place6907 (.A(net6907),
    .X(net6906));
 sg13g2_buf_1 place6908 (.A(_09387_),
    .X(net6907));
 sg13g2_buf_1 place6909 (.A(net6909),
    .X(net6908));
 sg13g2_buf_1 place6910 (.A(net6912),
    .X(net6909));
 sg13g2_buf_1 place6911 (.A(net6911),
    .X(net6910));
 sg13g2_buf_1 place6912 (.A(net6912),
    .X(net6911));
 sg13g2_buf_1 place6913 (.A(_09386_),
    .X(net6912));
 sg13g2_buf_1 place6914 (.A(net6916),
    .X(net6913));
 sg13g2_buf_1 place6915 (.A(net6915),
    .X(net6914));
 sg13g2_buf_1 place6916 (.A(net6916),
    .X(net6915));
 sg13g2_buf_1 place6917 (.A(_08874_),
    .X(net6916));
 sg13g2_buf_1 place6918 (.A(_08251_),
    .X(net6917));
 sg13g2_buf_1 place6919 (.A(net6919),
    .X(net6918));
 sg13g2_buf_1 place6920 (.A(_08251_),
    .X(net6919));
 sg13g2_buf_1 place6921 (.A(net6921),
    .X(net6920));
 sg13g2_buf_1 place6922 (.A(net6922),
    .X(net6921));
 sg13g2_buf_1 place6923 (.A(_07704_),
    .X(net6922));
 sg13g2_buf_1 place6924 (.A(net6924),
    .X(net6923));
 sg13g2_buf_1 place6925 (.A(net6925),
    .X(net6924));
 sg13g2_buf_1 place6926 (.A(_07690_),
    .X(net6925));
 sg13g2_buf_1 place6927 (.A(net6927),
    .X(net6926));
 sg13g2_buf_1 place6928 (.A(_07686_),
    .X(net6927));
 sg13g2_buf_1 place6929 (.A(net6929),
    .X(net6928));
 sg13g2_buf_1 place6930 (.A(_07686_),
    .X(net6929));
 sg13g2_buf_1 place6931 (.A(net6931),
    .X(net6930));
 sg13g2_buf_1 place6932 (.A(net6932),
    .X(net6931));
 sg13g2_buf_1 place6933 (.A(_06786_),
    .X(net6932));
 sg13g2_buf_1 place6934 (.A(_05792_),
    .X(net6933));
 sg13g2_buf_1 place6935 (.A(_05498_),
    .X(net6934));
 sg13g2_buf_1 place6936 (.A(net6936),
    .X(net6935));
 sg13g2_buf_1 place6937 (.A(net6939),
    .X(net6936));
 sg13g2_buf_1 place6938 (.A(net6938),
    .X(net6937));
 sg13g2_buf_1 place6939 (.A(net6939),
    .X(net6938));
 sg13g2_buf_1 place6940 (.A(_05185_),
    .X(net6939));
 sg13g2_buf_1 place6941 (.A(net6942),
    .X(net6940));
 sg13g2_buf_1 place6942 (.A(net6942),
    .X(net6941));
 sg13g2_buf_1 place6943 (.A(net6943),
    .X(net6942));
 sg13g2_buf_1 place6944 (.A(_05184_),
    .X(net6943));
 sg13g2_buf_1 place6945 (.A(net6945),
    .X(net6944));
 sg13g2_buf_1 place6946 (.A(_05184_),
    .X(net6945));
 sg13g2_buf_1 place6947 (.A(_04556_),
    .X(net6946));
 sg13g2_buf_1 place6948 (.A(_04294_),
    .X(net6947));
 sg13g2_buf_1 place6949 (.A(_13840_),
    .X(net6948));
 sg13g2_buf_1 place6950 (.A(_12822_),
    .X(net6949));
 sg13g2_buf_1 place6951 (.A(net6951),
    .X(net6950));
 sg13g2_buf_1 place6952 (.A(_12819_),
    .X(net6951));
 sg13g2_buf_1 place6953 (.A(net6953),
    .X(net6952));
 sg13g2_buf_1 place6954 (.A(_11682_),
    .X(net6953));
 sg13g2_buf_1 place6955 (.A(net6958),
    .X(net6954));
 sg13g2_buf_1 place6956 (.A(net6956),
    .X(net6955));
 sg13g2_buf_1 place6957 (.A(net6957),
    .X(net6956));
 sg13g2_buf_1 place6958 (.A(net6958),
    .X(net6957));
 sg13g2_buf_1 place6959 (.A(_09400_),
    .X(net6958));
 sg13g2_buf_1 place6960 (.A(net6960),
    .X(net6959));
 sg13g2_buf_1 place6961 (.A(_09400_),
    .X(net6960));
 sg13g2_buf_1 place6962 (.A(net6963),
    .X(net6961));
 sg13g2_buf_1 place6963 (.A(net6963),
    .X(net6962));
 sg13g2_buf_1 place6964 (.A(net6964),
    .X(net6963));
 sg13g2_buf_1 place6965 (.A(_09399_),
    .X(net6964));
 sg13g2_buf_1 place6966 (.A(net6969),
    .X(net6965));
 sg13g2_buf_1 place6967 (.A(net6968),
    .X(net6966));
 sg13g2_buf_1 place6968 (.A(net6968),
    .X(net6967));
 sg13g2_buf_1 place6969 (.A(net6969),
    .X(net6968));
 sg13g2_buf_1 place6970 (.A(_09399_),
    .X(net6969));
 sg13g2_buf_1 place6971 (.A(net6971),
    .X(net6970));
 sg13g2_buf_1 place6972 (.A(_09390_),
    .X(net6971));
 sg13g2_buf_1 place6973 (.A(_09390_),
    .X(net6972));
 sg13g2_buf_1 place6974 (.A(net6976),
    .X(net6973));
 sg13g2_buf_1 place6975 (.A(net6976),
    .X(net6974));
 sg13g2_buf_1 place6976 (.A(net6976),
    .X(net6975));
 sg13g2_buf_1 place6977 (.A(net6977),
    .X(net6976));
 sg13g2_buf_1 place6978 (.A(_08873_),
    .X(net6977));
 sg13g2_buf_1 place6979 (.A(net6979),
    .X(net6978));
 sg13g2_buf_1 place6980 (.A(net6980),
    .X(net6979));
 sg13g2_buf_1 place6981 (.A(net6981),
    .X(net6980));
 sg13g2_buf_1 place6982 (.A(_08228_),
    .X(net6981));
 sg13g2_buf_1 place6983 (.A(_08222_),
    .X(net6982));
 sg13g2_buf_1 place6984 (.A(net6984),
    .X(net6983));
 sg13g2_buf_1 place6985 (.A(_08222_),
    .X(net6984));
 sg13g2_buf_1 place6986 (.A(_07762_),
    .X(net6985));
 sg13g2_buf_1 place6987 (.A(net6987),
    .X(net6986));
 sg13g2_buf_1 place6988 (.A(net6988),
    .X(net6987));
 sg13g2_buf_1 place6989 (.A(_07762_),
    .X(net6988));
 sg13g2_buf_1 place6990 (.A(_05924_),
    .X(net6989));
 sg13g2_buf_1 place6991 (.A(_05488_),
    .X(net6990));
 sg13g2_buf_1 place6992 (.A(_05182_),
    .X(net6991));
 sg13g2_buf_1 place6993 (.A(_05176_),
    .X(net6992));
 sg13g2_buf_1 place6994 (.A(_05027_),
    .X(net6993));
 sg13g2_buf_1 place6995 (.A(_05027_),
    .X(net6994));
 sg13g2_buf_1 place6996 (.A(net6996),
    .X(net6995));
 sg13g2_buf_1 place6997 (.A(_05027_),
    .X(net6996));
 sg13g2_buf_1 place6998 (.A(_04919_),
    .X(net6997));
 sg13g2_buf_1 place6999 (.A(net6999),
    .X(net6998));
 sg13g2_buf_1 place7000 (.A(_04919_),
    .X(net6999));
 sg13g2_buf_1 place7001 (.A(net7002),
    .X(net7000));
 sg13g2_buf_1 place7002 (.A(net7002),
    .X(net7001));
 sg13g2_buf_1 place7003 (.A(net7004),
    .X(net7002));
 sg13g2_buf_1 place7004 (.A(net7004),
    .X(net7003));
 sg13g2_buf_2 place7005 (.A(_04918_),
    .X(net7004));
 sg13g2_buf_1 place7006 (.A(_04916_),
    .X(net7005));
 sg13g2_buf_1 place7007 (.A(_03805_),
    .X(net7006));
 sg13g2_buf_1 place7008 (.A(_03800_),
    .X(net7007));
 sg13g2_buf_1 place7009 (.A(_03789_),
    .X(net7008));
 sg13g2_buf_1 place7010 (.A(_03779_),
    .X(net7009));
 sg13g2_buf_1 place7011 (.A(_03774_),
    .X(net7010));
 sg13g2_buf_1 place7012 (.A(_03769_),
    .X(net7011));
 sg13g2_buf_1 place7013 (.A(_03749_),
    .X(net7012));
 sg13g2_buf_1 place7014 (.A(_03744_),
    .X(net7013));
 sg13g2_buf_1 place7015 (.A(_03739_),
    .X(net7014));
 sg13g2_buf_1 place7016 (.A(_03735_),
    .X(net7015));
 sg13g2_buf_1 place7017 (.A(_03724_),
    .X(net7016));
 sg13g2_buf_1 place7018 (.A(_03719_),
    .X(net7017));
 sg13g2_buf_1 place7019 (.A(_03714_),
    .X(net7018));
 sg13g2_buf_1 place7020 (.A(_03709_),
    .X(net7019));
 sg13g2_buf_1 place7021 (.A(_03704_),
    .X(net7020));
 sg13g2_buf_1 place7022 (.A(_03699_),
    .X(net7021));
 sg13g2_buf_1 place7023 (.A(_03694_),
    .X(net7022));
 sg13g2_buf_1 place7024 (.A(_03689_),
    .X(net7023));
 sg13g2_buf_1 place7025 (.A(_03684_),
    .X(net7024));
 sg13g2_buf_1 place7026 (.A(_03679_),
    .X(net7025));
 sg13g2_buf_1 place7027 (.A(_03674_),
    .X(net7026));
 sg13g2_buf_1 place7028 (.A(_03668_),
    .X(net7027));
 sg13g2_buf_1 place7029 (.A(_03662_),
    .X(net7028));
 sg13g2_buf_1 place7030 (.A(_03657_),
    .X(net7029));
 sg13g2_buf_1 place7031 (.A(_03123_),
    .X(net7030));
 sg13g2_buf_1 place7032 (.A(net7032),
    .X(net7031));
 sg13g2_buf_1 place7033 (.A(_02254_),
    .X(net7032));
 sg13g2_buf_1 place7034 (.A(_02173_),
    .X(net7033));
 sg13g2_buf_1 place7035 (.A(net7035),
    .X(net7034));
 sg13g2_buf_1 place7036 (.A(net7036),
    .X(net7035));
 sg13g2_buf_1 place7037 (.A(_13895_),
    .X(net7036));
 sg13g2_buf_1 place7038 (.A(net7038),
    .X(net7037));
 sg13g2_buf_1 place7039 (.A(_13895_),
    .X(net7038));
 sg13g2_buf_1 place7040 (.A(_13410_),
    .X(net7039));
 sg13g2_buf_1 place7041 (.A(net7043),
    .X(net7040));
 sg13g2_buf_1 place7042 (.A(net7043),
    .X(net7041));
 sg13g2_buf_1 place7043 (.A(net7043),
    .X(net7042));
 sg13g2_buf_1 place7044 (.A(_08687_),
    .X(net7043));
 sg13g2_buf_1 place7045 (.A(net7045),
    .X(net7044));
 sg13g2_buf_1 place7046 (.A(_08687_),
    .X(net7045));
 sg13g2_buf_1 place7047 (.A(_08126_),
    .X(net7046));
 sg13g2_buf_1 place7048 (.A(net7048),
    .X(net7047));
 sg13g2_buf_1 place7049 (.A(net7049),
    .X(net7048));
 sg13g2_buf_1 place7050 (.A(_07696_),
    .X(net7049));
 sg13g2_buf_1 place7051 (.A(_07228_),
    .X(net7050));
 sg13g2_buf_1 place7052 (.A(_07215_),
    .X(net7051));
 sg13g2_buf_1 place7053 (.A(_05355_),
    .X(net7052));
 sg13g2_buf_1 place7054 (.A(_05026_),
    .X(net7053));
 sg13g2_buf_1 place7055 (.A(net7056),
    .X(net7054));
 sg13g2_buf_1 place7056 (.A(net7056),
    .X(net7055));
 sg13g2_buf_1 place7057 (.A(net7058),
    .X(net7056));
 sg13g2_buf_1 place7058 (.A(net7058),
    .X(net7057));
 sg13g2_buf_1 place7059 (.A(_05026_),
    .X(net7058));
 sg13g2_buf_1 place7060 (.A(_05025_),
    .X(net7059));
 sg13g2_buf_1 place7061 (.A(_05025_),
    .X(net7060));
 sg13g2_buf_1 place7062 (.A(_04793_),
    .X(net7061));
 sg13g2_buf_1 place7063 (.A(net7063),
    .X(net7062));
 sg13g2_buf_1 place7064 (.A(_04743_),
    .X(net7063));
 sg13g2_buf_1 place7065 (.A(_04743_),
    .X(net7064));
 sg13g2_buf_1 place7066 (.A(_04734_),
    .X(net7065));
 sg13g2_buf_1 place7067 (.A(_04131_),
    .X(net7066));
 sg13g2_buf_2 place7068 (.A(_04130_),
    .X(net7067));
 sg13g2_buf_1 place7069 (.A(_04015_),
    .X(net7068));
 sg13g2_buf_1 place7070 (.A(net7070),
    .X(net7069));
 sg13g2_buf_1 place7071 (.A(_03835_),
    .X(net7070));
 sg13g2_buf_1 place7072 (.A(_03826_),
    .X(net7071));
 sg13g2_buf_1 place7073 (.A(_03649_),
    .X(net7072));
 sg13g2_buf_1 place7074 (.A(_02852_),
    .X(net7073));
 sg13g2_buf_2 place7075 (.A(_13803_),
    .X(net7074));
 sg13g2_buf_1 place7076 (.A(_13570_),
    .X(net7075));
 sg13g2_buf_1 place7077 (.A(_10370_),
    .X(net7076));
 sg13g2_buf_2 place7078 (.A(_09924_),
    .X(net7077));
 sg13g2_buf_1 place7079 (.A(_09321_),
    .X(net7078));
 sg13g2_buf_1 place7080 (.A(_09320_),
    .X(net7079));
 sg13g2_buf_1 place7081 (.A(_08753_),
    .X(net7080));
 sg13g2_buf_1 place7082 (.A(_08742_),
    .X(net7081));
 sg13g2_buf_1 place7083 (.A(_08742_),
    .X(net7082));
 sg13g2_buf_1 place7084 (.A(_08709_),
    .X(net7083));
 sg13g2_buf_1 place7085 (.A(net7089),
    .X(net7084));
 sg13g2_buf_1 place7086 (.A(net7086),
    .X(net7085));
 sg13g2_buf_1 place7087 (.A(net7089),
    .X(net7086));
 sg13g2_buf_1 place7088 (.A(net7089),
    .X(net7087));
 sg13g2_buf_1 place7089 (.A(net7089),
    .X(net7088));
 sg13g2_buf_1 place7090 (.A(_08707_),
    .X(net7089));
 sg13g2_buf_1 place7091 (.A(net7091),
    .X(net7090));
 sg13g2_buf_1 place7092 (.A(net7092),
    .X(net7091));
 sg13g2_buf_1 place7093 (.A(_08695_),
    .X(net7092));
 sg13g2_buf_1 place7094 (.A(net7095),
    .X(net7093));
 sg13g2_buf_1 place7095 (.A(net7095),
    .X(net7094));
 sg13g2_buf_1 place7096 (.A(_08695_),
    .X(net7095));
 sg13g2_buf_1 place7097 (.A(net7097),
    .X(net7096));
 sg13g2_buf_1 place7098 (.A(_08694_),
    .X(net7097));
 sg13g2_buf_1 place7099 (.A(net7100),
    .X(net7098));
 sg13g2_buf_1 place7100 (.A(net7100),
    .X(net7099));
 sg13g2_buf_1 place7101 (.A(_08690_),
    .X(net7100));
 sg13g2_buf_1 place7102 (.A(_08690_),
    .X(net7101));
 sg13g2_buf_1 place7103 (.A(_08688_),
    .X(net7102));
 sg13g2_buf_1 place7104 (.A(_08586_),
    .X(net7103));
 sg13g2_buf_1 place7105 (.A(_08195_),
    .X(net7104));
 sg13g2_buf_1 place7106 (.A(_06775_),
    .X(net7105));
 sg13g2_buf_1 place7107 (.A(net7108),
    .X(net7106));
 sg13g2_buf_1 place7108 (.A(net7108),
    .X(net7107));
 sg13g2_buf_1 place7109 (.A(_06568_),
    .X(net7108));
 sg13g2_buf_1 place7110 (.A(_06363_),
    .X(net7109));
 sg13g2_buf_1 place7111 (.A(_06160_),
    .X(net7110));
 sg13g2_buf_1 place7112 (.A(_06121_),
    .X(net7111));
 sg13g2_buf_1 place7113 (.A(_06010_),
    .X(net7112));
 sg13g2_buf_1 place7114 (.A(_05754_),
    .X(net7113));
 sg13g2_buf_1 place7115 (.A(net7116),
    .X(net7114));
 sg13g2_buf_1 place7116 (.A(net7116),
    .X(net7115));
 sg13g2_buf_1 place7117 (.A(_04798_),
    .X(net7116));
 sg13g2_buf_1 place7118 (.A(_04798_),
    .X(net7117));
 sg13g2_buf_1 place7119 (.A(_04797_),
    .X(net7118));
 sg13g2_buf_1 place7120 (.A(_04797_),
    .X(net7119));
 sg13g2_buf_1 place7121 (.A(_04794_),
    .X(net7120));
 sg13g2_buf_1 place7122 (.A(_04742_),
    .X(net7121));
 sg13g2_buf_1 place7123 (.A(_04742_),
    .X(net7122));
 sg13g2_buf_1 place7124 (.A(net7124),
    .X(net7123));
 sg13g2_buf_1 place7125 (.A(_04742_),
    .X(net7124));
 sg13g2_buf_1 place7126 (.A(net7126),
    .X(net7125));
 sg13g2_buf_1 place7127 (.A(net7129),
    .X(net7126));
 sg13g2_buf_1 place7128 (.A(net7128),
    .X(net7127));
 sg13g2_buf_1 place7129 (.A(net7129),
    .X(net7128));
 sg13g2_buf_1 place7130 (.A(_04736_),
    .X(net7129));
 sg13g2_buf_1 place7131 (.A(net7132),
    .X(net7130));
 sg13g2_buf_1 place7132 (.A(net7132),
    .X(net7131));
 sg13g2_buf_1 place7133 (.A(_04678_),
    .X(net7132));
 sg13g2_buf_1 place7134 (.A(_04677_),
    .X(net7133));
 sg13g2_buf_2 place7135 (.A(net7135),
    .X(net7134));
 sg13g2_buf_1 place7136 (.A(_04649_),
    .X(net7135));
 sg13g2_buf_1 place7137 (.A(net7137),
    .X(net7136));
 sg13g2_buf_1 place7138 (.A(net7139),
    .X(net7137));
 sg13g2_buf_1 place7139 (.A(net7139),
    .X(net7138));
 sg13g2_buf_1 place7140 (.A(_04576_),
    .X(net7139));
 sg13g2_buf_1 place7141 (.A(net7143),
    .X(net7140));
 sg13g2_buf_1 place7142 (.A(net7142),
    .X(net7141));
 sg13g2_buf_1 place7143 (.A(net7143),
    .X(net7142));
 sg13g2_buf_2 place7144 (.A(_04560_),
    .X(net7143));
 sg13g2_buf_1 place7145 (.A(net7147),
    .X(net7144));
 sg13g2_buf_1 place7146 (.A(net7146),
    .X(net7145));
 sg13g2_buf_1 place7147 (.A(net7147),
    .X(net7146));
 sg13g2_buf_2 place7148 (.A(_04503_),
    .X(net7147));
 sg13g2_buf_1 place7149 (.A(net7149),
    .X(net7148));
 sg13g2_buf_1 place7150 (.A(net7151),
    .X(net7149));
 sg13g2_buf_1 place7151 (.A(net7151),
    .X(net7150));
 sg13g2_buf_2 place7152 (.A(_04446_),
    .X(net7151));
 sg13g2_buf_1 place7153 (.A(net7153),
    .X(net7152));
 sg13g2_buf_1 place7154 (.A(net7155),
    .X(net7153));
 sg13g2_buf_1 place7155 (.A(net7155),
    .X(net7154));
 sg13g2_buf_1 place7156 (.A(_04414_),
    .X(net7155));
 sg13g2_buf_1 place7157 (.A(net7158),
    .X(net7156));
 sg13g2_buf_1 place7158 (.A(net7158),
    .X(net7157));
 sg13g2_buf_1 place7159 (.A(_04367_),
    .X(net7158));
 sg13g2_buf_2 place7160 (.A(net7161),
    .X(net7159));
 sg13g2_buf_1 place7161 (.A(net7161),
    .X(net7160));
 sg13g2_buf_2 place7162 (.A(_04336_),
    .X(net7161));
 sg13g2_buf_1 place7163 (.A(_04297_),
    .X(net7162));
 sg13g2_buf_1 place7164 (.A(net7165),
    .X(net7163));
 sg13g2_buf_1 place7165 (.A(net7165),
    .X(net7164));
 sg13g2_buf_1 place7166 (.A(_04297_),
    .X(net7165));
 sg13g2_buf_1 place7167 (.A(_04297_),
    .X(net7166));
 sg13g2_buf_1 place7168 (.A(net7172),
    .X(net7167));
 sg13g2_buf_1 place7169 (.A(net7172),
    .X(net7168));
 sg13g2_buf_1 place7170 (.A(net7172),
    .X(net7169));
 sg13g2_buf_1 place7171 (.A(net7171),
    .X(net7170));
 sg13g2_buf_1 place7172 (.A(net7172),
    .X(net7171));
 sg13g2_buf_2 place7173 (.A(_04243_),
    .X(net7172));
 sg13g2_buf_1 place7174 (.A(net7174),
    .X(net7173));
 sg13g2_buf_1 place7175 (.A(_04215_),
    .X(net7174));
 sg13g2_buf_1 place7176 (.A(_04215_),
    .X(net7175));
 sg13g2_buf_1 place7177 (.A(_04215_),
    .X(net7176));
 sg13g2_buf_1 place7178 (.A(net7180),
    .X(net7177));
 sg13g2_buf_1 place7179 (.A(net7179),
    .X(net7178));
 sg13g2_buf_2 place7180 (.A(net7180),
    .X(net7179));
 sg13g2_buf_8 place7181 (.A(_04178_),
    .X(net7180));
 sg13g2_buf_1 place7182 (.A(net7183),
    .X(net7181));
 sg13g2_buf_1 place7183 (.A(net7183),
    .X(net7182));
 sg13g2_buf_2 place7184 (.A(_04142_),
    .X(net7183));
 sg13g2_buf_1 place7185 (.A(net7187),
    .X(net7184));
 sg13g2_buf_1 place7186 (.A(net7186),
    .X(net7185));
 sg13g2_buf_1 place7187 (.A(net7187),
    .X(net7186));
 sg13g2_buf_4 place7188 (.X(net7187),
    .A(_04129_));
 sg13g2_buf_1 place7189 (.A(net7190),
    .X(net7188));
 sg13g2_buf_1 place7190 (.A(net7190),
    .X(net7189));
 sg13g2_buf_2 place7191 (.A(_04078_),
    .X(net7190));
 sg13g2_buf_1 place7192 (.A(net7194),
    .X(net7191));
 sg13g2_buf_1 place7193 (.A(net7194),
    .X(net7192));
 sg13g2_buf_1 place7194 (.A(net7194),
    .X(net7193));
 sg13g2_buf_2 place7195 (.A(_04041_),
    .X(net7194));
 sg13g2_buf_1 place7196 (.A(_04021_),
    .X(net7195));
 sg13g2_buf_1 place7197 (.A(net7197),
    .X(net7196));
 sg13g2_buf_1 place7198 (.A(_04021_),
    .X(net7197));
 sg13g2_buf_1 place7199 (.A(net7199),
    .X(net7198));
 sg13g2_buf_1 place7200 (.A(_03981_),
    .X(net7199));
 sg13g2_buf_1 place7201 (.A(_03981_),
    .X(net7200));
 sg13g2_buf_2 place7202 (.A(_03970_),
    .X(net7201));
 sg13g2_buf_1 place7203 (.A(net7203),
    .X(net7202));
 sg13g2_buf_1 place7204 (.A(_03970_),
    .X(net7203));
 sg13g2_buf_1 place7205 (.A(net7208),
    .X(net7204));
 sg13g2_buf_1 place7206 (.A(net7208),
    .X(net7205));
 sg13g2_buf_1 place7207 (.A(net7207),
    .X(net7206));
 sg13g2_buf_1 place7208 (.A(net7208),
    .X(net7207));
 sg13g2_buf_1 place7209 (.A(_03952_),
    .X(net7208));
 sg13g2_buf_1 place7210 (.A(_03931_),
    .X(net7209));
 sg13g2_buf_1 place7211 (.A(_03931_),
    .X(net7210));
 sg13g2_buf_1 place7212 (.A(_03908_),
    .X(net7211));
 sg13g2_buf_1 place7213 (.A(_03908_),
    .X(net7212));
 sg13g2_buf_1 place7214 (.A(net7214),
    .X(net7213));
 sg13g2_buf_1 place7215 (.A(net7216),
    .X(net7214));
 sg13g2_buf_1 place7216 (.A(net7216),
    .X(net7215));
 sg13g2_buf_2 place7217 (.A(_03904_),
    .X(net7216));
 sg13g2_buf_1 place7218 (.A(net7218),
    .X(net7217));
 sg13g2_buf_1 place7219 (.A(net7220),
    .X(net7218));
 sg13g2_buf_1 place7220 (.A(net7220),
    .X(net7219));
 sg13g2_buf_2 place7221 (.A(_03883_),
    .X(net7220));
 sg13g2_buf_1 place7222 (.A(net7224),
    .X(net7221));
 sg13g2_buf_1 place7223 (.A(net7223),
    .X(net7222));
 sg13g2_buf_1 place7224 (.A(net7224),
    .X(net7223));
 sg13g2_buf_1 place7225 (.A(_03869_),
    .X(net7224));
 sg13g2_buf_1 place7226 (.A(net7226),
    .X(net7225));
 sg13g2_buf_1 place7227 (.A(_03862_),
    .X(net7226));
 sg13g2_buf_1 place7228 (.A(net7228),
    .X(net7227));
 sg13g2_buf_1 place7229 (.A(_03862_),
    .X(net7228));
 sg13g2_buf_1 place7230 (.A(_03846_),
    .X(net7229));
 sg13g2_buf_1 place7231 (.A(_03846_),
    .X(net7230));
 sg13g2_buf_1 place7232 (.A(_03846_),
    .X(net7231));
 sg13g2_buf_1 place7233 (.A(_03846_),
    .X(net7232));
 sg13g2_buf_1 place7234 (.A(_03846_),
    .X(net7233));
 sg13g2_buf_1 place7235 (.A(net7239),
    .X(net7234));
 sg13g2_buf_1 place7236 (.A(net7239),
    .X(net7235));
 sg13g2_buf_1 place7237 (.A(net7239),
    .X(net7236));
 sg13g2_buf_1 place7238 (.A(net7238),
    .X(net7237));
 sg13g2_buf_1 place7239 (.A(net7239),
    .X(net7238));
 sg13g2_buf_1 place7240 (.A(net7240),
    .X(net7239));
 sg13g2_buf_2 place7241 (.A(_03839_),
    .X(net7240));
 sg13g2_buf_1 place7242 (.A(_03834_),
    .X(net7241));
 sg13g2_buf_1 place7243 (.A(net7246),
    .X(net7242));
 sg13g2_buf_1 place7244 (.A(net7246),
    .X(net7243));
 sg13g2_buf_1 place7245 (.A(net7246),
    .X(net7244));
 sg13g2_buf_1 place7246 (.A(net7246),
    .X(net7245));
 sg13g2_buf_4 place7247 (.X(net7246),
    .A(_03829_));
 sg13g2_buf_1 place7248 (.A(net7248),
    .X(net7247));
 sg13g2_buf_1 place7249 (.A(net7250),
    .X(net7248));
 sg13g2_buf_1 place7250 (.A(net7250),
    .X(net7249));
 sg13g2_buf_1 place7251 (.A(_03825_),
    .X(net7250));
 sg13g2_buf_1 place7252 (.A(_03653_),
    .X(net7251));
 sg13g2_buf_1 place7253 (.A(net7254),
    .X(net7252));
 sg13g2_buf_1 place7254 (.A(net7254),
    .X(net7253));
 sg13g2_buf_1 place7255 (.A(_03653_),
    .X(net7254));
 sg13g2_buf_1 place7256 (.A(net7256),
    .X(net7255));
 sg13g2_buf_1 place7257 (.A(net7258),
    .X(net7256));
 sg13g2_buf_1 place7258 (.A(net7258),
    .X(net7257));
 sg13g2_buf_1 place7259 (.A(_03646_),
    .X(net7258));
 sg13g2_buf_1 place7260 (.A(_03538_),
    .X(net7259));
 sg13g2_buf_1 place7261 (.A(_03404_),
    .X(net7260));
 sg13g2_buf_1 place7262 (.A(_02851_),
    .X(net7261));
 sg13g2_buf_1 place7263 (.A(_02779_),
    .X(net7262));
 sg13g2_buf_1 place7264 (.A(_02714_),
    .X(net7263));
 sg13g2_buf_1 place7265 (.A(_02534_),
    .X(net7264));
 sg13g2_buf_1 place7266 (.A(_02400_),
    .X(net7265));
 sg13g2_buf_1 place7267 (.A(_02325_),
    .X(net7266));
 sg13g2_buf_1 place7268 (.A(net7268),
    .X(net7267));
 sg13g2_buf_1 place7269 (.A(_02290_),
    .X(net7268));
 sg13g2_buf_1 place7270 (.A(_02253_),
    .X(net7269));
 sg13g2_buf_1 place7271 (.A(_02103_),
    .X(net7270));
 sg13g2_buf_2 place7272 (.A(_02030_),
    .X(net7271));
 sg13g2_buf_1 place7273 (.A(_15458_),
    .X(net7272));
 sg13g2_buf_1 place7274 (.A(_15072_),
    .X(net7273));
 sg13g2_buf_1 place7275 (.A(_14722_),
    .X(net7274));
 sg13g2_buf_1 place7276 (.A(_14252_),
    .X(net7275));
 sg13g2_buf_1 place7277 (.A(net7280),
    .X(net7276));
 sg13g2_buf_1 place7278 (.A(net7280),
    .X(net7277));
 sg13g2_buf_1 place7279 (.A(net7279),
    .X(net7278));
 sg13g2_buf_1 place7280 (.A(net7280),
    .X(net7279));
 sg13g2_buf_1 place7281 (.A(_13569_),
    .X(net7280));
 sg13g2_buf_1 place7282 (.A(_12788_),
    .X(net7281));
 sg13g2_buf_1 place7283 (.A(_12228_),
    .X(net7282));
 sg13g2_buf_1 place7284 (.A(_11147_),
    .X(net7283));
 sg13g2_buf_1 place7285 (.A(_09254_),
    .X(net7284));
 sg13g2_buf_1 place7286 (.A(_08662_),
    .X(net7285));
 sg13g2_buf_1 place7287 (.A(net7287),
    .X(net7286));
 sg13g2_buf_1 place7288 (.A(net7290),
    .X(net7287));
 sg13g2_buf_1 place7289 (.A(net7289),
    .X(net7288));
 sg13g2_buf_1 place7290 (.A(net7290),
    .X(net7289));
 sg13g2_buf_1 place7291 (.A(_08657_),
    .X(net7290));
 sg13g2_buf_1 place7292 (.A(_08641_),
    .X(net7291));
 sg13g2_buf_1 place7293 (.A(_08639_),
    .X(net7292));
 sg13g2_buf_1 place7294 (.A(net7295),
    .X(net7293));
 sg13g2_buf_1 place7295 (.A(net7295),
    .X(net7294));
 sg13g2_buf_1 place7296 (.A(net7296),
    .X(net7295));
 sg13g2_buf_1 place7297 (.A(_08202_),
    .X(net7296));
 sg13g2_buf_1 place7298 (.A(net7299),
    .X(net7297));
 sg13g2_buf_1 place7299 (.A(net7299),
    .X(net7298));
 sg13g2_buf_1 place7300 (.A(_08081_),
    .X(net7299));
 sg13g2_buf_1 place7301 (.A(_08081_),
    .X(net7300));
 sg13g2_buf_1 place7302 (.A(_07180_),
    .X(net7301));
 sg13g2_buf_1 place7303 (.A(_07179_),
    .X(net7302));
 sg13g2_buf_1 place7304 (.A(net7305),
    .X(net7303));
 sg13g2_buf_1 place7305 (.A(net7305),
    .X(net7304));
 sg13g2_buf_1 place7306 (.A(_07178_),
    .X(net7305));
 sg13g2_buf_1 place7307 (.A(_07134_),
    .X(net7306));
 sg13g2_buf_1 place7308 (.A(_07133_),
    .X(net7307));
 sg13g2_buf_1 place7309 (.A(_07130_),
    .X(net7308));
 sg13g2_buf_1 place7310 (.A(net7312),
    .X(net7309));
 sg13g2_buf_1 place7311 (.A(net7311),
    .X(net7310));
 sg13g2_buf_1 place7312 (.A(net7312),
    .X(net7311));
 sg13g2_buf_1 place7313 (.A(_06970_),
    .X(net7312));
 sg13g2_buf_1 place7314 (.A(_06778_),
    .X(net7313));
 sg13g2_buf_1 place7315 (.A(net7315),
    .X(net7314));
 sg13g2_buf_1 place7316 (.A(_05018_),
    .X(net7315));
 sg13g2_buf_1 place7317 (.A(net7317),
    .X(net7316));
 sg13g2_buf_1 place7318 (.A(_05018_),
    .X(net7317));
 sg13g2_buf_1 place7319 (.A(_04796_),
    .X(net7318));
 sg13g2_buf_1 place7320 (.A(net7324),
    .X(net7319));
 sg13g2_buf_1 place7321 (.A(net7323),
    .X(net7320));
 sg13g2_buf_1 place7322 (.A(net7322),
    .X(net7321));
 sg13g2_buf_1 place7323 (.A(net7323),
    .X(net7322));
 sg13g2_buf_1 place7324 (.A(net7324),
    .X(net7323));
 sg13g2_buf_1 place7325 (.A(_03819_),
    .X(net7324));
 sg13g2_buf_1 place7326 (.A(_03818_),
    .X(net7325));
 sg13g2_buf_1 place7327 (.A(net7327),
    .X(net7326));
 sg13g2_buf_1 place7328 (.A(_03817_),
    .X(net7327));
 sg13g2_buf_1 place7329 (.A(_03574_),
    .X(net7328));
 sg13g2_buf_1 place7330 (.A(_03505_),
    .X(net7329));
 sg13g2_buf_2 place7331 (.A(_03472_),
    .X(net7330));
 sg13g2_buf_1 place7332 (.A(_03437_),
    .X(net7331));
 sg13g2_buf_1 place7333 (.A(_03292_),
    .X(net7332));
 sg13g2_buf_1 place7334 (.A(_03226_),
    .X(net7333));
 sg13g2_buf_1 place7335 (.A(_03158_),
    .X(net7334));
 sg13g2_buf_1 place7336 (.A(_03121_),
    .X(net7335));
 sg13g2_buf_1 place7337 (.A(_03085_),
    .X(net7336));
 sg13g2_buf_1 place7338 (.A(_03052_),
    .X(net7337));
 sg13g2_buf_1 place7339 (.A(_03018_),
    .X(net7338));
 sg13g2_buf_1 place7340 (.A(_02985_),
    .X(net7339));
 sg13g2_buf_1 place7341 (.A(_02951_),
    .X(net7340));
 sg13g2_buf_1 place7342 (.A(_02886_),
    .X(net7341));
 sg13g2_buf_1 place7343 (.A(_02849_),
    .X(net7342));
 sg13g2_buf_1 place7344 (.A(_02746_),
    .X(net7343));
 sg13g2_buf_1 place7345 (.A(_02682_),
    .X(net7344));
 sg13g2_buf_1 place7346 (.A(_02651_),
    .X(net7345));
 sg13g2_buf_1 place7347 (.A(_02615_),
    .X(net7346));
 sg13g2_buf_1 place7348 (.A(_02503_),
    .X(net7347));
 sg13g2_buf_1 place7349 (.A(_02206_),
    .X(net7348));
 sg13g2_buf_1 place7350 (.A(_02140_),
    .X(net7349));
 sg13g2_buf_1 place7351 (.A(_13660_),
    .X(net7350));
 sg13g2_buf_1 place7352 (.A(_13660_),
    .X(net7351));
 sg13g2_buf_1 place7353 (.A(net7353),
    .X(net7352));
 sg13g2_buf_1 place7354 (.A(_09275_),
    .X(net7353));
 sg13g2_buf_1 place7355 (.A(_09275_),
    .X(net7354));
 sg13g2_buf_1 place7356 (.A(net7359),
    .X(net7355));
 sg13g2_buf_1 place7357 (.A(net7359),
    .X(net7356));
 sg13g2_buf_1 place7358 (.A(net7358),
    .X(net7357));
 sg13g2_buf_1 place7359 (.A(net7359),
    .X(net7358));
 sg13g2_buf_1 place7360 (.A(net7362),
    .X(net7359));
 sg13g2_buf_1 place7361 (.A(net7362),
    .X(net7360));
 sg13g2_buf_1 place7362 (.A(net7362),
    .X(net7361));
 sg13g2_buf_1 place7363 (.A(_08636_),
    .X(net7362));
 sg13g2_buf_1 place7364 (.A(_08614_),
    .X(net7363));
 sg13g2_buf_1 place7365 (.A(_08250_),
    .X(net7364));
 sg13g2_buf_1 place7366 (.A(net7366),
    .X(net7365));
 sg13g2_buf_1 place7367 (.A(_08250_),
    .X(net7366));
 sg13g2_buf_1 place7368 (.A(net7368),
    .X(net7367));
 sg13g2_buf_1 place7369 (.A(net7369),
    .X(net7368));
 sg13g2_buf_1 place7370 (.A(net7371),
    .X(net7369));
 sg13g2_buf_1 place7371 (.A(net7371),
    .X(net7370));
 sg13g2_buf_1 place7372 (.A(net7372),
    .X(net7371));
 sg13g2_buf_1 place7373 (.A(net7373),
    .X(net7372));
 sg13g2_buf_1 place7374 (.A(_08250_),
    .X(net7373));
 sg13g2_buf_1 place7375 (.A(net7375),
    .X(net7374));
 sg13g2_buf_1 place7376 (.A(net7376),
    .X(net7375));
 sg13g2_buf_1 place7377 (.A(_08250_),
    .X(net7376));
 sg13g2_buf_1 place7378 (.A(net7384),
    .X(net7377));
 sg13g2_buf_1 place7379 (.A(net7379),
    .X(net7378));
 sg13g2_buf_1 place7380 (.A(net7380),
    .X(net7379));
 sg13g2_buf_1 place7381 (.A(net7384),
    .X(net7380));
 sg13g2_buf_1 place7382 (.A(net7383),
    .X(net7381));
 sg13g2_buf_1 place7383 (.A(net7383),
    .X(net7382));
 sg13g2_buf_1 place7384 (.A(net7384),
    .X(net7383));
 sg13g2_buf_2 place7385 (.A(_08249_),
    .X(net7384));
 sg13g2_buf_1 place7386 (.A(_08239_),
    .X(net7385));
 sg13g2_buf_1 place7387 (.A(net7387),
    .X(net7386));
 sg13g2_buf_1 place7388 (.A(_07195_),
    .X(net7387));
 sg13g2_buf_1 place7389 (.A(_07194_),
    .X(net7388));
 sg13g2_buf_1 place7390 (.A(_07194_),
    .X(net7389));
 sg13g2_buf_1 place7391 (.A(_07129_),
    .X(net7390));
 sg13g2_buf_1 place7392 (.A(_07129_),
    .X(net7391));
 sg13g2_buf_1 place7393 (.A(_07128_),
    .X(net7392));
 sg13g2_buf_1 place7394 (.A(net7394),
    .X(net7393));
 sg13g2_buf_1 place7395 (.A(_07128_),
    .X(net7394));
 sg13g2_buf_1 place7396 (.A(net7397),
    .X(net7395));
 sg13g2_buf_1 place7397 (.A(net7397),
    .X(net7396));
 sg13g2_buf_1 place7398 (.A(_07121_),
    .X(net7397));
 sg13g2_buf_1 place7399 (.A(_07121_),
    .X(net7398));
 sg13g2_buf_1 place7400 (.A(net7400),
    .X(net7399));
 sg13g2_buf_1 place7401 (.A(_07115_),
    .X(net7400));
 sg13g2_buf_1 place7402 (.A(net7402),
    .X(net7401));
 sg13g2_buf_1 place7403 (.A(net7403),
    .X(net7402));
 sg13g2_buf_1 place7404 (.A(_07114_),
    .X(net7403));
 sg13g2_buf_1 place7405 (.A(net7405),
    .X(net7404));
 sg13g2_buf_1 place7406 (.A(_07109_),
    .X(net7405));
 sg13g2_buf_1 place7407 (.A(net7407),
    .X(net7406));
 sg13g2_buf_1 place7408 (.A(_07108_),
    .X(net7407));
 sg13g2_buf_1 place7409 (.A(_07108_),
    .X(net7408));
 sg13g2_buf_1 place7410 (.A(_07103_),
    .X(net7409));
 sg13g2_buf_1 place7411 (.A(_07102_),
    .X(net7410));
 sg13g2_buf_1 place7412 (.A(net7412),
    .X(net7411));
 sg13g2_buf_1 place7413 (.A(_07102_),
    .X(net7412));
 sg13g2_buf_1 place7414 (.A(_07102_),
    .X(net7413));
 sg13g2_buf_1 place7415 (.A(_06968_),
    .X(net7414));
 sg13g2_buf_1 place7416 (.A(net7416),
    .X(net7415));
 sg13g2_buf_1 place7417 (.A(net7417),
    .X(net7416));
 sg13g2_buf_1 place7418 (.A(_06968_),
    .X(net7417));
 sg13g2_buf_1 place7419 (.A(_02604_),
    .X(net7418));
 sg13g2_buf_1 place7420 (.A(net7420),
    .X(net7419));
 sg13g2_buf_1 place7421 (.A(_13579_),
    .X(net7420));
 sg13g2_buf_2 place7422 (.A(_12139_),
    .X(net7421));
 sg13g2_buf_1 place7423 (.A(_10463_),
    .X(net7422));
 sg13g2_buf_1 place7424 (.A(_10463_),
    .X(net7423));
 sg13g2_buf_2 place7425 (.A(_10449_),
    .X(net7424));
 sg13g2_buf_1 place7426 (.A(net7426),
    .X(net7425));
 sg13g2_buf_1 place7427 (.A(net7427),
    .X(net7426));
 sg13g2_buf_1 place7428 (.A(net7429),
    .X(net7427));
 sg13g2_buf_1 place7429 (.A(net7429),
    .X(net7428));
 sg13g2_buf_1 place7430 (.A(_09263_),
    .X(net7429));
 sg13g2_buf_1 place7431 (.A(_08850_),
    .X(net7430));
 sg13g2_buf_1 place7432 (.A(_08725_),
    .X(net7431));
 sg13g2_buf_1 place7433 (.A(_08634_),
    .X(net7432));
 sg13g2_buf_2 place7434 (.A(net7434),
    .X(net7433));
 sg13g2_buf_4 place7435 (.X(net7434),
    .A(_08387_));
 sg13g2_buf_1 place7436 (.A(_08288_),
    .X(net7435));
 sg13g2_buf_1 place7437 (.A(_08288_),
    .X(net7436));
 sg13g2_buf_1 place7438 (.A(_07672_),
    .X(net7437));
 sg13g2_buf_1 place7439 (.A(_07602_),
    .X(net7438));
 sg13g2_buf_1 place7440 (.A(_07201_),
    .X(net7439));
 sg13g2_buf_1 place7441 (.A(_03827_),
    .X(net7440));
 sg13g2_buf_1 place7442 (.A(_03827_),
    .X(net7441));
 sg13g2_buf_1 place7443 (.A(_14476_),
    .X(net7442));
 sg13g2_buf_1 place7444 (.A(_12187_),
    .X(net7443));
 sg13g2_buf_1 place7445 (.A(net7445),
    .X(net7444));
 sg13g2_buf_2 place7446 (.A(_12187_),
    .X(net7445));
 sg13g2_buf_1 place7447 (.A(_11477_),
    .X(net7446));
 sg13g2_buf_1 place7448 (.A(_11158_),
    .X(net7447));
 sg13g2_buf_1 place7449 (.A(_10982_),
    .X(net7448));
 sg13g2_buf_1 place7450 (.A(_10982_),
    .X(net7449));
 sg13g2_buf_1 place7451 (.A(_10980_),
    .X(net7450));
 sg13g2_buf_1 place7452 (.A(net7455),
    .X(net7451));
 sg13g2_buf_1 place7453 (.A(net7453),
    .X(net7452));
 sg13g2_buf_1 place7454 (.A(net7454),
    .X(net7453));
 sg13g2_buf_1 place7455 (.A(net7455),
    .X(net7454));
 sg13g2_buf_1 place7456 (.A(_10215_),
    .X(net7455));
 sg13g2_buf_1 place7457 (.A(_10191_),
    .X(net7456));
 sg13g2_buf_1 place7458 (.A(net7458),
    .X(net7457));
 sg13g2_buf_1 place7459 (.A(net7460),
    .X(net7458));
 sg13g2_buf_1 place7460 (.A(net7460),
    .X(net7459));
 sg13g2_buf_1 place7461 (.A(_10191_),
    .X(net7460));
 sg13g2_buf_1 place7462 (.A(_10191_),
    .X(net7461));
 sg13g2_buf_1 place7463 (.A(_10189_),
    .X(net7462));
 sg13g2_buf_1 place7464 (.A(_10189_),
    .X(net7463));
 sg13g2_buf_1 place7465 (.A(_10189_),
    .X(net7464));
 sg13g2_buf_1 place7466 (.A(net7466),
    .X(net7465));
 sg13g2_buf_1 place7467 (.A(net7470),
    .X(net7466));
 sg13g2_buf_1 place7468 (.A(net7470),
    .X(net7467));
 sg13g2_buf_1 place7469 (.A(net7469),
    .X(net7468));
 sg13g2_buf_1 place7470 (.A(net7470),
    .X(net7469));
 sg13g2_buf_1 place7471 (.A(_10182_),
    .X(net7470));
 sg13g2_buf_1 place7472 (.A(_10179_),
    .X(net7471));
 sg13g2_buf_1 place7473 (.A(_10179_),
    .X(net7472));
 sg13g2_buf_1 place7474 (.A(_10179_),
    .X(net7473));
 sg13g2_buf_1 place7475 (.A(_09679_),
    .X(net7474));
 sg13g2_buf_1 place7476 (.A(net7476),
    .X(net7475));
 sg13g2_buf_1 place7477 (.A(_09366_),
    .X(net7476));
 sg13g2_buf_1 place7478 (.A(_09282_),
    .X(net7477));
 sg13g2_buf_1 place7479 (.A(net7481),
    .X(net7478));
 sg13g2_buf_1 place7480 (.A(net7480),
    .X(net7479));
 sg13g2_buf_1 place7481 (.A(net7481),
    .X(net7480));
 sg13g2_buf_1 place7482 (.A(_09260_),
    .X(net7481));
 sg13g2_buf_1 place7483 (.A(_09244_),
    .X(net7482));
 sg13g2_buf_1 place7484 (.A(_09153_),
    .X(net7483));
 sg13g2_buf_1 place7485 (.A(net7485),
    .X(net7484));
 sg13g2_buf_1 place7486 (.A(_09153_),
    .X(net7485));
 sg13g2_buf_1 place7487 (.A(_09153_),
    .X(net7486));
 sg13g2_buf_1 place7488 (.A(net7489),
    .X(net7487));
 sg13g2_buf_1 place7489 (.A(net7489),
    .X(net7488));
 sg13g2_buf_1 place7490 (.A(_09152_),
    .X(net7489));
 sg13g2_buf_1 place7491 (.A(_09152_),
    .X(net7490));
 sg13g2_buf_1 place7492 (.A(net7492),
    .X(net7491));
 sg13g2_buf_1 place7493 (.A(_09152_),
    .X(net7492));
 sg13g2_buf_1 place7494 (.A(net7495),
    .X(net7493));
 sg13g2_buf_1 place7495 (.A(net7495),
    .X(net7494));
 sg13g2_buf_1 place7496 (.A(net7496),
    .X(net7495));
 sg13g2_buf_1 place7497 (.A(_09150_),
    .X(net7496));
 sg13g2_buf_1 place7498 (.A(_09150_),
    .X(net7497));
 sg13g2_buf_1 place7499 (.A(_09150_),
    .X(net7498));
 sg13g2_buf_1 place7500 (.A(_09073_),
    .X(net7499));
 sg13g2_buf_1 place7501 (.A(_09073_),
    .X(net7500));
 sg13g2_buf_1 place7502 (.A(net7503),
    .X(net7501));
 sg13g2_buf_1 place7503 (.A(net7503),
    .X(net7502));
 sg13g2_buf_1 place7504 (.A(_09070_),
    .X(net7503));
 sg13g2_buf_1 place7505 (.A(_09028_),
    .X(net7504));
 sg13g2_buf_1 place7506 (.A(net7508),
    .X(net7505));
 sg13g2_buf_1 place7507 (.A(net7508),
    .X(net7506));
 sg13g2_buf_1 place7508 (.A(net7508),
    .X(net7507));
 sg13g2_buf_1 place7509 (.A(_09028_),
    .X(net7508));
 sg13g2_buf_1 place7510 (.A(net7510),
    .X(net7509));
 sg13g2_buf_1 place7511 (.A(_09028_),
    .X(net7510));
 sg13g2_buf_1 place7512 (.A(_09026_),
    .X(net7511));
 sg13g2_buf_1 place7513 (.A(_09026_),
    .X(net7512));
 sg13g2_buf_1 place7514 (.A(net7515),
    .X(net7513));
 sg13g2_buf_2 place7515 (.A(net7515),
    .X(net7514));
 sg13g2_buf_1 place7516 (.A(_09026_),
    .X(net7515));
 sg13g2_buf_1 place7517 (.A(net7517),
    .X(net7516));
 sg13g2_buf_1 place7518 (.A(_09011_),
    .X(net7517));
 sg13g2_buf_1 place7519 (.A(net7519),
    .X(net7518));
 sg13g2_buf_2 place7520 (.A(_09011_),
    .X(net7519));
 sg13g2_buf_1 place7521 (.A(net7521),
    .X(net7520));
 sg13g2_buf_1 place7522 (.A(_09004_),
    .X(net7521));
 sg13g2_buf_1 place7523 (.A(net7523),
    .X(net7522));
 sg13g2_buf_1 place7524 (.A(_09004_),
    .X(net7523));
 sg13g2_buf_1 place7525 (.A(_09004_),
    .X(net7524));
 sg13g2_buf_1 place7526 (.A(_09001_),
    .X(net7525));
 sg13g2_buf_1 place7527 (.A(_09001_),
    .X(net7526));
 sg13g2_buf_1 place7528 (.A(_08988_),
    .X(net7527));
 sg13g2_buf_1 place7529 (.A(_08974_),
    .X(net7528));
 sg13g2_buf_1 place7530 (.A(_08974_),
    .X(net7529));
 sg13g2_buf_1 place7531 (.A(_08973_),
    .X(net7530));
 sg13g2_buf_1 place7532 (.A(_08946_),
    .X(net7531));
 sg13g2_buf_1 place7533 (.A(_08946_),
    .X(net7532));
 sg13g2_buf_1 place7534 (.A(net7534),
    .X(net7533));
 sg13g2_buf_1 place7535 (.A(_08946_),
    .X(net7534));
 sg13g2_buf_1 place7536 (.A(net7540),
    .X(net7535));
 sg13g2_buf_1 place7537 (.A(net7540),
    .X(net7536));
 sg13g2_buf_1 place7538 (.A(net7539),
    .X(net7537));
 sg13g2_buf_1 place7539 (.A(net7539),
    .X(net7538));
 sg13g2_buf_1 place7540 (.A(net7540),
    .X(net7539));
 sg13g2_buf_1 place7541 (.A(_08892_),
    .X(net7540));
 sg13g2_buf_1 place7542 (.A(net7542),
    .X(net7541));
 sg13g2_buf_1 place7543 (.A(_08889_),
    .X(net7542));
 sg13g2_buf_1 place7544 (.A(net7544),
    .X(net7543));
 sg13g2_buf_1 place7545 (.A(net7545),
    .X(net7544));
 sg13g2_buf_1 place7546 (.A(net7546),
    .X(net7545));
 sg13g2_buf_1 place7547 (.A(_08889_),
    .X(net7546));
 sg13g2_buf_1 place7548 (.A(net7549),
    .X(net7547));
 sg13g2_buf_1 place7549 (.A(net7549),
    .X(net7548));
 sg13g2_buf_1 place7550 (.A(_08889_),
    .X(net7549));
 sg13g2_buf_1 place7551 (.A(_08527_),
    .X(net7550));
 sg13g2_buf_1 place7552 (.A(net7553),
    .X(net7551));
 sg13g2_buf_1 place7553 (.A(net7553),
    .X(net7552));
 sg13g2_buf_2 place7554 (.A(net7554),
    .X(net7553));
 sg13g2_buf_2 place7555 (.A(_08527_),
    .X(net7554));
 sg13g2_buf_1 place7556 (.A(net7556),
    .X(net7555));
 sg13g2_buf_2 place7557 (.A(_08527_),
    .X(net7556));
 sg13g2_buf_1 place7558 (.A(net7558),
    .X(net7557));
 sg13g2_buf_4 place7559 (.X(net7558),
    .A(_08503_));
 sg13g2_buf_1 place7560 (.A(_08503_),
    .X(net7559));
 sg13g2_buf_4 place7561 (.X(net7560),
    .A(_08503_));
 sg13g2_buf_1 place7562 (.A(_08485_),
    .X(net7561));
 sg13g2_buf_1 place7563 (.A(_08485_),
    .X(net7562));
 sg13g2_buf_1 place7564 (.A(_08485_),
    .X(net7563));
 sg13g2_buf_1 place7565 (.A(_08485_),
    .X(net7564));
 sg13g2_buf_1 place7566 (.A(_08485_),
    .X(net7565));
 sg13g2_buf_1 place7567 (.A(_08485_),
    .X(net7566));
 sg13g2_buf_1 place7568 (.A(net7569),
    .X(net7567));
 sg13g2_buf_1 place7569 (.A(net7569),
    .X(net7568));
 sg13g2_buf_1 place7570 (.A(_08464_),
    .X(net7569));
 sg13g2_buf_1 place7571 (.A(_08464_),
    .X(net7570));
 sg13g2_buf_1 place7572 (.A(_08464_),
    .X(net7571));
 sg13g2_buf_1 place7573 (.A(net7574),
    .X(net7572));
 sg13g2_buf_1 place7574 (.A(net7574),
    .X(net7573));
 sg13g2_buf_1 place7575 (.A(_08462_),
    .X(net7574));
 sg13g2_buf_1 place7576 (.A(_08462_),
    .X(net7575));
 sg13g2_buf_1 place7577 (.A(_08462_),
    .X(net7576));
 sg13g2_buf_1 place7578 (.A(net7578),
    .X(net7577));
 sg13g2_buf_1 place7579 (.A(net7585),
    .X(net7578));
 sg13g2_buf_1 place7580 (.A(net7582),
    .X(net7579));
 sg13g2_buf_1 place7581 (.A(net7582),
    .X(net7580));
 sg13g2_buf_1 place7582 (.A(net7582),
    .X(net7581));
 sg13g2_buf_1 place7583 (.A(net7585),
    .X(net7582));
 sg13g2_buf_1 place7584 (.A(net7584),
    .X(net7583));
 sg13g2_buf_1 place7585 (.A(net7585),
    .X(net7584));
 sg13g2_buf_2 place7586 (.A(_08462_),
    .X(net7585));
 sg13g2_buf_1 place7587 (.A(net7587),
    .X(net7586));
 sg13g2_buf_1 place7588 (.A(_08424_),
    .X(net7587));
 sg13g2_buf_1 place7589 (.A(_08424_),
    .X(net7588));
 sg13g2_buf_1 place7590 (.A(net7590),
    .X(net7589));
 sg13g2_buf_1 place7591 (.A(_08384_),
    .X(net7590));
 sg13g2_buf_1 place7592 (.A(net7592),
    .X(net7591));
 sg13g2_buf_1 place7593 (.A(_08384_),
    .X(net7592));
 sg13g2_buf_1 place7594 (.A(_08313_),
    .X(net7593));
 sg13g2_buf_1 place7595 (.A(_08313_),
    .X(net7594));
 sg13g2_buf_1 place7596 (.A(net7596),
    .X(net7595));
 sg13g2_buf_2 place7597 (.A(_08313_),
    .X(net7596));
 sg13g2_buf_1 place7598 (.A(_08307_),
    .X(net7597));
 sg13g2_buf_2 place7599 (.A(_08306_),
    .X(net7598));
 sg13g2_buf_1 place7600 (.A(_08305_),
    .X(net7599));
 sg13g2_buf_1 place7601 (.A(_08291_),
    .X(net7600));
 sg13g2_buf_1 place7602 (.A(_08291_),
    .X(net7601));
 sg13g2_buf_1 place7603 (.A(_08255_),
    .X(net7602));
 sg13g2_buf_1 place7604 (.A(net7604),
    .X(net7603));
 sg13g2_buf_1 place7605 (.A(_08255_),
    .X(net7604));
 sg13g2_buf_1 place7606 (.A(_08255_),
    .X(net7605));
 sg13g2_buf_1 place7607 (.A(_08255_),
    .X(net7606));
 sg13g2_buf_1 place7608 (.A(_07790_),
    .X(net7607));
 sg13g2_buf_1 place7609 (.A(_07593_),
    .X(net7608));
 sg13g2_buf_1 place7610 (.A(_07567_),
    .X(net7609));
 sg13g2_buf_1 place7611 (.A(_07559_),
    .X(net7610));
 sg13g2_buf_1 place7612 (.A(_07202_),
    .X(net7611));
 sg13g2_buf_1 place7613 (.A(_07200_),
    .X(net7612));
 sg13g2_buf_1 place7614 (.A(_07188_),
    .X(net7613));
 sg13g2_buf_1 place7615 (.A(net7615),
    .X(net7614));
 sg13g2_buf_1 place7616 (.A(_07168_),
    .X(net7615));
 sg13g2_buf_1 place7617 (.A(_07154_),
    .X(net7616));
 sg13g2_buf_1 place7618 (.A(_07144_),
    .X(net7617));
 sg13g2_buf_1 place7619 (.A(_07141_),
    .X(net7618));
 sg13g2_buf_1 place7620 (.A(_07140_),
    .X(net7619));
 sg13g2_buf_1 place7621 (.A(_07132_),
    .X(net7620));
 sg13g2_buf_1 place7622 (.A(_07123_),
    .X(net7621));
 sg13g2_buf_1 place7623 (.A(net7624),
    .X(net7622));
 sg13g2_buf_1 place7624 (.A(net7624),
    .X(net7623));
 sg13g2_buf_1 place7625 (.A(net7625),
    .X(net7624));
 sg13g2_buf_1 place7626 (.A(_06902_),
    .X(net7625));
 sg13g2_buf_1 place7627 (.A(_06896_),
    .X(net7626));
 sg13g2_buf_1 place7628 (.A(_06619_),
    .X(net7627));
 sg13g2_buf_1 place7629 (.A(_06077_),
    .X(net7628));
 sg13g2_buf_1 place7630 (.A(_05186_),
    .X(net7629));
 sg13g2_buf_1 place7631 (.A(net7631),
    .X(net7630));
 sg13g2_buf_1 place7632 (.A(_05180_),
    .X(net7631));
 sg13g2_buf_1 place7633 (.A(net7633),
    .X(net7632));
 sg13g2_buf_1 place7634 (.A(net7634),
    .X(net7633));
 sg13g2_buf_1 place7635 (.A(_03823_),
    .X(net7634));
 sg13g2_buf_1 place7636 (.A(net7636),
    .X(net7635));
 sg13g2_buf_1 place7637 (.A(_03822_),
    .X(net7636));
 sg13g2_buf_1 place7638 (.A(net7638),
    .X(net7637));
 sg13g2_buf_1 place7639 (.A(_03815_),
    .X(net7638));
 sg13g2_buf_1 place7640 (.A(_03815_),
    .X(net7639));
 sg13g2_buf_1 place7641 (.A(_02462_),
    .X(net7640));
 sg13g2_buf_1 place7642 (.A(net7642),
    .X(net7641));
 sg13g2_buf_1 place7643 (.A(_01987_),
    .X(net7642));
 sg13g2_buf_1 place7644 (.A(net7644),
    .X(net7643));
 sg13g2_buf_1 place7645 (.A(net7648),
    .X(net7644));
 sg13g2_buf_1 place7646 (.A(net7646),
    .X(net7645));
 sg13g2_buf_1 place7647 (.A(net7647),
    .X(net7646));
 sg13g2_buf_1 place7648 (.A(net7648),
    .X(net7647));
 sg13g2_buf_1 place7649 (.A(_01987_),
    .X(net7648));
 sg13g2_buf_1 place7650 (.A(net7650),
    .X(net7649));
 sg13g2_buf_1 place7651 (.A(_01986_),
    .X(net7650));
 sg13g2_buf_1 place7652 (.A(net7656),
    .X(net7651));
 sg13g2_buf_1 place7653 (.A(net7654),
    .X(net7652));
 sg13g2_buf_1 place7654 (.A(net7654),
    .X(net7653));
 sg13g2_buf_1 place7655 (.A(net7655),
    .X(net7654));
 sg13g2_buf_1 place7656 (.A(net7656),
    .X(net7655));
 sg13g2_buf_1 place7657 (.A(_01986_),
    .X(net7656));
 sg13g2_buf_1 place7658 (.A(_01985_),
    .X(net7657));
 sg13g2_buf_1 place7659 (.A(net7659),
    .X(net7658));
 sg13g2_buf_1 place7660 (.A(_01984_),
    .X(net7659));
 sg13g2_buf_1 place7661 (.A(_01983_),
    .X(net7660));
 sg13g2_buf_1 place7662 (.A(_01982_),
    .X(net7661));
 sg13g2_buf_1 place7663 (.A(net7663),
    .X(net7662));
 sg13g2_buf_1 place7664 (.A(net7664),
    .X(net7663));
 sg13g2_buf_1 place7665 (.A(_00007_),
    .X(net7664));
 sg13g2_buf_1 place7666 (.A(\id_stage_i.controller_i.instr_valid_i ),
    .X(net7665));
 sg13g2_buf_1 place7667 (.A(_01917_),
    .X(net7666));
 sg13g2_buf_1 place7668 (.A(net7668),
    .X(net7667));
 sg13g2_buf_1 place7669 (.A(net7671),
    .X(net7668));
 sg13g2_buf_1 place7670 (.A(net7670),
    .X(net7669));
 sg13g2_buf_1 place7671 (.A(net7671),
    .X(net7670));
 sg13g2_buf_1 place7672 (.A(_01916_),
    .X(net7671));
 sg13g2_buf_1 place7673 (.A(_01914_),
    .X(net7672));
 sg13g2_buf_1 place7674 (.A(_01913_),
    .X(net7673));
 sg13g2_buf_1 place7675 (.A(_01913_),
    .X(net7674));
 sg13g2_buf_1 place7676 (.A(_01912_),
    .X(net7675));
 sg13g2_buf_1 place7677 (.A(_01911_),
    .X(net7676));
 sg13g2_buf_1 place7678 (.A(_01910_),
    .X(net7677));
 sg13g2_buf_1 place7679 (.A(_01909_),
    .X(net7678));
 sg13g2_buf_1 place7680 (.A(_01908_),
    .X(net7679));
 sg13g2_buf_1 place7681 (.A(_01907_),
    .X(net7680));
 sg13g2_buf_1 place7682 (.A(_01906_),
    .X(net7681));
 sg13g2_buf_1 place7683 (.A(_01905_),
    .X(net7682));
 sg13g2_buf_1 place7684 (.A(_01904_),
    .X(net7683));
 sg13g2_buf_1 place7685 (.A(_01903_),
    .X(net7684));
 sg13g2_buf_1 place7686 (.A(net7688),
    .X(net7685));
 sg13g2_buf_1 place7687 (.A(net7687),
    .X(net7686));
 sg13g2_buf_1 place7688 (.A(net7688),
    .X(net7687));
 sg13g2_buf_1 place7689 (.A(net7689),
    .X(net7688));
 sg13g2_buf_1 place7690 (.A(_01902_),
    .X(net7689));
 sg13g2_buf_1 place7691 (.A(net7691),
    .X(net7690));
 sg13g2_buf_1 place7692 (.A(_01902_),
    .X(net7691));
 sg13g2_buf_1 place7693 (.A(net7693),
    .X(net7692));
 sg13g2_buf_1 place7694 (.A(_01901_),
    .X(net7693));
 sg13g2_buf_1 place7695 (.A(net7695),
    .X(net7694));
 sg13g2_buf_1 place7696 (.A(net7696),
    .X(net7695));
 sg13g2_buf_1 place7697 (.A(_01901_),
    .X(net7696));
 sg13g2_buf_1 place7698 (.A(_01901_),
    .X(net7697));
 sg13g2_buf_1 place7699 (.A(net7702),
    .X(net7698));
 sg13g2_buf_1 place7700 (.A(net7700),
    .X(net7699));
 sg13g2_buf_1 place7701 (.A(net7701),
    .X(net7700));
 sg13g2_buf_1 place7702 (.A(net7702),
    .X(net7701));
 sg13g2_buf_1 place7703 (.A(_01900_),
    .X(net7702));
 sg13g2_buf_1 place7704 (.A(net7705),
    .X(net7703));
 sg13g2_buf_1 place7705 (.A(net7705),
    .X(net7704));
 sg13g2_buf_1 place7706 (.A(net7706),
    .X(net7705));
 sg13g2_buf_1 place7707 (.A(_01900_),
    .X(net7706));
 sg13g2_buf_1 place7708 (.A(net7708),
    .X(net7707));
 sg13g2_buf_1 place7709 (.A(net7710),
    .X(net7708));
 sg13g2_buf_1 place7710 (.A(net7710),
    .X(net7709));
 sg13g2_buf_1 place7711 (.A(net7711),
    .X(net7710));
 sg13g2_buf_1 place7712 (.A(net7712),
    .X(net7711));
 sg13g2_buf_1 place7713 (.A(net7715),
    .X(net7712));
 sg13g2_buf_1 place7714 (.A(net7714),
    .X(net7713));
 sg13g2_buf_1 place7715 (.A(net7715),
    .X(net7714));
 sg13g2_buf_1 place7716 (.A(_01900_),
    .X(net7715));
 sg13g2_buf_1 place7717 (.A(net7717),
    .X(net7716));
 sg13g2_buf_1 place7718 (.A(_01900_),
    .X(net7717));
 sg13g2_buf_1 place7719 (.A(net7721),
    .X(net7718));
 sg13g2_buf_1 place7720 (.A(net7720),
    .X(net7719));
 sg13g2_buf_1 place7721 (.A(net7721),
    .X(net7720));
 sg13g2_buf_1 place7722 (.A(net7732),
    .X(net7721));
 sg13g2_buf_1 place7723 (.A(net7730),
    .X(net7722));
 sg13g2_buf_1 place7724 (.A(net7725),
    .X(net7723));
 sg13g2_buf_1 place7725 (.A(net7725),
    .X(net7724));
 sg13g2_buf_1 place7726 (.A(net7730),
    .X(net7725));
 sg13g2_buf_1 place7727 (.A(net7728),
    .X(net7726));
 sg13g2_buf_1 place7728 (.A(net7728),
    .X(net7727));
 sg13g2_buf_1 place7729 (.A(net7729),
    .X(net7728));
 sg13g2_buf_2 place7730 (.A(net7730),
    .X(net7729));
 sg13g2_buf_2 place7731 (.A(net7732),
    .X(net7730));
 sg13g2_buf_1 place7732 (.A(net7732),
    .X(net7731));
 sg13g2_buf_1 place7733 (.A(_01899_),
    .X(net7732));
 sg13g2_buf_1 place7734 (.A(net7735),
    .X(net7733));
 sg13g2_buf_1 place7735 (.A(net7735),
    .X(net7734));
 sg13g2_buf_1 place7736 (.A(_01899_),
    .X(net7735));
 sg13g2_buf_1 place7737 (.A(net7743),
    .X(net7736));
 sg13g2_buf_1 place7738 (.A(net7739),
    .X(net7737));
 sg13g2_buf_1 place7739 (.A(net7739),
    .X(net7738));
 sg13g2_buf_1 place7740 (.A(net7743),
    .X(net7739));
 sg13g2_buf_1 place7741 (.A(net7742),
    .X(net7740));
 sg13g2_buf_1 place7742 (.A(net7742),
    .X(net7741));
 sg13g2_buf_1 place7743 (.A(net7743),
    .X(net7742));
 sg13g2_buf_1 place7744 (.A(_01899_),
    .X(net7743));
 sg13g2_buf_1 place7745 (.A(_01899_),
    .X(net7744));
 sg13g2_buf_1 place7746 (.A(net7747),
    .X(net7745));
 sg13g2_buf_1 place7747 (.A(net7747),
    .X(net7746));
 sg13g2_buf_1 place7748 (.A(_01899_),
    .X(net7747));
 sg13g2_buf_1 place7749 (.A(_01898_),
    .X(net7748));
 sg13g2_buf_1 place7750 (.A(net7753),
    .X(net7749));
 sg13g2_buf_1 place7751 (.A(net7752),
    .X(net7750));
 sg13g2_buf_1 place7752 (.A(net7752),
    .X(net7751));
 sg13g2_buf_1 place7753 (.A(net7753),
    .X(net7752));
 sg13g2_buf_2 place7754 (.A(net7762),
    .X(net7753));
 sg13g2_buf_1 place7755 (.A(net7757),
    .X(net7754));
 sg13g2_buf_1 place7756 (.A(net7757),
    .X(net7755));
 sg13g2_buf_1 place7757 (.A(net7757),
    .X(net7756));
 sg13g2_buf_1 place7758 (.A(net7759),
    .X(net7757));
 sg13g2_buf_1 place7759 (.A(net7759),
    .X(net7758));
 sg13g2_buf_1 place7760 (.A(net7762),
    .X(net7759));
 sg13g2_buf_1 place7761 (.A(net7761),
    .X(net7760));
 sg13g2_buf_1 place7762 (.A(net7762),
    .X(net7761));
 sg13g2_buf_1 place7763 (.A(_01898_),
    .X(net7762));
 sg13g2_buf_1 place7764 (.A(net7764),
    .X(net7763));
 sg13g2_buf_1 place7765 (.A(net7780),
    .X(net7764));
 sg13g2_buf_1 place7766 (.A(net7773),
    .X(net7765));
 sg13g2_buf_1 place7767 (.A(net7770),
    .X(net7766));
 sg13g2_buf_1 place7768 (.A(net7770),
    .X(net7767));
 sg13g2_buf_1 place7769 (.A(net7769),
    .X(net7768));
 sg13g2_buf_1 place7770 (.A(net7770),
    .X(net7769));
 sg13g2_buf_1 place7771 (.A(net7773),
    .X(net7770));
 sg13g2_buf_1 place7772 (.A(net7772),
    .X(net7771));
 sg13g2_buf_1 place7773 (.A(net7773),
    .X(net7772));
 sg13g2_buf_1 place7774 (.A(net7780),
    .X(net7773));
 sg13g2_buf_1 place7775 (.A(net7775),
    .X(net7774));
 sg13g2_buf_1 place7776 (.A(net7776),
    .X(net7775));
 sg13g2_buf_1 place7777 (.A(net7779),
    .X(net7776));
 sg13g2_buf_1 place7778 (.A(net7778),
    .X(net7777));
 sg13g2_buf_1 place7779 (.A(net7779),
    .X(net7778));
 sg13g2_buf_1 place7780 (.A(net7780),
    .X(net7779));
 sg13g2_buf_1 place7781 (.A(_01898_),
    .X(net7780));
 sg13g2_buf_1 place7782 (.A(net7788),
    .X(net7781));
 sg13g2_buf_1 place7783 (.A(net7788),
    .X(net7782));
 sg13g2_buf_1 place7784 (.A(net7785),
    .X(net7783));
 sg13g2_buf_1 place7785 (.A(net7785),
    .X(net7784));
 sg13g2_buf_1 place7786 (.A(net7787),
    .X(net7785));
 sg13g2_buf_1 place7787 (.A(net7787),
    .X(net7786));
 sg13g2_buf_2 place7788 (.A(net7788),
    .X(net7787));
 sg13g2_buf_2 place7789 (.A(net7804),
    .X(net7788));
 sg13g2_buf_1 place7790 (.A(net7804),
    .X(net7789));
 sg13g2_buf_1 place7791 (.A(net7804),
    .X(net7790));
 sg13g2_buf_1 place7792 (.A(net7792),
    .X(net7791));
 sg13g2_buf_1 place7793 (.A(net7804),
    .X(net7792));
 sg13g2_buf_1 place7794 (.A(net7794),
    .X(net7793));
 sg13g2_buf_1 place7795 (.A(net7795),
    .X(net7794));
 sg13g2_buf_1 place7796 (.A(net7796),
    .X(net7795));
 sg13g2_buf_1 place7797 (.A(net7797),
    .X(net7796));
 sg13g2_buf_1 place7798 (.A(net7804),
    .X(net7797));
 sg13g2_buf_1 place7799 (.A(net7803),
    .X(net7798));
 sg13g2_buf_1 place7800 (.A(net7800),
    .X(net7799));
 sg13g2_buf_1 place7801 (.A(net7802),
    .X(net7800));
 sg13g2_buf_1 place7802 (.A(net7802),
    .X(net7801));
 sg13g2_buf_1 place7803 (.A(net7803),
    .X(net7802));
 sg13g2_buf_1 place7804 (.A(net7804),
    .X(net7803));
 sg13g2_buf_2 place7805 (.A(_01898_),
    .X(net7804));
 sg13g2_buf_1 place7806 (.A(_01896_),
    .X(net7805));
 sg13g2_buf_1 place7807 (.A(_01896_),
    .X(net7806));
 sg13g2_buf_1 place7808 (.A(_01895_),
    .X(net7807));
 sg13g2_buf_1 place7809 (.A(_01895_),
    .X(net7808));
 sg13g2_buf_1 place7810 (.A(_01894_),
    .X(net7809));
 sg13g2_buf_1 place7811 (.A(net7813),
    .X(net7810));
 sg13g2_buf_1 place7812 (.A(net7812),
    .X(net7811));
 sg13g2_buf_1 place7813 (.A(net7813),
    .X(net7812));
 sg13g2_buf_1 place7814 (.A(_01894_),
    .X(net7813));
 sg13g2_buf_1 place7815 (.A(net7816),
    .X(net7814));
 sg13g2_buf_1 place7816 (.A(net7816),
    .X(net7815));
 sg13g2_buf_2 place7817 (.A(_01894_),
    .X(net7816));
 sg13g2_buf_1 place7818 (.A(net7818),
    .X(net7817));
 sg13g2_buf_1 place7819 (.A(net7819),
    .X(net7818));
 sg13g2_buf_1 place7820 (.A(net7831),
    .X(net7819));
 sg13g2_buf_1 place7821 (.A(net7821),
    .X(net7820));
 sg13g2_buf_1 place7822 (.A(net7823),
    .X(net7821));
 sg13g2_buf_1 place7823 (.A(net7823),
    .X(net7822));
 sg13g2_buf_1 place7824 (.A(net7827),
    .X(net7823));
 sg13g2_buf_1 place7825 (.A(net7825),
    .X(net7824));
 sg13g2_buf_1 place7826 (.A(net7826),
    .X(net7825));
 sg13g2_buf_1 place7827 (.A(net7827),
    .X(net7826));
 sg13g2_buf_1 place7828 (.A(net7831),
    .X(net7827));
 sg13g2_buf_1 place7829 (.A(net7829),
    .X(net7828));
 sg13g2_buf_1 place7830 (.A(net7831),
    .X(net7829));
 sg13g2_buf_1 place7831 (.A(net7831),
    .X(net7830));
 sg13g2_buf_2 place7832 (.A(_01893_),
    .X(net7831));
 sg13g2_buf_1 place7833 (.A(_01893_),
    .X(net7832));
 sg13g2_buf_1 place7834 (.A(net7834),
    .X(net7833));
 sg13g2_buf_1 place7835 (.A(net7835),
    .X(net7834));
 sg13g2_buf_1 place7836 (.A(_01893_),
    .X(net7835));
 sg13g2_buf_1 place7837 (.A(net7837),
    .X(net7836));
 sg13g2_buf_1 place7838 (.A(net7838),
    .X(net7837));
 sg13g2_buf_1 place7839 (.A(net7862),
    .X(net7838));
 sg13g2_buf_1 place7840 (.A(net7841),
    .X(net7839));
 sg13g2_buf_1 place7841 (.A(net7841),
    .X(net7840));
 sg13g2_buf_1 place7842 (.A(net7842),
    .X(net7841));
 sg13g2_buf_1 place7843 (.A(net7862),
    .X(net7842));
 sg13g2_buf_1 place7844 (.A(net7862),
    .X(net7843));
 sg13g2_buf_1 place7845 (.A(net7855),
    .X(net7844));
 sg13g2_buf_1 place7846 (.A(net7855),
    .X(net7845));
 sg13g2_buf_1 place7847 (.A(net7847),
    .X(net7846));
 sg13g2_buf_1 place7848 (.A(net7850),
    .X(net7847));
 sg13g2_buf_1 place7849 (.A(net7849),
    .X(net7848));
 sg13g2_buf_1 place7850 (.A(net7850),
    .X(net7849));
 sg13g2_buf_1 place7851 (.A(net7852),
    .X(net7850));
 sg13g2_buf_1 place7852 (.A(net7852),
    .X(net7851));
 sg13g2_buf_1 place7853 (.A(net7855),
    .X(net7852));
 sg13g2_buf_1 place7854 (.A(net7854),
    .X(net7853));
 sg13g2_buf_1 place7855 (.A(net7855),
    .X(net7854));
 sg13g2_buf_2 place7856 (.A(net7862),
    .X(net7855));
 sg13g2_buf_1 place7857 (.A(net7862),
    .X(net7856));
 sg13g2_buf_1 place7858 (.A(net7861),
    .X(net7857));
 sg13g2_buf_1 place7859 (.A(net7860),
    .X(net7858));
 sg13g2_buf_1 place7860 (.A(net7860),
    .X(net7859));
 sg13g2_buf_1 place7861 (.A(net7861),
    .X(net7860));
 sg13g2_buf_1 place7862 (.A(net7862),
    .X(net7861));
 sg13g2_buf_1 place7863 (.A(_01892_),
    .X(net7862));
 sg13g2_buf_1 place7864 (.A(_01892_),
    .X(net7863));
 sg13g2_buf_1 place7865 (.A(net7865),
    .X(net7864));
 sg13g2_buf_1 place7866 (.A(_01892_),
    .X(net7865));
 sg13g2_buf_1 place7867 (.A(_01892_),
    .X(net7866));
 sg13g2_buf_1 place7868 (.A(net7880),
    .X(net7867));
 sg13g2_buf_1 place7869 (.A(net7875),
    .X(net7868));
 sg13g2_buf_1 place7870 (.A(net7870),
    .X(net7869));
 sg13g2_buf_1 place7871 (.A(net7871),
    .X(net7870));
 sg13g2_buf_1 place7872 (.A(net7875),
    .X(net7871));
 sg13g2_buf_1 place7873 (.A(net7875),
    .X(net7872));
 sg13g2_buf_1 place7874 (.A(net7875),
    .X(net7873));
 sg13g2_buf_1 place7875 (.A(net7875),
    .X(net7874));
 sg13g2_buf_1 place7876 (.A(net7880),
    .X(net7875));
 sg13g2_buf_1 place7877 (.A(net7877),
    .X(net7876));
 sg13g2_buf_1 place7878 (.A(net7878),
    .X(net7877));
 sg13g2_buf_1 place7879 (.A(net7879),
    .X(net7878));
 sg13g2_buf_1 place7880 (.A(net7880),
    .X(net7879));
 sg13g2_buf_1 place7881 (.A(net7895),
    .X(net7880));
 sg13g2_buf_1 place7882 (.A(net7882),
    .X(net7881));
 sg13g2_buf_1 place7883 (.A(net7894),
    .X(net7882));
 sg13g2_buf_1 place7884 (.A(net7884),
    .X(net7883));
 sg13g2_buf_1 place7885 (.A(net7885),
    .X(net7884));
 sg13g2_buf_1 place7886 (.A(net7894),
    .X(net7885));
 sg13g2_buf_1 place7887 (.A(net7887),
    .X(net7886));
 sg13g2_buf_1 place7888 (.A(net7893),
    .X(net7887));
 sg13g2_buf_1 place7889 (.A(net7889),
    .X(net7888));
 sg13g2_buf_1 place7890 (.A(net7891),
    .X(net7889));
 sg13g2_buf_1 place7891 (.A(net7891),
    .X(net7890));
 sg13g2_buf_1 place7892 (.A(net7893),
    .X(net7891));
 sg13g2_buf_1 place7893 (.A(net7893),
    .X(net7892));
 sg13g2_buf_1 place7894 (.A(net7894),
    .X(net7893));
 sg13g2_buf_1 place7895 (.A(net7895),
    .X(net7894));
 sg13g2_buf_1 place7896 (.A(_01892_),
    .X(net7895));
 sg13g2_buf_1 place7897 (.A(net7897),
    .X(net7896));
 sg13g2_buf_1 place7898 (.A(net7900),
    .X(net7897));
 sg13g2_buf_1 place7899 (.A(net7900),
    .X(net7898));
 sg13g2_buf_2 place7900 (.A(net7900),
    .X(net7899));
 sg13g2_buf_2 place7901 (.A(net7919),
    .X(net7900));
 sg13g2_buf_1 place7902 (.A(net7906),
    .X(net7901));
 sg13g2_buf_1 place7903 (.A(net7906),
    .X(net7902));
 sg13g2_buf_1 place7904 (.A(net7904),
    .X(net7903));
 sg13g2_buf_1 place7905 (.A(net7906),
    .X(net7904));
 sg13g2_buf_1 place7906 (.A(net7906),
    .X(net7905));
 sg13g2_buf_1 place7907 (.A(net7919),
    .X(net7906));
 sg13g2_buf_1 place7908 (.A(net7912),
    .X(net7907));
 sg13g2_buf_1 place7909 (.A(net7909),
    .X(net7908));
 sg13g2_buf_1 place7910 (.A(net7912),
    .X(net7909));
 sg13g2_buf_1 place7911 (.A(net7911),
    .X(net7910));
 sg13g2_buf_1 place7912 (.A(net7912),
    .X(net7911));
 sg13g2_buf_1 place7913 (.A(net7919),
    .X(net7912));
 sg13g2_buf_1 place7914 (.A(net7914),
    .X(net7913));
 sg13g2_buf_1 place7915 (.A(net7919),
    .X(net7914));
 sg13g2_buf_1 place7916 (.A(net7916),
    .X(net7915));
 sg13g2_buf_1 place7917 (.A(net7919),
    .X(net7916));
 sg13g2_buf_1 place7918 (.A(net7918),
    .X(net7917));
 sg13g2_buf_2 place7919 (.A(net7919),
    .X(net7918));
 sg13g2_buf_1 place7920 (.A(_01892_),
    .X(net7919));
 sg13g2_buf_1 place7921 (.A(net7921),
    .X(net7920));
 sg13g2_buf_1 place7922 (.A(net7925),
    .X(net7921));
 sg13g2_buf_1 place7923 (.A(net7923),
    .X(net7922));
 sg13g2_buf_1 place7924 (.A(net7924),
    .X(net7923));
 sg13g2_buf_1 place7925 (.A(net7925),
    .X(net7924));
 sg13g2_buf_1 place7926 (.A(_01891_),
    .X(net7925));
 sg13g2_buf_1 place7927 (.A(net7928),
    .X(net7926));
 sg13g2_buf_1 place7928 (.A(net7928),
    .X(net7927));
 sg13g2_buf_1 place7929 (.A(_01890_),
    .X(net7928));
 sg13g2_buf_1 place7930 (.A(net7931),
    .X(net7929));
 sg13g2_buf_1 place7931 (.A(net7931),
    .X(net7930));
 sg13g2_buf_1 place7932 (.A(_01889_),
    .X(net7931));
 sg13g2_buf_1 place7933 (.A(_01887_),
    .X(net7932));
 sg13g2_buf_1 place7934 (.A(net7934),
    .X(net7933));
 sg13g2_buf_1 place7935 (.A(\id_stage_i.controller_i.instr_is_compressed_i ),
    .X(net7934));
 sg13g2_buf_1 place7936 (.A(net7936),
    .X(net7935));
 sg13g2_buf_1 place7937 (.A(\id_stage_i.controller_i.instr_is_compressed_i ),
    .X(net7936));
 sg13g2_buf_1 place7938 (.A(_01838_),
    .X(net7937));
 sg13g2_buf_1 place7939 (.A(_01837_),
    .X(net7938));
 sg13g2_buf_1 place7940 (.A(net7940),
    .X(net7939));
 sg13g2_buf_1 place7941 (.A(net7941),
    .X(net7940));
 sg13g2_buf_1 place7942 (.A(net7947),
    .X(net7941));
 sg13g2_buf_1 place7943 (.A(net7943),
    .X(net7942));
 sg13g2_buf_1 place7944 (.A(net7944),
    .X(net7943));
 sg13g2_buf_1 place7945 (.A(net7947),
    .X(net7944));
 sg13g2_buf_1 place7946 (.A(net7946),
    .X(net7945));
 sg13g2_buf_1 place7947 (.A(net7947),
    .X(net7946));
 sg13g2_buf_1 place7948 (.A(_01837_),
    .X(net7947));
 sg13g2_buf_1 place7949 (.A(net7949),
    .X(net7948));
 sg13g2_buf_1 place7950 (.A(net7956),
    .X(net7949));
 sg13g2_buf_1 place7951 (.A(net7955),
    .X(net7950));
 sg13g2_buf_1 place7952 (.A(net7955),
    .X(net7951));
 sg13g2_buf_1 place7953 (.A(net7953),
    .X(net7952));
 sg13g2_buf_1 place7954 (.A(net7954),
    .X(net7953));
 sg13g2_buf_1 place7955 (.A(net7955),
    .X(net7954));
 sg13g2_buf_1 place7956 (.A(net7956),
    .X(net7955));
 sg13g2_buf_1 place7957 (.A(_01836_),
    .X(net7956));
 sg13g2_buf_1 place7958 (.A(net7966),
    .X(net7957));
 sg13g2_buf_1 place7959 (.A(net7965),
    .X(net7958));
 sg13g2_buf_1 place7960 (.A(net7965),
    .X(net7959));
 sg13g2_buf_1 place7961 (.A(net7964),
    .X(net7960));
 sg13g2_buf_1 place7962 (.A(net7963),
    .X(net7961));
 sg13g2_buf_1 place7963 (.A(net7963),
    .X(net7962));
 sg13g2_buf_1 place7964 (.A(net7964),
    .X(net7963));
 sg13g2_buf_1 place7965 (.A(net7965),
    .X(net7964));
 sg13g2_buf_1 place7966 (.A(net7966),
    .X(net7965));
 sg13g2_buf_1 place7967 (.A(_01835_),
    .X(net7966));
 sg13g2_buf_1 place7968 (.A(net7968),
    .X(net7967));
 sg13g2_buf_1 place7969 (.A(net7976),
    .X(net7968));
 sg13g2_buf_1 place7970 (.A(net7970),
    .X(net7969));
 sg13g2_buf_1 place7971 (.A(net7974),
    .X(net7970));
 sg13g2_buf_1 place7972 (.A(net7972),
    .X(net7971));
 sg13g2_buf_1 place7973 (.A(net7973),
    .X(net7972));
 sg13g2_buf_1 place7974 (.A(net7974),
    .X(net7973));
 sg13g2_buf_1 place7975 (.A(net7975),
    .X(net7974));
 sg13g2_buf_1 place7976 (.A(net7976),
    .X(net7975));
 sg13g2_buf_1 place7977 (.A(_01718_),
    .X(net7976));
 sg13g2_buf_1 place7978 (.A(_01666_),
    .X(net7977));
 sg13g2_buf_1 place7979 (.A(_01657_),
    .X(net7978));
 sg13g2_buf_1 place7980 (.A(_01655_),
    .X(net7979));
 sg13g2_buf_1 place7981 (.A(_01654_),
    .X(net7980));
 sg13g2_buf_1 place7982 (.A(\id_stage_i.id_fsm_q ),
    .X(net7981));
 sg13g2_buf_1 place7983 (.A(net7983),
    .X(net7982));
 sg13g2_buf_1 place7984 (.A(\cs_registers_i.nmi_mode_i ),
    .X(net7983));
 sg13g2_buf_1 place7985 (.A(\cs_registers_i.debug_mode_i ),
    .X(net7984));
 sg13g2_buf_1 place7986 (.A(_01603_),
    .X(net7985));
 sg13g2_buf_1 place7987 (.A(_01603_),
    .X(net7986));
 sg13g2_buf_1 place7988 (.A(net7991),
    .X(net7987));
 sg13g2_buf_1 place7989 (.A(net7989),
    .X(net7988));
 sg13g2_buf_1 place7990 (.A(net7990),
    .X(net7989));
 sg13g2_buf_1 place7991 (.A(net7991),
    .X(net7990));
 sg13g2_buf_1 place7992 (.A(_00543_),
    .X(net7991));
 sg13g2_buf_1 place7993 (.A(net7994),
    .X(net7992));
 sg13g2_buf_1 place7994 (.A(net7994),
    .X(net7993));
 sg13g2_buf_1 place7995 (.A(net7995),
    .X(net7994));
 sg13g2_buf_1 place7996 (.A(net7996),
    .X(net7995));
 sg13g2_buf_1 place7997 (.A(net7997),
    .X(net7996));
 sg13g2_buf_1 place7998 (.A(net8002),
    .X(net7997));
 sg13g2_buf_1 place7999 (.A(net7999),
    .X(net7998));
 sg13g2_buf_1 place8000 (.A(net8001),
    .X(net7999));
 sg13g2_buf_1 place8001 (.A(net8001),
    .X(net8000));
 sg13g2_buf_1 place8002 (.A(net8002),
    .X(net8001));
 sg13g2_buf_1 place8003 (.A(_00542_),
    .X(net8002));
 sg13g2_buf_1 place8004 (.A(_00541_),
    .X(net8003));
 sg13g2_buf_1 place8005 (.A(net8005),
    .X(net8004));
 sg13g2_buf_1 place8006 (.A(net8008),
    .X(net8005));
 sg13g2_buf_1 place8007 (.A(net8007),
    .X(net8006));
 sg13g2_buf_1 place8008 (.A(net8008),
    .X(net8007));
 sg13g2_buf_1 place8009 (.A(_00541_),
    .X(net8008));
 sg13g2_buf_1 place8010 (.A(net8010),
    .X(net8009));
 sg13g2_buf_1 place8011 (.A(_00539_),
    .X(net8010));
 sg13g2_buf_1 place8012 (.A(net8013),
    .X(net8011));
 sg13g2_buf_1 place8013 (.A(net8013),
    .X(net8012));
 sg13g2_buf_1 place8014 (.A(net8014),
    .X(net8013));
 sg13g2_buf_1 place8015 (.A(net8015),
    .X(net8014));
 sg13g2_buf_1 place8016 (.A(_00005_),
    .X(net8015));
 sg13g2_buf_1 place8017 (.A(_00538_),
    .X(net8016));
 sg13g2_buf_1 place8018 (.A(_00535_),
    .X(net8017));
 sg13g2_buf_1 place8019 (.A(_00533_),
    .X(net8018));
 sg13g2_buf_1 place8020 (.A(net8020),
    .X(net8019));
 sg13g2_buf_1 place8021 (.A(_00532_),
    .X(net8020));
 sg13g2_buf_1 place8022 (.A(net8022),
    .X(net8021));
 sg13g2_buf_1 place8023 (.A(_00531_),
    .X(net8022));
 sg13g2_buf_1 place8024 (.A(net8082),
    .X(net8023));
 sg13g2_buf_1 place8025 (.A(net8027),
    .X(net8024));
 sg13g2_buf_1 place8026 (.A(net8026),
    .X(net8025));
 sg13g2_buf_1 place8027 (.A(net8027),
    .X(net8026));
 sg13g2_buf_1 place8028 (.A(net8082),
    .X(net8027));
 sg13g2_buf_1 place8029 (.A(net8033),
    .X(net8028));
 sg13g2_buf_1 place8030 (.A(net8033),
    .X(net8029));
 sg13g2_buf_1 place8031 (.A(net8031),
    .X(net8030));
 sg13g2_buf_1 place8032 (.A(net8032),
    .X(net8031));
 sg13g2_buf_1 place8033 (.A(net8033),
    .X(net8032));
 sg13g2_buf_1 place8034 (.A(net8082),
    .X(net8033));
 sg13g2_buf_1 place8035 (.A(net8081),
    .X(net8034));
 sg13g2_buf_1 place8036 (.A(net8040),
    .X(net8035));
 sg13g2_buf_1 place8037 (.A(net8040),
    .X(net8036));
 sg13g2_buf_1 place8038 (.A(net8039),
    .X(net8037));
 sg13g2_buf_1 place8039 (.A(net8039),
    .X(net8038));
 sg13g2_buf_1 place8040 (.A(net8040),
    .X(net8039));
 sg13g2_buf_1 place8041 (.A(net8081),
    .X(net8040));
 sg13g2_buf_1 place8042 (.A(net8050),
    .X(net8041));
 sg13g2_buf_1 place8043 (.A(net8043),
    .X(net8042));
 sg13g2_buf_1 place8044 (.A(net8050),
    .X(net8043));
 sg13g2_buf_1 place8045 (.A(net8048),
    .X(net8044));
 sg13g2_buf_1 place8046 (.A(net8047),
    .X(net8045));
 sg13g2_buf_1 place8047 (.A(net8047),
    .X(net8046));
 sg13g2_buf_1 place8048 (.A(net8048),
    .X(net8047));
 sg13g2_buf_1 place8049 (.A(net8049),
    .X(net8048));
 sg13g2_buf_1 place8050 (.A(net8050),
    .X(net8049));
 sg13g2_buf_1 place8051 (.A(net8081),
    .X(net8050));
 sg13g2_buf_1 place8052 (.A(net8079),
    .X(net8051));
 sg13g2_buf_1 place8053 (.A(net8053),
    .X(net8052));
 sg13g2_buf_1 place8054 (.A(net8064),
    .X(net8053));
 sg13g2_buf_1 place8055 (.A(net8055),
    .X(net8054));
 sg13g2_buf_1 place8056 (.A(net8064),
    .X(net8055));
 sg13g2_buf_1 place8057 (.A(net8057),
    .X(net8056));
 sg13g2_buf_1 place8058 (.A(net8063),
    .X(net8057));
 sg13g2_buf_1 place8059 (.A(net8059),
    .X(net8058));
 sg13g2_buf_1 place8060 (.A(net8062),
    .X(net8059));
 sg13g2_buf_1 place8061 (.A(net8061),
    .X(net8060));
 sg13g2_buf_1 place8062 (.A(net8062),
    .X(net8061));
 sg13g2_buf_1 place8063 (.A(net8063),
    .X(net8062));
 sg13g2_buf_1 place8064 (.A(net8064),
    .X(net8063));
 sg13g2_buf_1 place8065 (.A(net8079),
    .X(net8064));
 sg13g2_buf_1 place8066 (.A(net8066),
    .X(net8065));
 sg13g2_buf_1 place8067 (.A(net8067),
    .X(net8066));
 sg13g2_buf_1 place8068 (.A(net8078),
    .X(net8067));
 sg13g2_buf_1 place8069 (.A(net8069),
    .X(net8068));
 sg13g2_buf_1 place8070 (.A(net8078),
    .X(net8069));
 sg13g2_buf_1 place8071 (.A(net8078),
    .X(net8070));
 sg13g2_buf_1 place8072 (.A(net8072),
    .X(net8071));
 sg13g2_buf_1 place8073 (.A(net8076),
    .X(net8072));
 sg13g2_buf_1 place8074 (.A(net8075),
    .X(net8073));
 sg13g2_buf_1 place8075 (.A(net8075),
    .X(net8074));
 sg13g2_buf_1 place8076 (.A(net8076),
    .X(net8075));
 sg13g2_buf_1 place8077 (.A(net8078),
    .X(net8076));
 sg13g2_buf_1 place8078 (.A(net8078),
    .X(net8077));
 sg13g2_buf_1 place8079 (.A(net8079),
    .X(net8078));
 sg13g2_buf_1 place8080 (.A(net8080),
    .X(net8079));
 sg13g2_buf_1 place8081 (.A(net8081),
    .X(net8080));
 sg13g2_buf_1 place8082 (.A(net8082),
    .X(net8081));
 sg13g2_buf_1 place8083 (.A(net437),
    .X(net8082));
 sg13g2_buf_1 place8084 (.A(net8084),
    .X(net8083));
 sg13g2_buf_1 place8085 (.A(net8094),
    .X(net8084));
 sg13g2_buf_1 place8086 (.A(net8086),
    .X(net8085));
 sg13g2_buf_1 place8087 (.A(net8093),
    .X(net8086));
 sg13g2_buf_1 place8088 (.A(net8088),
    .X(net8087));
 sg13g2_buf_1 place8089 (.A(net8089),
    .X(net8088));
 sg13g2_buf_1 place8090 (.A(net8093),
    .X(net8089));
 sg13g2_buf_1 place8091 (.A(net8091),
    .X(net8090));
 sg13g2_buf_1 place8092 (.A(net8092),
    .X(net8091));
 sg13g2_buf_1 place8093 (.A(net8093),
    .X(net8092));
 sg13g2_buf_1 place8094 (.A(net8094),
    .X(net8093));
 sg13g2_buf_1 place8095 (.A(net8095),
    .X(net8094));
 sg13g2_buf_1 place8096 (.A(net8109),
    .X(net8095));
 sg13g2_buf_1 place8097 (.A(net8097),
    .X(net8096));
 sg13g2_buf_1 place8098 (.A(net8109),
    .X(net8097));
 sg13g2_buf_1 place8099 (.A(net8101),
    .X(net8098));
 sg13g2_buf_1 place8100 (.A(net8100),
    .X(net8099));
 sg13g2_buf_1 place8101 (.A(net8101),
    .X(net8100));
 sg13g2_buf_1 place8102 (.A(net8109),
    .X(net8101));
 sg13g2_buf_1 place8103 (.A(net8108),
    .X(net8102));
 sg13g2_buf_1 place8104 (.A(net8107),
    .X(net8103));
 sg13g2_buf_1 place8105 (.A(net8106),
    .X(net8104));
 sg13g2_buf_1 place8106 (.A(net8106),
    .X(net8105));
 sg13g2_buf_1 place8107 (.A(net8107),
    .X(net8106));
 sg13g2_buf_1 place8108 (.A(net8108),
    .X(net8107));
 sg13g2_buf_1 place8109 (.A(net8109),
    .X(net8108));
 sg13g2_buf_1 place8110 (.A(net437),
    .X(net8109));
 sg13g2_buf_1 place8111 (.A(net8124),
    .X(net8110));
 sg13g2_buf_1 place8112 (.A(net8118),
    .X(net8111));
 sg13g2_buf_1 place8113 (.A(net8113),
    .X(net8112));
 sg13g2_buf_1 place8114 (.A(net8118),
    .X(net8113));
 sg13g2_buf_1 place8115 (.A(net8118),
    .X(net8114));
 sg13g2_buf_1 place8116 (.A(net8116),
    .X(net8115));
 sg13g2_buf_1 place8117 (.A(net8117),
    .X(net8116));
 sg13g2_buf_1 place8118 (.A(net8118),
    .X(net8117));
 sg13g2_buf_1 place8119 (.A(net8124),
    .X(net8118));
 sg13g2_buf_1 place8120 (.A(net8120),
    .X(net8119));
 sg13g2_buf_1 place8121 (.A(net8123),
    .X(net8120));
 sg13g2_buf_1 place8122 (.A(net8123),
    .X(net8121));
 sg13g2_buf_1 place8123 (.A(net8123),
    .X(net8122));
 sg13g2_buf_1 place8124 (.A(net8124),
    .X(net8123));
 sg13g2_buf_1 place8125 (.A(net437),
    .X(net8124));
 sg13g2_buf_1 place8126 (.A(net8207),
    .X(net8125));
 sg13g2_buf_1 place8127 (.A(net8128),
    .X(net8126));
 sg13g2_buf_1 place8128 (.A(net8128),
    .X(net8127));
 sg13g2_buf_1 place8129 (.A(net8207),
    .X(net8128));
 sg13g2_buf_1 place8130 (.A(net8130),
    .X(net8129));
 sg13g2_buf_1 place8131 (.A(net8131),
    .X(net8130));
 sg13g2_buf_1 place8132 (.A(net8140),
    .X(net8131));
 sg13g2_buf_1 place8133 (.A(net8140),
    .X(net8132));
 sg13g2_buf_1 place8134 (.A(net8134),
    .X(net8133));
 sg13g2_buf_1 place8135 (.A(net8138),
    .X(net8134));
 sg13g2_buf_1 place8136 (.A(net8137),
    .X(net8135));
 sg13g2_buf_1 place8137 (.A(net8137),
    .X(net8136));
 sg13g2_buf_1 place8138 (.A(net8138),
    .X(net8137));
 sg13g2_buf_1 place8139 (.A(net8140),
    .X(net8138));
 sg13g2_buf_1 place8140 (.A(net8140),
    .X(net8139));
 sg13g2_buf_1 place8141 (.A(net8207),
    .X(net8140));
 sg13g2_buf_1 place8142 (.A(net8142),
    .X(net8141));
 sg13g2_buf_1 place8143 (.A(net8156),
    .X(net8142));
 sg13g2_buf_1 place8144 (.A(net8156),
    .X(net8143));
 sg13g2_buf_1 place8145 (.A(net8146),
    .X(net8144));
 sg13g2_buf_1 place8146 (.A(net8146),
    .X(net8145));
 sg13g2_buf_1 place8147 (.A(net8147),
    .X(net8146));
 sg13g2_buf_1 place8148 (.A(net8148),
    .X(net8147));
 sg13g2_buf_1 place8149 (.A(net8155),
    .X(net8148));
 sg13g2_buf_1 place8150 (.A(net8150),
    .X(net8149));
 sg13g2_buf_1 place8151 (.A(net8155),
    .X(net8150));
 sg13g2_buf_1 place8152 (.A(net8152),
    .X(net8151));
 sg13g2_buf_1 place8153 (.A(net8153),
    .X(net8152));
 sg13g2_buf_1 place8154 (.A(net8154),
    .X(net8153));
 sg13g2_buf_1 place8155 (.A(net8155),
    .X(net8154));
 sg13g2_buf_1 place8156 (.A(net8156),
    .X(net8155));
 sg13g2_buf_1 place8157 (.A(net8207),
    .X(net8156));
 sg13g2_buf_1 place8158 (.A(net8162),
    .X(net8157));
 sg13g2_buf_1 place8159 (.A(net8161),
    .X(net8158));
 sg13g2_buf_1 place8160 (.A(net8160),
    .X(net8159));
 sg13g2_buf_1 place8161 (.A(net8161),
    .X(net8160));
 sg13g2_buf_1 place8162 (.A(net8162),
    .X(net8161));
 sg13g2_buf_1 place8163 (.A(net8163),
    .X(net8162));
 sg13g2_buf_1 place8164 (.A(net8207),
    .X(net8163));
 sg13g2_buf_1 place8165 (.A(net8165),
    .X(net8164));
 sg13g2_buf_1 place8166 (.A(net8167),
    .X(net8165));
 sg13g2_buf_1 place8167 (.A(net8167),
    .X(net8166));
 sg13g2_buf_1 place8168 (.A(net8188),
    .X(net8167));
 sg13g2_buf_1 place8169 (.A(net8169),
    .X(net8168));
 sg13g2_buf_1 place8170 (.A(net8170),
    .X(net8169));
 sg13g2_buf_1 place8171 (.A(net8171),
    .X(net8170));
 sg13g2_buf_1 place8172 (.A(net8188),
    .X(net8171));
 sg13g2_buf_1 place8173 (.A(net8173),
    .X(net8172));
 sg13g2_buf_1 place8174 (.A(net8188),
    .X(net8173));
 sg13g2_buf_1 place8175 (.A(net8180),
    .X(net8174));
 sg13g2_buf_1 place8176 (.A(net8176),
    .X(net8175));
 sg13g2_buf_1 place8177 (.A(net8180),
    .X(net8176));
 sg13g2_buf_1 place8178 (.A(net8178),
    .X(net8177));
 sg13g2_buf_1 place8179 (.A(net8180),
    .X(net8178));
 sg13g2_buf_1 place8180 (.A(net8180),
    .X(net8179));
 sg13g2_buf_1 place8181 (.A(net8188),
    .X(net8180));
 sg13g2_buf_1 place8182 (.A(net8188),
    .X(net8181));
 sg13g2_buf_1 place8183 (.A(net8187),
    .X(net8182));
 sg13g2_buf_1 place8184 (.A(net8184),
    .X(net8183));
 sg13g2_buf_1 place8185 (.A(net8186),
    .X(net8184));
 sg13g2_buf_1 place8186 (.A(net8186),
    .X(net8185));
 sg13g2_buf_1 place8187 (.A(net8187),
    .X(net8186));
 sg13g2_buf_1 place8188 (.A(net8188),
    .X(net8187));
 sg13g2_buf_1 place8189 (.A(net8206),
    .X(net8188));
 sg13g2_buf_1 place8190 (.A(net8206),
    .X(net8189));
 sg13g2_buf_1 place8191 (.A(net8191),
    .X(net8190));
 sg13g2_buf_1 place8192 (.A(net8206),
    .X(net8191));
 sg13g2_buf_1 place8193 (.A(net8206),
    .X(net8192));
 sg13g2_buf_1 place8194 (.A(net8205),
    .X(net8193));
 sg13g2_buf_1 place8195 (.A(net8195),
    .X(net8194));
 sg13g2_buf_1 place8196 (.A(net8205),
    .X(net8195));
 sg13g2_buf_1 place8197 (.A(net8205),
    .X(net8196));
 sg13g2_buf_1 place8198 (.A(net8198),
    .X(net8197));
 sg13g2_buf_1 place8199 (.A(net8204),
    .X(net8198));
 sg13g2_buf_1 place8200 (.A(net8204),
    .X(net8199));
 sg13g2_buf_1 place8201 (.A(net8203),
    .X(net8200));
 sg13g2_buf_1 place8202 (.A(net8202),
    .X(net8201));
 sg13g2_buf_1 place8203 (.A(net8203),
    .X(net8202));
 sg13g2_buf_1 place8204 (.A(net8204),
    .X(net8203));
 sg13g2_buf_1 place8205 (.A(net8205),
    .X(net8204));
 sg13g2_buf_1 place8206 (.A(net8206),
    .X(net8205));
 sg13g2_buf_1 place8207 (.A(net8207),
    .X(net8206));
 sg13g2_buf_4 place8208 (.X(net8207),
    .A(net437));
 sg13g2_buf_1 place8209 (.A(net8226),
    .X(net8208));
 sg13g2_buf_1 place8210 (.A(net8212),
    .X(net8209));
 sg13g2_buf_1 place8211 (.A(net8212),
    .X(net8210));
 sg13g2_buf_1 place8212 (.A(net8212),
    .X(net8211));
 sg13g2_buf_1 place8213 (.A(net8213),
    .X(net8212));
 sg13g2_buf_1 place8214 (.A(net8226),
    .X(net8213));
 sg13g2_buf_1 place8215 (.A(net8215),
    .X(net8214));
 sg13g2_buf_1 place8216 (.A(net8225),
    .X(net8215));
 sg13g2_buf_1 place8217 (.A(net8225),
    .X(net8216));
 sg13g2_buf_1 place8218 (.A(net8219),
    .X(net8217));
 sg13g2_buf_1 place8219 (.A(net8219),
    .X(net8218));
 sg13g2_buf_1 place8220 (.A(net8225),
    .X(net8219));
 sg13g2_buf_1 place8221 (.A(net8224),
    .X(net8220));
 sg13g2_buf_1 place8222 (.A(net8222),
    .X(net8221));
 sg13g2_buf_1 place8223 (.A(net8223),
    .X(net8222));
 sg13g2_buf_1 place8224 (.A(net8224),
    .X(net8223));
 sg13g2_buf_1 place8225 (.A(net8225),
    .X(net8224));
 sg13g2_buf_1 place8226 (.A(net8226),
    .X(net8225));
 sg13g2_buf_1 place8227 (.A(net8285),
    .X(net8226));
 sg13g2_buf_1 place8228 (.A(net8228),
    .X(net8227));
 sg13g2_buf_1 place8229 (.A(net8237),
    .X(net8228));
 sg13g2_buf_1 place8230 (.A(net8235),
    .X(net8229));
 sg13g2_buf_1 place8231 (.A(net8231),
    .X(net8230));
 sg13g2_buf_1 place8232 (.A(net8232),
    .X(net8231));
 sg13g2_buf_1 place8233 (.A(net8233),
    .X(net8232));
 sg13g2_buf_1 place8234 (.A(net8234),
    .X(net8233));
 sg13g2_buf_1 place8235 (.A(net8235),
    .X(net8234));
 sg13g2_buf_1 place8236 (.A(net8236),
    .X(net8235));
 sg13g2_buf_1 place8237 (.A(net8237),
    .X(net8236));
 sg13g2_buf_1 place8238 (.A(net8285),
    .X(net8237));
 sg13g2_buf_1 place8239 (.A(net8284),
    .X(net8238));
 sg13g2_buf_1 place8240 (.A(net8240),
    .X(net8239));
 sg13g2_buf_1 place8241 (.A(net8242),
    .X(net8240));
 sg13g2_buf_1 place8242 (.A(net8242),
    .X(net8241));
 sg13g2_buf_1 place8243 (.A(net8284),
    .X(net8242));
 sg13g2_buf_1 place8244 (.A(net8252),
    .X(net8243));
 sg13g2_buf_1 place8245 (.A(net8252),
    .X(net8244));
 sg13g2_buf_1 place8246 (.A(net8246),
    .X(net8245));
 sg13g2_buf_1 place8247 (.A(net8252),
    .X(net8246));
 sg13g2_buf_1 place8248 (.A(net8252),
    .X(net8247));
 sg13g2_buf_1 place8249 (.A(net8251),
    .X(net8248));
 sg13g2_buf_1 place8250 (.A(net8250),
    .X(net8249));
 sg13g2_buf_1 place8251 (.A(net8251),
    .X(net8250));
 sg13g2_buf_1 place8252 (.A(net8252),
    .X(net8251));
 sg13g2_buf_1 place8253 (.A(net8283),
    .X(net8252));
 sg13g2_buf_1 place8254 (.A(net8256),
    .X(net8253));
 sg13g2_buf_1 place8255 (.A(net8256),
    .X(net8254));
 sg13g2_buf_1 place8256 (.A(net8256),
    .X(net8255));
 sg13g2_buf_1 place8257 (.A(net8257),
    .X(net8256));
 sg13g2_buf_1 place8258 (.A(net8283),
    .X(net8257));
 sg13g2_buf_1 place8259 (.A(net8282),
    .X(net8258));
 sg13g2_buf_1 place8260 (.A(net8260),
    .X(net8259));
 sg13g2_buf_1 place8261 (.A(net8282),
    .X(net8260));
 sg13g2_buf_1 place8262 (.A(net8266),
    .X(net8261));
 sg13g2_buf_1 place8263 (.A(net8265),
    .X(net8262));
 sg13g2_buf_1 place8264 (.A(net8264),
    .X(net8263));
 sg13g2_buf_1 place8265 (.A(net8265),
    .X(net8264));
 sg13g2_buf_1 place8266 (.A(net8266),
    .X(net8265));
 sg13g2_buf_1 place8267 (.A(net8282),
    .X(net8266));
 sg13g2_buf_1 place8268 (.A(net8282),
    .X(net8267));
 sg13g2_buf_1 place8269 (.A(net8269),
    .X(net8268));
 sg13g2_buf_1 place8270 (.A(net8281),
    .X(net8269));
 sg13g2_buf_1 place8271 (.A(net8271),
    .X(net8270));
 sg13g2_buf_1 place8272 (.A(net8273),
    .X(net8271));
 sg13g2_buf_1 place8273 (.A(net8273),
    .X(net8272));
 sg13g2_buf_1 place8274 (.A(net8281),
    .X(net8273));
 sg13g2_buf_1 place8275 (.A(net8275),
    .X(net8274));
 sg13g2_buf_1 place8276 (.A(net8280),
    .X(net8275));
 sg13g2_buf_1 place8277 (.A(net8279),
    .X(net8276));
 sg13g2_buf_1 place8278 (.A(net8279),
    .X(net8277));
 sg13g2_buf_1 place8279 (.A(net8279),
    .X(net8278));
 sg13g2_buf_1 place8280 (.A(net8280),
    .X(net8279));
 sg13g2_buf_1 place8281 (.A(net8281),
    .X(net8280));
 sg13g2_buf_1 place8282 (.A(net8282),
    .X(net8281));
 sg13g2_buf_1 place8283 (.A(net8283),
    .X(net8282));
 sg13g2_buf_1 place8284 (.A(net8284),
    .X(net8283));
 sg13g2_buf_1 place8285 (.A(net8285),
    .X(net8284));
 sg13g2_buf_2 place8286 (.A(net437),
    .X(net8285));
endmodule
module \ALU_33_0_33_0_33_unused_CO_X_Y[0]_KOGGE_STONE  (A,
    B,
    BI,
    CI,
    \Y[32:1] );
 input [32:0] A;
 input [32:0] B;
 input BI;
 input CI;
 output [31:0] \Y[32:1] ;

 wire _203_;
 wire _202_;
 wire _201_;
 wire _200_;
 wire _199_;
 wire _198_;
 wire _197_;
 wire _196_;
 wire _195_;
 wire _194_;
 wire _193_;
 wire _192_;
 wire _191_;
 wire _190_;
 wire _189_;
 wire _188_;
 wire _187_;
 wire _186_;
 wire _185_;
 wire _184_;
 wire _183_;
 wire _182_;
 wire _181_;
 wire _180_;
 wire _179_;
 wire _178_;
 wire _177_;
 wire _176_;
 wire _175_;
 wire _174_;
 wire _173_;
 wire _172_;
 wire _171_;
 wire _170_;
 wire _169_;
 wire _168_;
 wire _167_;
 wire _166_;
 wire _165_;
 wire _164_;
 wire _163_;
 wire _162_;
 wire _161_;
 wire _160_;
 wire _159_;
 wire _158_;
 wire _157_;
 wire _156_;
 wire _155_;
 wire _154_;
 wire _153_;
 wire _152_;
 wire _151_;
 wire _150_;
 wire _149_;
 wire _148_;
 wire _147_;
 wire _146_;
 wire _145_;
 wire _144_;
 wire _143_;
 wire _142_;
 wire _141_;
 wire _140_;
 wire _139_;
 wire _138_;
 wire _137_;
 wire _136_;
 wire _135_;
 wire _134_;
 wire _133_;
 wire _132_;
 wire _131_;
 wire _130_;
 wire _129_;
 wire _128_;
 wire _127_;
 wire _126_;
 wire _125_;
 wire _124_;
 wire _123_;
 wire _122_;
 wire _121_;
 wire _120_;
 wire _119_;
 wire _118_;
 wire _117_;
 wire _116_;
 wire _115_;
 wire _114_;
 wire _113_;
 wire _112_;
 wire _111_;
 wire _110_;
 wire _109_;
 wire _108_;
 wire _107_;
 wire _106_;
 wire _105_;
 wire _104_;
 wire _103_;
 wire _102_;
 wire _101_;
 wire _100_;
 wire _099_;
 wire _098_;
 wire _097_;
 wire _096_;
 wire _095_;
 wire _094_;
 wire _093_;
 wire _092_;
 wire _091_;
 wire _090_;
 wire _089_;
 wire _088_;
 wire _307_;
 wire _087_;
 wire _086_;
 wire _085_;
 wire _084_;
 wire _083_;
 wire _082_;
 wire _081_;
 wire _080_;
 wire _079_;
 wire _078_;
 wire _077_;
 wire _076_;
 wire _075_;
 wire _074_;
 wire _297_;
 wire _073_;
 wire _072_;
 wire _071_;
 wire _070_;
 wire _069_;
 wire _068_;
 wire _067_;
 wire _066_;
 wire _065_;
 wire _064_;
 wire _063_;
 wire _062_;
 wire _061_;
 wire _284_;
 wire _060_;
 wire _059_;
 wire _058_;
 wire _057_;
 wire _056_;
 wire _055_;
 wire _054_;
 wire _053_;
 wire _052_;
 wire _051_;
 wire _275_;
 wire _050_;
 wire _049_;
 wire _048_;
 wire _047_;
 wire _046_;
 wire _045_;
 wire _044_;
 wire _043_;
 wire _042_;
 wire _041_;
 wire _040_;
 wire _265_;
 wire _039_;
 wire _304_;
 wire _303_;
 wire _038_;
 wire _037_;
 wire _036_;
 wire _035_;
 wire _034_;
 wire _033_;
 wire _032_;
 wire _031_;
 wire _030_;
 wire _029_;
 wire _257_;
 wire _028_;
 wire _294_;
 wire _293_;
 wire _027_;
 wire _026_;
 wire _025_;
 wire _024_;
 wire _023_;
 wire _022_;
 wire _021_;
 wire _020_;
 wire _019_;
 wire _018_;
 wire _249_;
 wire _017_;
 wire _281_;
 wire _016_;
 wire _302_;
 wire _015_;
 wire _282_;
 wire _014_;
 wire _013_;
 wire _012_;
 wire _287_;
 wire _011_;
 wire _010_;
 wire _241_;
 wire _009_;
 wire _273_;
 wire _008_;
 wire _271_;
 wire _007_;
 wire _006_;
 wire _291_;
 wire _005_;
 wire _292_;
 wire _289_;
 wire _004_;
 wire _299_;
 wire _003_;
 wire _300_;
 wire _290_;
 wire _002_;
 wire _001_;
 wire _000_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _272_;
 wire _274_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _283_;
 wire _285_;
 wire _286_;
 wire _288_;
 wire _295_;
 wire _296_;
 wire _298_;
 wire _301_;
 wire _305_;
 wire _306_;

 sg13g2_xor2_1 _308_ (.B(BI),
    .A(B[15]),
    .X(_000_));
 sg13g2_nand2_1 _309_ (.Y(_001_),
    .A(A[15]),
    .B(_000_));
 sg13g2_xnor2_1 _310_ (.Y(_002_),
    .A(A[15]),
    .B(_000_));
 sg13g2_nor2_1 _311_ (.A(_290_),
    .B(_300_),
    .Y(_003_));
 sg13g2_o21ai_1 _312_ (.B1(_299_),
    .Y(_004_),
    .A1(_289_),
    .A2(_300_));
 sg13g2_a21o_1 _313_ (.A2(_003_),
    .A1(_292_),
    .B1(_004_),
    .X(_005_));
 sg13g2_and2_1 _314_ (.A(_291_),
    .B(_003_),
    .X(_006_));
 sg13g2_nand2_1 _315_ (.Y(_007_),
    .A(_291_),
    .B(_003_));
 sg13g2_a21o_1 _316_ (.A2(_006_),
    .A1(_271_),
    .B1(_005_),
    .X(_008_));
 sg13g2_nor2_1 _317_ (.A(_273_),
    .B(_007_),
    .Y(_009_));
 sg13g2_a21oi_1 _318_ (.A1(_241_),
    .A2(_009_),
    .Y(_010_),
    .B1(_008_));
 sg13g2_xor2_1 _319_ (.B(_010_),
    .A(_002_),
    .X(\Y[32:1] [14]));
 sg13g2_nor2_1 _320_ (.A(_300_),
    .B(_002_),
    .Y(_011_));
 sg13g2_nor4_1 _321_ (.A(_287_),
    .B(_290_),
    .C(_300_),
    .D(_002_),
    .Y(_012_));
 sg13g2_inv_1 _322_ (.Y(_013_),
    .A(_014_));
 sg13g2_nand2_1 _323_ (.Y(_014_),
    .A(_282_),
    .B(_012_));
 sg13g2_o21ai_1 _324_ (.B1(_001_),
    .Y(_015_),
    .A1(_299_),
    .A2(_002_));
 sg13g2_a21o_1 _325_ (.A2(_011_),
    .A1(_302_),
    .B1(_015_),
    .X(_016_));
 sg13g2_a21o_1 _326_ (.A2(_012_),
    .A1(_281_),
    .B1(_016_),
    .X(_017_));
 sg13g2_a21oi_1 _327_ (.A1(_249_),
    .A2(_013_),
    .Y(_018_),
    .B1(_017_));
 sg13g2_xor2_1 _328_ (.B(BI),
    .A(B[16]),
    .X(_019_));
 sg13g2_nand2_1 _329_ (.Y(_020_),
    .A(A[16]),
    .B(_019_));
 sg13g2_xnor2_1 _330_ (.Y(_021_),
    .A(A[16]),
    .B(_019_));
 sg13g2_xor2_1 _331_ (.B(_021_),
    .A(_018_),
    .X(\Y[32:1] [15]));
 sg13g2_nor2_1 _332_ (.A(_002_),
    .B(_021_),
    .Y(_022_));
 sg13g2_nand2_1 _333_ (.Y(_023_),
    .A(_003_),
    .B(_022_));
 sg13g2_o21ai_1 _334_ (.B1(_020_),
    .Y(_024_),
    .A1(_001_),
    .A2(_021_));
 sg13g2_a21oi_1 _335_ (.A1(_004_),
    .A2(_022_),
    .Y(_025_),
    .B1(_024_));
 sg13g2_inv_1 _336_ (.Y(_026_),
    .A(_025_));
 sg13g2_o21ai_1 _337_ (.B1(_025_),
    .Y(_027_),
    .A1(_293_),
    .A2(_023_));
 sg13g2_nor2_1 _338_ (.A(_294_),
    .B(_023_),
    .Y(_028_));
 sg13g2_a21oi_1 _339_ (.A1(_257_),
    .A2(_028_),
    .Y(_029_),
    .B1(_027_));
 sg13g2_xor2_1 _340_ (.B(BI),
    .A(B[17]),
    .X(_030_));
 sg13g2_nand2_1 _341_ (.Y(_031_),
    .A(A[17]),
    .B(_030_));
 sg13g2_xnor2_1 _342_ (.Y(_032_),
    .A(A[17]),
    .B(_030_));
 sg13g2_xor2_1 _343_ (.B(_032_),
    .A(_029_),
    .X(\Y[32:1] [16]));
 sg13g2_nor2_1 _344_ (.A(_021_),
    .B(_032_),
    .Y(_033_));
 sg13g2_nand2_1 _345_ (.Y(_034_),
    .A(_011_),
    .B(_033_));
 sg13g2_o21ai_1 _346_ (.B1(_031_),
    .Y(_035_),
    .A1(_020_),
    .A2(_032_));
 sg13g2_a21oi_1 _347_ (.A1(_015_),
    .A2(_033_),
    .Y(_036_),
    .B1(_035_));
 sg13g2_inv_1 _348_ (.Y(_037_),
    .A(_036_));
 sg13g2_o21ai_1 _349_ (.B1(_036_),
    .Y(_038_),
    .A1(_303_),
    .A2(_034_));
 sg13g2_nor2_1 _350_ (.A(_304_),
    .B(_034_),
    .Y(_039_));
 sg13g2_a21oi_1 _351_ (.A1(_265_),
    .A2(_039_),
    .Y(_040_),
    .B1(_038_));
 sg13g2_xor2_1 _352_ (.B(BI),
    .A(B[18]),
    .X(_041_));
 sg13g2_nand2_1 _353_ (.Y(_042_),
    .A(A[18]),
    .B(_041_));
 sg13g2_xnor2_1 _354_ (.Y(_043_),
    .A(A[18]),
    .B(_041_));
 sg13g2_xor2_1 _355_ (.B(_043_),
    .A(_040_),
    .X(\Y[32:1] [17]));
 sg13g2_nor2_1 _356_ (.A(_032_),
    .B(_043_),
    .Y(_044_));
 sg13g2_nor4_1 _357_ (.A(_002_),
    .B(_021_),
    .C(_032_),
    .D(_043_),
    .Y(_045_));
 sg13g2_o21ai_1 _358_ (.B1(_042_),
    .Y(_046_),
    .A1(_031_),
    .A2(_043_));
 sg13g2_a21oi_1 _359_ (.A1(_024_),
    .A2(_044_),
    .Y(_047_),
    .B1(_046_));
 sg13g2_a221oi_1 _360_ (.B2(_005_),
    .C1(_046_),
    .B1(_045_),
    .A1(_024_),
    .Y(_048_),
    .A2(_044_));
 sg13g2_nand3_1 _361_ (.B(_003_),
    .C(_045_),
    .A(_291_),
    .Y(_049_));
 sg13g2_o21ai_1 _362_ (.B1(_048_),
    .Y(_050_),
    .A1(_275_),
    .A2(_049_));
 sg13g2_xor2_1 _363_ (.B(BI),
    .A(B[19]),
    .X(_051_));
 sg13g2_nand2_1 _364_ (.Y(_052_),
    .A(A[19]),
    .B(_051_));
 sg13g2_xnor2_1 _365_ (.Y(_053_),
    .A(A[19]),
    .B(_051_));
 sg13g2_xnor2_1 _366_ (.Y(\Y[32:1] [18]),
    .A(_050_),
    .B(_053_));
 sg13g2_nor2_1 _367_ (.A(_043_),
    .B(_053_),
    .Y(_054_));
 sg13g2_o21ai_1 _368_ (.B1(_052_),
    .Y(_055_),
    .A1(_042_),
    .A2(_053_));
 sg13g2_a21oi_1 _369_ (.A1(_035_),
    .A2(_054_),
    .Y(_056_),
    .B1(_055_));
 sg13g2_nor4_1 _370_ (.A(_021_),
    .B(_032_),
    .C(_043_),
    .D(_053_),
    .Y(_057_));
 sg13g2_a221oi_1 _371_ (.B2(_016_),
    .C1(_055_),
    .B1(_057_),
    .A1(_035_),
    .Y(_058_),
    .A2(_054_));
 sg13g2_nand2_1 _372_ (.Y(_059_),
    .A(_012_),
    .B(_057_));
 sg13g2_o21ai_1 _373_ (.B1(_058_),
    .Y(_060_),
    .A1(_284_),
    .A2(_059_));
 sg13g2_xor2_1 _374_ (.B(BI),
    .A(B[20]),
    .X(_061_));
 sg13g2_nand2_1 _375_ (.Y(_062_),
    .A(A[20]),
    .B(_061_));
 sg13g2_xnor2_1 _376_ (.Y(_063_),
    .A(A[20]),
    .B(_061_));
 sg13g2_xnor2_1 _377_ (.Y(\Y[32:1] [19]),
    .A(_060_),
    .B(_063_));
 sg13g2_nor2_1 _378_ (.A(_053_),
    .B(_063_),
    .Y(_064_));
 sg13g2_o21ai_1 _379_ (.B1(_062_),
    .Y(_065_),
    .A1(_052_),
    .A2(_063_));
 sg13g2_a21oi_1 _380_ (.A1(_046_),
    .A2(_064_),
    .Y(_066_),
    .B1(_065_));
 sg13g2_a21o_1 _381_ (.A2(_064_),
    .A1(_046_),
    .B1(_065_),
    .X(_067_));
 sg13g2_nor4_1 _382_ (.A(_032_),
    .B(_043_),
    .C(_053_),
    .D(_063_),
    .Y(_068_));
 sg13g2_inv_1 _383_ (.Y(_069_),
    .A(_068_));
 sg13g2_a21oi_1 _384_ (.A1(_026_),
    .A2(_068_),
    .Y(_070_),
    .B1(_067_));
 sg13g2_o21ai_1 _385_ (.B1(_066_),
    .Y(_071_),
    .A1(_025_),
    .A2(_069_));
 sg13g2_nand3_1 _386_ (.B(_022_),
    .C(_068_),
    .A(_003_),
    .Y(_072_));
 sg13g2_o21ai_1 _387_ (.B1(_070_),
    .Y(_073_),
    .A1(_297_),
    .A2(_072_));
 sg13g2_xor2_1 _388_ (.B(BI),
    .A(B[21]),
    .X(_074_));
 sg13g2_nand2_1 _389_ (.Y(_075_),
    .A(A[21]),
    .B(_074_));
 sg13g2_xnor2_1 _390_ (.Y(_076_),
    .A(A[21]),
    .B(_074_));
 sg13g2_xnor2_1 _391_ (.Y(\Y[32:1] [20]),
    .A(_073_),
    .B(_076_));
 sg13g2_nor2_1 _392_ (.A(_063_),
    .B(_076_),
    .Y(_077_));
 sg13g2_xor2_1 _393_ (.B(BI),
    .A(B[1]),
    .X(_078_));
 sg13g2_o21ai_1 _394_ (.B1(_075_),
    .Y(_079_),
    .A1(_062_),
    .A2(_076_));
 sg13g2_a21oi_1 _395_ (.A1(_055_),
    .A2(_077_),
    .Y(_080_),
    .B1(_079_));
 sg13g2_a21o_1 _396_ (.A2(_077_),
    .A1(_055_),
    .B1(_079_),
    .X(_081_));
 sg13g2_nor4_1 _397_ (.A(_043_),
    .B(_053_),
    .C(_063_),
    .D(_076_),
    .Y(_082_));
 sg13g2_inv_1 _398_ (.Y(_083_),
    .A(_082_));
 sg13g2_a21oi_1 _399_ (.A1(_037_),
    .A2(_082_),
    .Y(_084_),
    .B1(_081_));
 sg13g2_o21ai_1 _400_ (.B1(_080_),
    .Y(_085_),
    .A1(_036_),
    .A2(_083_));
 sg13g2_nand3_1 _401_ (.B(_033_),
    .C(_082_),
    .A(_011_),
    .Y(_086_));
 sg13g2_o21ai_1 _402_ (.B1(_084_),
    .Y(_087_),
    .A1(_307_),
    .A2(_086_));
 sg13g2_nand2_1 _403_ (.Y(_088_),
    .A(A[1]),
    .B(_078_));
 sg13g2_xor2_1 _404_ (.B(BI),
    .A(B[22]),
    .X(_089_));
 sg13g2_nand2_1 _405_ (.Y(_090_),
    .A(A[22]),
    .B(_089_));
 sg13g2_xnor2_1 _406_ (.Y(_091_),
    .A(A[22]),
    .B(_089_));
 sg13g2_xnor2_1 _407_ (.Y(\Y[32:1] [21]),
    .A(_087_),
    .B(_091_));
 sg13g2_nor2_1 _408_ (.A(_076_),
    .B(_091_),
    .Y(_092_));
 sg13g2_o21ai_1 _409_ (.B1(_090_),
    .Y(_093_),
    .A1(_075_),
    .A2(_091_));
 sg13g2_a21oi_1 _410_ (.A1(_065_),
    .A2(_092_),
    .Y(_094_),
    .B1(_093_));
 sg13g2_nand2_1 _411_ (.Y(_095_),
    .A(_064_),
    .B(_092_));
 sg13g2_o21ai_1 _412_ (.B1(_094_),
    .Y(_096_),
    .A1(_047_),
    .A2(_095_));
 sg13g2_inv_1 _413_ (.Y(_097_),
    .A(_098_));
 sg13g2_nand3_1 _414_ (.B(_064_),
    .C(_092_),
    .A(_045_),
    .Y(_098_));
 sg13g2_nor3_1 _415_ (.A(_273_),
    .B(_007_),
    .C(_098_),
    .Y(_099_));
 sg13g2_a221oi_1 _416_ (.B2(_241_),
    .C1(_096_),
    .B1(_099_),
    .A1(_008_),
    .Y(_100_),
    .A2(_097_));
 sg13g2_xor2_1 _417_ (.B(BI),
    .A(B[23]),
    .X(_101_));
 sg13g2_nand2_1 _418_ (.Y(_102_),
    .A(A[23]),
    .B(_101_));
 sg13g2_xnor2_1 _419_ (.Y(_103_),
    .A(A[23]),
    .B(_101_));
 sg13g2_xnor2_1 _420_ (.Y(_104_),
    .A(A[1]),
    .B(_078_));
 sg13g2_xor2_1 _421_ (.B(_103_),
    .A(_100_),
    .X(\Y[32:1] [22]));
 sg13g2_nor2_1 _422_ (.A(_091_),
    .B(_103_),
    .Y(_105_));
 sg13g2_o21ai_1 _423_ (.B1(_102_),
    .Y(_106_),
    .A1(_090_),
    .A2(_103_));
 sg13g2_a21oi_1 _424_ (.A1(_079_),
    .A2(_105_),
    .Y(_107_),
    .B1(_106_));
 sg13g2_nor4_1 _425_ (.A(_063_),
    .B(_076_),
    .C(_091_),
    .D(_103_),
    .Y(_108_));
 sg13g2_inv_1 _426_ (.Y(_109_),
    .A(_108_));
 sg13g2_nand2_1 _427_ (.Y(_110_),
    .A(A[0]),
    .B(CI));
 sg13g2_o21ai_1 _428_ (.B1(_107_),
    .Y(_111_),
    .A1(_056_),
    .A2(_109_));
 sg13g2_inv_1 _429_ (.Y(_112_),
    .A(_113_));
 sg13g2_nand2_1 _430_ (.Y(_113_),
    .A(_057_),
    .B(_108_));
 sg13g2_nor2_1 _431_ (.A(_014_),
    .B(_113_),
    .Y(_114_));
 sg13g2_a221oi_1 _432_ (.B2(_249_),
    .C1(_111_),
    .B1(_114_),
    .A1(_017_),
    .Y(_115_),
    .A2(_112_));
 sg13g2_xor2_1 _433_ (.B(BI),
    .A(B[24]),
    .X(_116_));
 sg13g2_nand2_1 _434_ (.Y(_117_),
    .A(A[24]),
    .B(_116_));
 sg13g2_xnor2_1 _435_ (.Y(_118_),
    .A(A[24]),
    .B(_116_));
 sg13g2_xor2_1 _436_ (.B(_118_),
    .A(_115_),
    .X(\Y[32:1] [23]));
 sg13g2_nor2_1 _437_ (.A(_103_),
    .B(_118_),
    .Y(_119_));
 sg13g2_o21ai_1 _438_ (.B1(_117_),
    .Y(_120_),
    .A1(_102_),
    .A2(_118_));
 sg13g2_a21o_1 _439_ (.A2(_119_),
    .A1(_093_),
    .B1(_120_),
    .X(_121_));
 sg13g2_and2_1 _440_ (.A(_092_),
    .B(_119_),
    .X(_122_));
 sg13g2_a21oi_1 _441_ (.A1(_067_),
    .A2(_122_),
    .Y(_123_),
    .B1(_121_));
 sg13g2_nand2_1 _442_ (.Y(_124_),
    .A(_068_),
    .B(_122_));
 sg13g2_o21ai_1 _443_ (.B1(_123_),
    .Y(_125_),
    .A1(_029_),
    .A2(_124_));
 sg13g2_xor2_1 _444_ (.B(BI),
    .A(B[25]),
    .X(_126_));
 sg13g2_nand2_1 _445_ (.Y(_127_),
    .A(A[25]),
    .B(_126_));
 sg13g2_xnor2_1 _446_ (.Y(_128_),
    .A(B[0]),
    .B(BI));
 sg13g2_xnor2_1 _447_ (.Y(_129_),
    .A(A[25]),
    .B(_126_));
 sg13g2_xnor2_1 _448_ (.Y(\Y[32:1] [24]),
    .A(_125_),
    .B(_129_));
 sg13g2_nor2_1 _449_ (.A(_118_),
    .B(_129_),
    .Y(_130_));
 sg13g2_nor2_1 _450_ (.A(A[0]),
    .B(CI),
    .Y(_131_));
 sg13g2_o21ai_1 _451_ (.B1(_127_),
    .Y(_132_),
    .A1(_117_),
    .A2(_129_));
 sg13g2_a21oi_1 _452_ (.A1(_106_),
    .A2(_130_),
    .Y(_133_),
    .B1(_132_));
 sg13g2_and2_1 _453_ (.A(_105_),
    .B(_130_),
    .X(_134_));
 sg13g2_a221oi_1 _454_ (.B2(_081_),
    .C1(_132_),
    .B1(_134_),
    .A1(_106_),
    .Y(_135_),
    .A2(_130_));
 sg13g2_nand2_1 _455_ (.Y(_136_),
    .A(_082_),
    .B(_134_));
 sg13g2_o21ai_1 _456_ (.B1(_135_),
    .Y(_137_),
    .A1(_040_),
    .A2(_136_));
 sg13g2_xor2_1 _457_ (.B(BI),
    .A(B[26]),
    .X(_138_));
 sg13g2_nand2_1 _458_ (.Y(_139_),
    .A(A[26]),
    .B(_138_));
 sg13g2_xnor2_1 _459_ (.Y(_140_),
    .A(A[26]),
    .B(_138_));
 sg13g2_xnor2_1 _460_ (.Y(\Y[32:1] [25]),
    .A(_137_),
    .B(_140_));
 sg13g2_nor2_1 _461_ (.A(_129_),
    .B(_140_),
    .Y(_141_));
 sg13g2_o21ai_1 _462_ (.B1(_139_),
    .Y(_142_),
    .A1(_127_),
    .A2(_140_));
 sg13g2_a21oi_1 _463_ (.A1(_120_),
    .A2(_141_),
    .Y(_143_),
    .B1(_142_));
 sg13g2_nand2_1 _464_ (.Y(_144_),
    .A(_119_),
    .B(_141_));
 sg13g2_o21ai_1 _465_ (.B1(_143_),
    .Y(_145_),
    .A1(_094_),
    .A2(_144_));
 sg13g2_nor2_1 _466_ (.A(_095_),
    .B(_144_),
    .Y(_146_));
 sg13g2_a21oi_1 _467_ (.A1(_050_),
    .A2(_146_),
    .Y(_147_),
    .B1(_145_));
 sg13g2_xor2_1 _468_ (.B(BI),
    .A(B[27]),
    .X(_148_));
 sg13g2_nand2_1 _469_ (.Y(_149_),
    .A(A[27]),
    .B(_148_));
 sg13g2_xnor2_1 _470_ (.Y(_150_),
    .A(A[27]),
    .B(_148_));
 sg13g2_xor2_1 _471_ (.B(_150_),
    .A(_147_),
    .X(\Y[32:1] [26]));
 sg13g2_nor2_1 _472_ (.A(_140_),
    .B(_150_),
    .Y(_151_));
 sg13g2_o21ai_1 _473_ (.B1(_149_),
    .Y(_152_),
    .A1(_139_),
    .A2(_150_));
 sg13g2_a21oi_1 _474_ (.A1(_132_),
    .A2(_151_),
    .Y(_153_),
    .B1(_152_));
 sg13g2_and2_1 _475_ (.A(_130_),
    .B(_151_),
    .X(_154_));
 sg13g2_inv_1 _476_ (.Y(_155_),
    .A(_154_));
 sg13g2_o21ai_1 _477_ (.B1(_153_),
    .Y(_156_),
    .A1(_107_),
    .A2(_155_));
 sg13g2_nor2_1 _478_ (.A(_109_),
    .B(_155_),
    .Y(_157_));
 sg13g2_a21oi_1 _479_ (.A1(_060_),
    .A2(_157_),
    .Y(_158_),
    .B1(_156_));
 sg13g2_xor2_1 _480_ (.B(BI),
    .A(B[28]),
    .X(_159_));
 sg13g2_nand2_1 _481_ (.Y(_160_),
    .A(A[28]),
    .B(_159_));
 sg13g2_a21o_1 _482_ (.A2(_128_),
    .A1(_110_),
    .B1(_131_),
    .X(_161_));
 sg13g2_xnor2_1 _483_ (.Y(_162_),
    .A(A[28]),
    .B(_159_));
 sg13g2_a21oi_1 _484_ (.A1(_110_),
    .A2(_128_),
    .Y(_163_),
    .B1(_131_));
 sg13g2_xor2_1 _485_ (.B(_162_),
    .A(_158_),
    .X(\Y[32:1] [27]));
 sg13g2_inv_1 _486_ (.Y(_164_),
    .A(_165_));
 sg13g2_o21ai_1 _487_ (.B1(_160_),
    .Y(_165_),
    .A1(_149_),
    .A2(_162_));
 sg13g2_nor2_1 _488_ (.A(_150_),
    .B(_162_),
    .Y(_166_));
 sg13g2_inv_1 _489_ (.Y(_167_),
    .A(_166_));
 sg13g2_a21o_1 _490_ (.A2(_141_),
    .A1(_121_),
    .B1(_142_),
    .X(_168_));
 sg13g2_and3_1 _491_ (.X(_169_),
    .A(_122_),
    .B(_141_),
    .C(_166_));
 sg13g2_a221oi_1 _492_ (.B2(_071_),
    .C1(_165_),
    .B1(_169_),
    .A1(_166_),
    .Y(_170_),
    .A2(_168_));
 sg13g2_nand2b_1 _493_ (.Y(_171_),
    .B(_169_),
    .A_N(_072_));
 sg13g2_o21ai_1 _494_ (.B1(_170_),
    .Y(_172_),
    .A1(_297_),
    .A2(_171_));
 sg13g2_xor2_1 _495_ (.B(BI),
    .A(B[29]),
    .X(_173_));
 sg13g2_nand2_1 _496_ (.Y(_174_),
    .A(A[29]),
    .B(_173_));
 sg13g2_xnor2_1 _497_ (.Y(_175_),
    .A(A[29]),
    .B(_173_));
 sg13g2_xnor2_1 _498_ (.Y(\Y[32:1] [28]),
    .A(_172_),
    .B(_175_));
 sg13g2_inv_1 _499_ (.Y(_176_),
    .A(_177_));
 sg13g2_o21ai_1 _500_ (.B1(_174_),
    .Y(_177_),
    .A1(_160_),
    .A2(_175_));
 sg13g2_nor2_1 _501_ (.A(_162_),
    .B(_175_),
    .Y(_178_));
 sg13g2_or2_1 _502_ (.X(_179_),
    .B(_175_),
    .A(_162_));
 sg13g2_nand2_1 _503_ (.Y(_180_),
    .A(_151_),
    .B(_178_));
 sg13g2_o21ai_1 _504_ (.B1(_176_),
    .Y(_181_),
    .A1(_133_),
    .A2(_180_));
 sg13g2_xnor2_1 _505_ (.Y(\Y[32:1] [0]),
    .A(_104_),
    .B(_163_));
 sg13g2_and3_1 _506_ (.X(_182_),
    .A(_134_),
    .B(_151_),
    .C(_178_));
 sg13g2_a221oi_1 _507_ (.B2(_085_),
    .C1(_181_),
    .B1(_182_),
    .A1(_152_),
    .Y(_183_),
    .A2(_178_));
 sg13g2_nand2b_1 _508_ (.Y(_184_),
    .B(_182_),
    .A_N(_086_));
 sg13g2_o21ai_1 _509_ (.B1(_183_),
    .Y(_185_),
    .A1(_307_),
    .A2(_184_));
 sg13g2_o21ai_1 _510_ (.B1(_088_),
    .Y(_186_),
    .A1(_104_),
    .A2(_161_));
 sg13g2_xor2_1 _511_ (.B(BI),
    .A(B[30]),
    .X(_187_));
 sg13g2_nand2_1 _512_ (.Y(_188_),
    .A(A[30]),
    .B(_187_));
 sg13g2_xnor2_1 _513_ (.Y(_189_),
    .A(A[30]),
    .B(_187_));
 sg13g2_xnor2_1 _514_ (.Y(\Y[32:1] [29]),
    .A(_185_),
    .B(_189_));
 sg13g2_o21ai_1 _515_ (.B1(_188_),
    .Y(_190_),
    .A1(_174_),
    .A2(_189_));
 sg13g2_nor2_1 _516_ (.A(_175_),
    .B(_189_),
    .Y(_191_));
 sg13g2_o21ai_1 _517_ (.B1(_164_),
    .Y(_192_),
    .A1(_143_),
    .A2(_167_));
 sg13g2_a21oi_1 _518_ (.A1(_191_),
    .A2(_192_),
    .Y(_193_),
    .B1(_190_));
 sg13g2_nand4_1 _519_ (.B(_141_),
    .C(_166_),
    .A(_119_),
    .Y(_194_),
    .D(_191_));
 sg13g2_o21ai_1 _520_ (.B1(_193_),
    .Y(_195_),
    .A1(_100_),
    .A2(_194_));
 sg13g2_xor2_1 _521_ (.B(BI),
    .A(B[31]),
    .X(_196_));
 sg13g2_xnor2_1 _522_ (.Y(_197_),
    .A(A[31]),
    .B(_196_));
 sg13g2_xor2_1 _523_ (.B(BI),
    .A(B[2]),
    .X(_198_));
 sg13g2_xnor2_1 _524_ (.Y(\Y[32:1] [30]),
    .A(_195_),
    .B(_197_));
 sg13g2_or2_1 _525_ (.X(_199_),
    .B(_197_),
    .A(_189_));
 sg13g2_nor3_1 _526_ (.A(_153_),
    .B(_179_),
    .C(_199_),
    .Y(_200_));
 sg13g2_nor2_1 _527_ (.A(_188_),
    .B(_197_),
    .Y(_201_));
 sg13g2_a21oi_1 _528_ (.A1(A[31]),
    .A2(_196_),
    .Y(_202_),
    .B1(_201_));
 sg13g2_o21ai_1 _529_ (.B1(_202_),
    .Y(_203_),
    .A1(_176_),
    .A2(_199_));
 sg13g2_nor2_1 _530_ (.A(_200_),
    .B(_203_),
    .Y(_204_));
 sg13g2_or3_1 _531_ (.A(_155_),
    .B(_179_),
    .C(_199_),
    .X(_205_));
 sg13g2_nand2_1 _532_ (.Y(_206_),
    .A(A[2]),
    .B(_198_));
 sg13g2_o21ai_1 _533_ (.B1(_204_),
    .Y(_207_),
    .A1(_115_),
    .A2(_205_));
 sg13g2_xor2_1 _534_ (.B(B[32]),
    .A(A[32]),
    .X(_208_));
 sg13g2_xnor2_1 _535_ (.Y(_209_),
    .A(BI),
    .B(_208_));
 sg13g2_xnor2_1 _536_ (.Y(\Y[32:1] [31]),
    .A(_207_),
    .B(_209_));
 sg13g2_xnor2_1 _537_ (.Y(_210_),
    .A(A[2]),
    .B(_198_));
 sg13g2_xnor2_1 _538_ (.Y(\Y[32:1] [1]),
    .A(_210_),
    .B(_186_));
 sg13g2_xor2_1 _539_ (.B(BI),
    .A(B[3]),
    .X(_211_));
 sg13g2_nand2_1 _540_ (.Y(_212_),
    .A(A[3]),
    .B(_211_));
 sg13g2_xnor2_1 _541_ (.Y(_213_),
    .A(A[3]),
    .B(_211_));
 sg13g2_o21ai_1 _542_ (.B1(_206_),
    .Y(_214_),
    .A1(_088_),
    .A2(_210_));
 sg13g2_nor3_1 _543_ (.A(_104_),
    .B(_161_),
    .C(_210_),
    .Y(_215_));
 sg13g2_or2_1 _544_ (.X(_216_),
    .B(_215_),
    .A(_214_));
 sg13g2_xnor2_1 _545_ (.Y(\Y[32:1] [2]),
    .A(_213_),
    .B(_216_));
 sg13g2_nor2_1 _546_ (.A(_210_),
    .B(_213_),
    .Y(_217_));
 sg13g2_o21ai_1 _547_ (.B1(_212_),
    .Y(_218_),
    .A1(_206_),
    .A2(_213_));
 sg13g2_a21o_1 _548_ (.A2(_217_),
    .A1(_186_),
    .B1(_218_),
    .X(_219_));
 sg13g2_xor2_1 _549_ (.B(BI),
    .A(B[4]),
    .X(_220_));
 sg13g2_nand2_1 _550_ (.Y(_221_),
    .A(A[4]),
    .B(_220_));
 sg13g2_xnor2_1 _551_ (.Y(_222_),
    .A(A[4]),
    .B(_220_));
 sg13g2_xnor2_1 _552_ (.Y(\Y[32:1] [3]),
    .A(_219_),
    .B(_222_));
 sg13g2_o21ai_1 _553_ (.B1(_221_),
    .Y(_223_),
    .A1(_212_),
    .A2(_222_));
 sg13g2_nor2_1 _554_ (.A(_213_),
    .B(_222_),
    .Y(_224_));
 sg13g2_nor4_1 _555_ (.A(_104_),
    .B(_210_),
    .C(_213_),
    .D(_222_),
    .Y(_225_));
 sg13g2_a221oi_1 _556_ (.B2(_163_),
    .C1(_223_),
    .B1(_225_),
    .A1(_214_),
    .Y(_226_),
    .A2(_224_));
 sg13g2_xor2_1 _557_ (.B(BI),
    .A(B[5]),
    .X(_227_));
 sg13g2_nand2_1 _558_ (.Y(_228_),
    .A(A[5]),
    .B(_227_));
 sg13g2_xnor2_1 _559_ (.Y(_229_),
    .A(A[5]),
    .B(_227_));
 sg13g2_xor2_1 _560_ (.B(_229_),
    .A(_226_),
    .X(\Y[32:1] [4]));
 sg13g2_xor2_1 _561_ (.B(BI),
    .A(B[6]),
    .X(_230_));
 sg13g2_nand2_1 _562_ (.Y(_231_),
    .A(A[6]),
    .B(_230_));
 sg13g2_xnor2_1 _563_ (.Y(_232_),
    .A(A[6]),
    .B(_230_));
 sg13g2_o21ai_1 _564_ (.B1(_228_),
    .Y(_233_),
    .A1(_221_),
    .A2(_229_));
 sg13g2_nor2_1 _565_ (.A(_222_),
    .B(_229_),
    .Y(_234_));
 sg13g2_nor4_1 _566_ (.A(_210_),
    .B(_213_),
    .C(_222_),
    .D(_229_),
    .Y(_235_));
 sg13g2_a221oi_1 _567_ (.B2(_186_),
    .C1(_233_),
    .B1(_235_),
    .A1(_218_),
    .Y(_236_),
    .A2(_234_));
 sg13g2_xor2_1 _568_ (.B(_236_),
    .A(_232_),
    .X(\Y[32:1] [5]));
 sg13g2_nor2_1 _569_ (.A(_229_),
    .B(_232_),
    .Y(_237_));
 sg13g2_and2_1 _570_ (.A(_224_),
    .B(_237_),
    .X(_238_));
 sg13g2_o21ai_1 _571_ (.B1(_231_),
    .Y(_239_),
    .A1(_228_),
    .A2(_232_));
 sg13g2_a21o_1 _572_ (.A2(_237_),
    .A1(_223_),
    .B1(_239_),
    .X(_240_));
 sg13g2_a21o_1 _573_ (.A2(_238_),
    .A1(_216_),
    .B1(_240_),
    .X(_241_));
 sg13g2_xor2_1 _574_ (.B(BI),
    .A(B[7]),
    .X(_242_));
 sg13g2_nand2_1 _575_ (.Y(_243_),
    .A(A[7]),
    .B(_242_));
 sg13g2_xnor2_1 _576_ (.Y(_244_),
    .A(A[7]),
    .B(_242_));
 sg13g2_xnor2_1 _577_ (.Y(\Y[32:1] [6]),
    .A(_241_),
    .B(_244_));
 sg13g2_nor2_1 _578_ (.A(_232_),
    .B(_244_),
    .Y(_245_));
 sg13g2_and2_1 _579_ (.A(_234_),
    .B(_245_),
    .X(_246_));
 sg13g2_o21ai_1 _580_ (.B1(_243_),
    .Y(_247_),
    .A1(_231_),
    .A2(_244_));
 sg13g2_a21o_1 _581_ (.A2(_245_),
    .A1(_233_),
    .B1(_247_),
    .X(_248_));
 sg13g2_a21o_1 _582_ (.A2(_246_),
    .A1(_219_),
    .B1(_248_),
    .X(_249_));
 sg13g2_xor2_1 _583_ (.B(BI),
    .A(B[8]),
    .X(_250_));
 sg13g2_nand2_1 _584_ (.Y(_251_),
    .A(A[8]),
    .B(_250_));
 sg13g2_xnor2_1 _585_ (.Y(_252_),
    .A(A[8]),
    .B(_250_));
 sg13g2_xnor2_1 _586_ (.Y(\Y[32:1] [7]),
    .A(_249_),
    .B(_252_));
 sg13g2_nor2_1 _587_ (.A(_244_),
    .B(_252_),
    .Y(_253_));
 sg13g2_o21ai_1 _588_ (.B1(_251_),
    .Y(_254_),
    .A1(_243_),
    .A2(_252_));
 sg13g2_a21oi_1 _589_ (.A1(_239_),
    .A2(_253_),
    .Y(_255_),
    .B1(_254_));
 sg13g2_nand2_1 _590_ (.Y(_256_),
    .A(_237_),
    .B(_253_));
 sg13g2_o21ai_1 _591_ (.B1(_255_),
    .Y(_257_),
    .A1(_226_),
    .A2(_256_));
 sg13g2_xor2_1 _592_ (.B(BI),
    .A(B[9]),
    .X(_258_));
 sg13g2_nand2_1 _593_ (.Y(_259_),
    .A(A[9]),
    .B(_258_));
 sg13g2_xnor2_1 _594_ (.Y(_260_),
    .A(A[9]),
    .B(_258_));
 sg13g2_xnor2_1 _595_ (.Y(\Y[32:1] [8]),
    .A(_257_),
    .B(_260_));
 sg13g2_nor2_1 _596_ (.A(_252_),
    .B(_260_),
    .Y(_261_));
 sg13g2_o21ai_1 _597_ (.B1(_259_),
    .Y(_262_),
    .A1(_251_),
    .A2(_260_));
 sg13g2_a21oi_1 _598_ (.A1(_247_),
    .A2(_261_),
    .Y(_263_),
    .B1(_262_));
 sg13g2_nand2_1 _599_ (.Y(_264_),
    .A(_245_),
    .B(_261_));
 sg13g2_o21ai_1 _600_ (.B1(_263_),
    .Y(_265_),
    .A1(_236_),
    .A2(_264_));
 sg13g2_xor2_1 _601_ (.B(BI),
    .A(B[10]),
    .X(_266_));
 sg13g2_nand2_1 _602_ (.Y(_267_),
    .A(A[10]),
    .B(_266_));
 sg13g2_xnor2_1 _603_ (.Y(_268_),
    .A(A[10]),
    .B(_266_));
 sg13g2_xnor2_1 _604_ (.Y(\Y[32:1] [9]),
    .A(_265_),
    .B(_268_));
 sg13g2_nor2_1 _605_ (.A(_260_),
    .B(_268_),
    .Y(_269_));
 sg13g2_o21ai_1 _606_ (.B1(_267_),
    .Y(_270_),
    .A1(_259_),
    .A2(_268_));
 sg13g2_a21o_1 _607_ (.A2(_269_),
    .A1(_254_),
    .B1(_270_),
    .X(_271_));
 sg13g2_nor4_1 _608_ (.A(_244_),
    .B(_252_),
    .C(_260_),
    .D(_268_),
    .Y(_272_));
 sg13g2_inv_1 _609_ (.Y(_273_),
    .A(_272_));
 sg13g2_and3_1 _610_ (.X(_274_),
    .A(_224_),
    .B(_237_),
    .C(_272_));
 sg13g2_a221oi_1 _611_ (.B2(_216_),
    .C1(_271_),
    .B1(_274_),
    .A1(_240_),
    .Y(_275_),
    .A2(_272_));
 sg13g2_xor2_1 _612_ (.B(BI),
    .A(B[11]),
    .X(_276_));
 sg13g2_nand2_1 _613_ (.Y(_277_),
    .A(A[11]),
    .B(_276_));
 sg13g2_xnor2_1 _614_ (.Y(_278_),
    .A(A[11]),
    .B(_276_));
 sg13g2_xor2_1 _615_ (.B(_278_),
    .A(_275_),
    .X(\Y[32:1] [10]));
 sg13g2_nor2_1 _616_ (.A(_268_),
    .B(_278_),
    .Y(_279_));
 sg13g2_o21ai_1 _617_ (.B1(_277_),
    .Y(_280_),
    .A1(_267_),
    .A2(_278_));
 sg13g2_a21o_1 _618_ (.A2(_279_),
    .A1(_262_),
    .B1(_280_),
    .X(_281_));
 sg13g2_nor4_1 _619_ (.A(_252_),
    .B(_260_),
    .C(_268_),
    .D(_278_),
    .Y(_282_));
 sg13g2_and3_1 _620_ (.X(_283_),
    .A(_234_),
    .B(_245_),
    .C(_282_));
 sg13g2_a221oi_1 _621_ (.B2(_219_),
    .C1(_281_),
    .B1(_283_),
    .A1(_248_),
    .Y(_284_),
    .A2(_282_));
 sg13g2_xor2_1 _622_ (.B(BI),
    .A(B[12]),
    .X(_285_));
 sg13g2_nand2_1 _623_ (.Y(_286_),
    .A(A[12]),
    .B(_285_));
 sg13g2_xnor2_1 _624_ (.Y(_287_),
    .A(A[12]),
    .B(_285_));
 sg13g2_xor2_1 _625_ (.B(_287_),
    .A(_284_),
    .X(\Y[32:1] [11]));
 sg13g2_xor2_1 _626_ (.B(BI),
    .A(B[13]),
    .X(_288_));
 sg13g2_nand2_1 _627_ (.Y(_289_),
    .A(A[13]),
    .B(_288_));
 sg13g2_xnor2_1 _628_ (.Y(_290_),
    .A(A[13]),
    .B(_288_));
 sg13g2_nor2_1 _629_ (.A(_278_),
    .B(_287_),
    .Y(_291_));
 sg13g2_o21ai_1 _630_ (.B1(_286_),
    .Y(_292_),
    .A1(_277_),
    .A2(_287_));
 sg13g2_a21oi_1 _631_ (.A1(_270_),
    .A2(_291_),
    .Y(_293_),
    .B1(_292_));
 sg13g2_nand2_1 _632_ (.Y(_294_),
    .A(_269_),
    .B(_291_));
 sg13g2_o21ai_1 _633_ (.B1(_293_),
    .Y(_295_),
    .A1(_255_),
    .A2(_294_));
 sg13g2_nor3_1 _634_ (.A(_226_),
    .B(_256_),
    .C(_294_),
    .Y(_296_));
 sg13g2_nor2_1 _635_ (.A(_295_),
    .B(_296_),
    .Y(_297_));
 sg13g2_xor2_1 _636_ (.B(_297_),
    .A(_290_),
    .X(\Y[32:1] [12]));
 sg13g2_xor2_1 _637_ (.B(BI),
    .A(B[14]),
    .X(_298_));
 sg13g2_nand2_1 _638_ (.Y(_299_),
    .A(A[14]),
    .B(_298_));
 sg13g2_xnor2_1 _639_ (.Y(_300_),
    .A(A[14]),
    .B(_298_));
 sg13g2_nor2_1 _640_ (.A(_287_),
    .B(_290_),
    .Y(_301_));
 sg13g2_o21ai_1 _641_ (.B1(_289_),
    .Y(_302_),
    .A1(_286_),
    .A2(_290_));
 sg13g2_a21oi_1 _642_ (.A1(_280_),
    .A2(_301_),
    .Y(_303_),
    .B1(_302_));
 sg13g2_nand2_1 _643_ (.Y(_304_),
    .A(_279_),
    .B(_301_));
 sg13g2_o21ai_1 _644_ (.B1(_303_),
    .Y(_305_),
    .A1(_263_),
    .A2(_304_));
 sg13g2_nor3_1 _645_ (.A(_236_),
    .B(_264_),
    .C(_304_),
    .Y(_306_));
 sg13g2_nor2_1 _646_ (.A(_305_),
    .B(_306_),
    .Y(_307_));
 sg13g2_xor2_1 _647_ (.B(_307_),
    .A(_300_),
    .X(\Y[32:1] [13]));
endmodule
module ALU_34_0_34_0_34_KOGGE_STONE (A,
    B,
    BI,
    CI,
    CO,
    X,
    Y);
 input [33:0] A;
 input [33:0] B;
 input BI;
 input CI;
 output [33:0] CO;
 output [33:0] X;
 output [33:0] Y;

 wire _267_;
 wire _265_;
 wire _264_;
 wire _263_;
 wire _260_;
 wire _257_;
 wire _255_;
 wire _254_;
 wire _253_;
 wire _252_;
 wire _251_;
 wire _250_;
 wire _249_;
 wire _248_;
 wire _247_;
 wire _246_;
 wire _245_;
 wire _244_;
 wire _242_;
 wire _241_;
 wire _240_;
 wire _239_;
 wire _238_;
 wire _237_;
 wire _236_;
 wire _235_;
 wire _234_;
 wire _232_;
 wire _231_;
 wire _230_;
 wire _229_;
 wire _228_;
 wire _226_;
 wire _225_;
 wire _224_;
 wire _223_;
 wire _222_;
 wire _221_;
 wire _220_;
 wire _219_;
 wire _218_;
 wire _216_;
 wire _215_;
 wire _214_;
 wire _213_;
 wire _212_;
 wire _210_;
 wire _209_;
 wire _208_;
 wire _207_;
 wire _206_;
 wire _205_;
 wire _204_;
 wire _203_;
 wire _202_;
 wire _200_;
 wire _199_;
 wire _198_;
 wire _197_;
 wire _196_;
 wire _195_;
 wire _194_;
 wire _193_;
 wire _191_;
 wire _190_;
 wire _189_;
 wire _188_;
 wire _187_;
 wire _186_;
 wire _184_;
 wire _183_;
 wire _182_;
 wire _181_;
 wire _180_;
 wire _179_;
 wire _178_;
 wire _176_;
 wire _175_;
 wire _174_;
 wire _172_;
 wire _171_;
 wire _170_;
 wire _169_;
 wire _167_;
 wire _166_;
 wire _165_;
 wire _164_;
 wire _266_;
 wire _256_;
 wire _227_;
 wire _217_;
 wire _211_;
 wire _201_;
 wire _162_;
 wire _185_;
 wire _177_;
 wire _161_;
 wire _173_;
 wire _168_;
 wire _163_;
 wire _160_;
 wire _159_;
 wire _158_;
 wire _157_;
 wire _156_;
 wire _155_;
 wire _154_;
 wire _153_;
 wire _152_;
 wire _151_;
 wire _150_;
 wire _149_;
 wire _148_;
 wire _147_;
 wire _146_;
 wire _145_;
 wire _144_;
 wire _143_;
 wire _142_;
 wire _141_;
 wire _140_;
 wire _139_;
 wire _138_;
 wire _137_;
 wire _136_;
 wire _135_;
 wire _134_;
 wire _133_;
 wire _132_;
 wire _131_;
 wire _130_;
 wire _129_;
 wire _128_;
 wire _127_;
 wire _126_;
 wire _125_;
 wire _124_;
 wire _123_;
 wire _122_;
 wire _121_;
 wire _120_;
 wire _119_;
 wire _118_;
 wire _117_;
 wire _116_;
 wire _115_;
 wire _114_;
 wire _113_;
 wire _112_;
 wire _111_;
 wire _110_;
 wire _109_;
 wire _108_;
 wire _107_;
 wire _106_;
 wire _105_;
 wire _104_;
 wire _103_;
 wire _102_;
 wire _101_;
 wire _100_;
 wire _099_;
 wire _098_;
 wire _097_;
 wire _096_;
 wire _095_;
 wire _094_;
 wire _093_;
 wire _092_;
 wire _091_;
 wire _090_;
 wire _089_;
 wire _088_;
 wire _087_;
 wire _086_;
 wire _085_;
 wire _084_;
 wire _083_;
 wire _082_;
 wire _081_;
 wire _080_;
 wire _079_;
 wire _078_;
 wire _077_;
 wire _076_;
 wire _075_;
 wire _074_;
 wire _073_;
 wire _072_;
 wire _071_;
 wire _070_;
 wire _284_;
 wire _069_;
 wire _068_;
 wire _067_;
 wire _066_;
 wire _065_;
 wire _064_;
 wire _063_;
 wire _062_;
 wire _061_;
 wire _273_;
 wire _060_;
 wire _059_;
 wire _058_;
 wire _057_;
 wire _056_;
 wire _055_;
 wire _054_;
 wire _053_;
 wire _052_;
 wire _051_;
 wire _050_;
 wire _259_;
 wire _192_;
 wire _049_;
 wire _262_;
 wire _048_;
 wire _047_;
 wire _046_;
 wire _045_;
 wire _044_;
 wire _043_;
 wire _042_;
 wire _041_;
 wire _040_;
 wire _039_;
 wire _291_;
 wire _038_;
 wire _290_;
 wire _037_;
 wire _036_;
 wire _035_;
 wire _034_;
 wire _033_;
 wire _032_;
 wire _031_;
 wire _030_;
 wire _243_;
 wire _281_;
 wire _029_;
 wire _028_;
 wire _027_;
 wire _280_;
 wire _026_;
 wire _025_;
 wire _024_;
 wire _023_;
 wire _022_;
 wire _021_;
 wire _020_;
 wire _233_;
 wire _268_;
 wire _019_;
 wire _018_;
 wire _272_;
 wire _017_;
 wire _288_;
 wire _289_;
 wire _016_;
 wire _015_;
 wire _014_;
 wire _013_;
 wire _012_;
 wire _011_;
 wire _010_;
 wire _009_;
 wire _258_;
 wire _261_;
 wire _008_;
 wire _007_;
 wire _006_;
 wire _278_;
 wire _005_;
 wire _279_;
 wire _004_;
 wire _003_;
 wire _287_;
 wire _286_;
 wire _002_;
 wire _001_;
 wire _000_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _282_;
 wire _283_;
 wire _285_;
 wire _292_;
 wire _293_;
 wire net6122;
 wire net6123;
 wire net6483;
 wire net6481;
 wire net6480;
 wire net6482;
 wire net6484;
 wire net6477;
 wire net6475;
 wire net6476;
 wire net6563;
 wire net6564;
 wire net6561;
 wire net6562;
 wire net6560;
 wire net6559;
 wire net6558;
 wire net6556;
 wire net6555;
 wire net6597;
 wire net6593;
 wire net6598;
 wire net6596;
 wire net6619;
 wire net6618;
 wire net5956;
 wire net6124;
 wire net6396;
 wire net6401;
 wire net6402;
 wire net6403;
 wire net6404;
 wire net6485;
 wire net6486;
 wire net6565;
 wire net6566;
 wire net6595;
 wire net6594;
 wire net6616;
 wire net6633;
 wire net6634;

 sg13g2_xor2_1 _294_ (.B(BI),
    .A(B[18]),
    .X(_000_));
 sg13g2_and2_1 _295_ (.A(A[18]),
    .B(_000_),
    .X(_001_));
 sg13g2_inv_1 _296_ (.Y(X[18]),
    .A(_002_));
 sg13g2_xnor2_1 _297_ (.Y(_002_),
    .A(A[18]),
    .B(_000_));
 sg13g2_nor3_1 _298_ (.A(_286_),
    .B(_287_),
    .C(_002_),
    .Y(_003_));
 sg13g2_a21o_1 _299_ (.A2(X[18]),
    .A1(_286_),
    .B1(_001_),
    .X(_004_));
 sg13g2_a21oi_1 _300_ (.A1(_279_),
    .A2(_003_),
    .Y(_005_),
    .B1(_004_));
 sg13g2_and2_1 _301_ (.A(_278_),
    .B(_003_),
    .X(_006_));
 sg13g2_inv_1 _302_ (.Y(_007_),
    .A(_006_));
 sg13g2_o21ai_1 _303_ (.B1(_005_),
    .Y(_008_),
    .A1(net6476),
    .A2(_007_));
 sg13g2_and2_1 _304_ (.A(_258_),
    .B(_006_),
    .X(_009_));
 sg13g2_a21o_1 _305_ (.A2(_009_),
    .A1(CO[10]),
    .B1(_008_),
    .X(CO[18]));
 sg13g2_xor2_1 _306_ (.B(BI),
    .A(B[19]),
    .X(_010_));
 sg13g2_and2_1 _307_ (.A(A[19]),
    .B(_010_),
    .X(_011_));
 sg13g2_nand2_1 _308_ (.Y(_012_),
    .A(A[19]),
    .B(_010_));
 sg13g2_inv_1 _309_ (.Y(X[19]),
    .A(_013_));
 sg13g2_xnor2_1 _310_ (.Y(_013_),
    .A(A[19]),
    .B(_010_));
 sg13g2_nand2b_1 _311_ (.Y(_014_),
    .B(X[19]),
    .A_N(net6566));
 sg13g2_a21oi_1 _312_ (.A1(_001_),
    .A2(X[19]),
    .Y(_015_),
    .B1(_011_));
 sg13g2_o21ai_1 _313_ (.B1(_015_),
    .Y(_016_),
    .A1(_289_),
    .A2(_014_));
 sg13g2_nor2_1 _314_ (.A(net6555),
    .B(_014_),
    .Y(_017_));
 sg13g2_a21oi_1 _315_ (.A1(_272_),
    .A2(_017_),
    .Y(_018_),
    .B1(_016_));
 sg13g2_nand2_1 _316_ (.Y(_019_),
    .A(_268_),
    .B(_017_));
 sg13g2_o21ai_1 _317_ (.B1(_018_),
    .Y(CO[19]),
    .A1(_233_),
    .A2(_019_));
 sg13g2_xor2_1 _318_ (.B(BI),
    .A(B[20]),
    .X(_020_));
 sg13g2_nand2_1 _319_ (.Y(_021_),
    .A(A[20]),
    .B(_020_));
 sg13g2_inv_1 _320_ (.Y(X[20]),
    .A(net6565));
 sg13g2_xnor2_1 _321_ (.Y(_022_),
    .A(A[20]),
    .B(_020_));
 sg13g2_nor2_1 _322_ (.A(_013_),
    .B(_022_),
    .Y(_023_));
 sg13g2_o21ai_1 _323_ (.B1(_021_),
    .Y(_024_),
    .A1(_012_),
    .A2(_022_));
 sg13g2_a21o_1 _324_ (.A2(_023_),
    .A1(_004_),
    .B1(_024_),
    .X(_025_));
 sg13g2_and2_1 _325_ (.A(_003_),
    .B(_023_),
    .X(_026_));
 sg13g2_nor2b_1 _326_ (.A(_280_),
    .B_N(_026_),
    .Y(_027_));
 sg13g2_nor2_1 _327_ (.A(_025_),
    .B(_027_),
    .Y(_028_));
 sg13g2_nand2b_1 _328_ (.Y(_029_),
    .B(_026_),
    .A_N(_281_));
 sg13g2_o21ai_1 _329_ (.B1(_028_),
    .Y(CO[20]),
    .A1(_243_),
    .A2(_029_));
 sg13g2_xor2_1 _330_ (.B(BI),
    .A(B[21]),
    .X(_030_));
 sg13g2_nand2_1 _331_ (.Y(_031_),
    .A(A[21]),
    .B(_030_));
 sg13g2_inv_1 _332_ (.Y(X[21]),
    .A(_032_));
 sg13g2_xnor2_1 _333_ (.Y(_032_),
    .A(A[21]),
    .B(_030_));
 sg13g2_nand2b_1 _334_ (.Y(_033_),
    .B(X[21]),
    .A_N(net6565));
 sg13g2_nor2_1 _335_ (.A(_021_),
    .B(_032_),
    .Y(_034_));
 sg13g2_a21oi_1 _336_ (.A1(A[21]),
    .A2(_030_),
    .Y(_035_),
    .B1(_034_));
 sg13g2_o21ai_1 _337_ (.B1(_035_),
    .Y(_036_),
    .A1(_015_),
    .A2(_033_));
 sg13g2_nor2_1 _338_ (.A(_014_),
    .B(_033_),
    .Y(_037_));
 sg13g2_a21o_1 _339_ (.A2(_037_),
    .A1(_290_),
    .B1(_036_),
    .X(_038_));
 sg13g2_and2_1 _340_ (.A(net6475),
    .B(_037_),
    .X(_039_));
 sg13g2_a21o_1 _341_ (.A2(_039_),
    .A1(CO[13]),
    .B1(_038_),
    .X(CO[21]));
 sg13g2_xor2_1 _342_ (.B(BI),
    .A(B[22]),
    .X(_040_));
 sg13g2_nand2_1 _343_ (.Y(_041_),
    .A(A[22]),
    .B(_040_));
 sg13g2_inv_1 _344_ (.Y(X[22]),
    .A(net6563));
 sg13g2_xnor2_1 _345_ (.Y(_042_),
    .A(A[22]),
    .B(_040_));
 sg13g2_nor2_1 _346_ (.A(_032_),
    .B(_042_),
    .Y(_043_));
 sg13g2_o21ai_1 _347_ (.B1(_041_),
    .Y(_044_),
    .A1(_031_),
    .A2(_042_));
 sg13g2_a21oi_1 _348_ (.A1(_024_),
    .A2(_043_),
    .Y(_045_),
    .B1(_044_));
 sg13g2_and2_1 _349_ (.A(_023_),
    .B(_043_),
    .X(_046_));
 sg13g2_nand2b_1 _350_ (.Y(_047_),
    .B(_046_),
    .A_N(_005_));
 sg13g2_nand2_1 _351_ (.Y(_048_),
    .A(_006_),
    .B(_046_));
 sg13g2_a21o_1 _352_ (.A2(net6396),
    .A1(net6476),
    .B1(_048_),
    .X(_049_));
 sg13g2_or3_1 _353_ (.A(net6597),
    .B(_259_),
    .C(_048_),
    .X(_050_));
 sg13g2_nand4_1 _354_ (.B(_047_),
    .C(_049_),
    .A(_045_),
    .Y(CO[22]),
    .D(_050_));
 sg13g2_xor2_1 _355_ (.B(BI),
    .A(B[23]),
    .X(_051_));
 sg13g2_nand2_1 _356_ (.Y(_052_),
    .A(A[23]),
    .B(_051_));
 sg13g2_inv_1 _357_ (.Y(X[23]),
    .A(net6562));
 sg13g2_xnor2_1 _358_ (.Y(_053_),
    .A(A[23]),
    .B(_051_));
 sg13g2_or2_1 _359_ (.X(_054_),
    .B(_053_),
    .A(_042_));
 sg13g2_nor2_1 _360_ (.A(_035_),
    .B(_054_),
    .Y(_055_));
 sg13g2_o21ai_1 _361_ (.B1(_052_),
    .Y(_056_),
    .A1(_041_),
    .A2(_053_));
 sg13g2_nor2_1 _362_ (.A(_033_),
    .B(_054_),
    .Y(_057_));
 sg13g2_and2_1 _363_ (.A(_016_),
    .B(_057_),
    .X(_058_));
 sg13g2_nor3_1 _364_ (.A(_055_),
    .B(_056_),
    .C(_058_),
    .Y(_059_));
 sg13g2_nand2_1 _365_ (.Y(_060_),
    .A(_017_),
    .B(net6124));
 sg13g2_o21ai_1 _366_ (.B1(_059_),
    .Y(CO[23]),
    .A1(net6123),
    .A2(_060_));
 sg13g2_xor2_1 _367_ (.B(BI),
    .A(B[24]),
    .X(_061_));
 sg13g2_nand2_1 _368_ (.Y(_062_),
    .A(A[24]),
    .B(_061_));
 sg13g2_inv_1 _369_ (.Y(X[24]),
    .A(net6561));
 sg13g2_xnor2_1 _370_ (.Y(_063_),
    .A(A[24]),
    .B(_061_));
 sg13g2_nor2_1 _371_ (.A(_053_),
    .B(_063_),
    .Y(_064_));
 sg13g2_o21ai_1 _372_ (.B1(_062_),
    .Y(_065_),
    .A1(_052_),
    .A2(_063_));
 sg13g2_a21o_1 _373_ (.A2(_064_),
    .A1(_044_),
    .B1(_065_),
    .X(_066_));
 sg13g2_and2_1 _374_ (.A(_043_),
    .B(_064_),
    .X(_067_));
 sg13g2_a21oi_1 _375_ (.A1(_025_),
    .A2(_067_),
    .Y(_068_),
    .B1(_066_));
 sg13g2_nand3b_1 _376_ (.B(net6404),
    .C(_067_),
    .Y(_069_),
    .A_N(net6122));
 sg13g2_nand2_1 _377_ (.Y(CO[24]),
    .A(_068_),
    .B(_069_));
 sg13g2_xor2_1 _378_ (.B(BI),
    .A(B[25]),
    .X(_070_));
 sg13g2_nand2_1 _379_ (.Y(_071_),
    .A(A[25]),
    .B(_070_));
 sg13g2_inv_1 _380_ (.Y(X[25]),
    .A(net6560));
 sg13g2_xnor2_1 _381_ (.Y(_072_),
    .A(A[25]),
    .B(_070_));
 sg13g2_nor2_1 _382_ (.A(_063_),
    .B(_072_),
    .Y(_073_));
 sg13g2_o21ai_1 _383_ (.B1(_071_),
    .Y(_074_),
    .A1(_062_),
    .A2(_072_));
 sg13g2_a21oi_1 _384_ (.A1(_056_),
    .A2(_073_),
    .Y(_075_),
    .B1(_074_));
 sg13g2_nor2b_1 _385_ (.A(_054_),
    .B_N(_073_),
    .Y(_076_));
 sg13g2_nand2_1 _386_ (.Y(_077_),
    .A(_036_),
    .B(_076_));
 sg13g2_nand3_1 _387_ (.B(_037_),
    .C(_076_),
    .A(CO[17]),
    .Y(_078_));
 sg13g2_and3_1 _388_ (.X(_079_),
    .A(_075_),
    .B(_077_),
    .C(_078_));
 sg13g2_inv_1 _389_ (.Y(CO[25]),
    .A(net5956));
 sg13g2_xor2_1 _390_ (.B(BI),
    .A(B[26]),
    .X(_080_));
 sg13g2_nand2_1 _391_ (.Y(_081_),
    .A(A[26]),
    .B(_080_));
 sg13g2_inv_1 _392_ (.Y(X[26]),
    .A(_082_));
 sg13g2_xnor2_1 _393_ (.Y(_082_),
    .A(A[26]),
    .B(_080_));
 sg13g2_nor2_1 _394_ (.A(_072_),
    .B(_082_),
    .Y(_083_));
 sg13g2_o21ai_1 _395_ (.B1(_081_),
    .Y(_084_),
    .A1(_071_),
    .A2(_082_));
 sg13g2_a21oi_1 _396_ (.A1(_065_),
    .A2(net6485),
    .Y(_085_),
    .B1(_084_));
 sg13g2_nand2_1 _397_ (.Y(_086_),
    .A(net6486),
    .B(net6485));
 sg13g2_xor2_1 _398_ (.B(BI),
    .A(B[0]),
    .X(_087_));
 sg13g2_o21ai_1 _399_ (.B1(_085_),
    .Y(_088_),
    .A1(_045_),
    .A2(_086_));
 sg13g2_and3_1 _400_ (.X(_089_),
    .A(_046_),
    .B(net6486),
    .C(net6485));
 sg13g2_a21o_1 _401_ (.A2(_089_),
    .A1(CO[18]),
    .B1(_088_),
    .X(CO[26]));
 sg13g2_and2_1 _402_ (.A(A[0]),
    .B(_087_),
    .X(_090_));
 sg13g2_xor2_1 _403_ (.B(BI),
    .A(B[27]),
    .X(_091_));
 sg13g2_nand2_1 _404_ (.Y(_092_),
    .A(net6593),
    .B(_091_));
 sg13g2_inv_1 _405_ (.Y(X[27]),
    .A(net6559));
 sg13g2_xnor2_1 _406_ (.Y(_093_),
    .A(net6593),
    .B(_091_));
 sg13g2_nor2_1 _407_ (.A(_082_),
    .B(net6559),
    .Y(_094_));
 sg13g2_o21ai_1 _408_ (.B1(_092_),
    .Y(_095_),
    .A1(_081_),
    .A2(net6559));
 sg13g2_a21oi_1 _409_ (.A1(_074_),
    .A2(_094_),
    .Y(_096_),
    .B1(_095_));
 sg13g2_and2_1 _410_ (.A(_073_),
    .B(_094_),
    .X(_097_));
 sg13g2_o21ai_1 _411_ (.B1(_097_),
    .Y(_098_),
    .A1(_055_),
    .A2(_056_));
 sg13g2_nand2_1 _412_ (.Y(_099_),
    .A(_096_),
    .B(_098_));
 sg13g2_and2_1 _413_ (.A(net6124),
    .B(_097_),
    .X(_100_));
 sg13g2_a21o_1 _414_ (.A2(_100_),
    .A1(CO[19]),
    .B1(_099_),
    .X(CO[27]));
 sg13g2_xor2_1 _415_ (.B(BI),
    .A(net6616),
    .X(_101_));
 sg13g2_nand2_1 _416_ (.Y(_102_),
    .A(A[28]),
    .B(net6598));
 sg13g2_inv_1 _417_ (.Y(X[28]),
    .A(net6558));
 sg13g2_xnor2_1 _418_ (.Y(_103_),
    .A(A[28]),
    .B(_101_));
 sg13g2_nor2_1 _419_ (.A(_093_),
    .B(_103_),
    .Y(_104_));
 sg13g2_o21ai_1 _420_ (.B1(_102_),
    .Y(_105_),
    .A1(_092_),
    .A2(_103_));
 sg13g2_a21o_1 _421_ (.A2(_104_),
    .A1(_084_),
    .B1(_105_),
    .X(_106_));
 sg13g2_and2_1 _422_ (.A(_083_),
    .B(_104_),
    .X(_107_));
 sg13g2_xor2_1 _423_ (.B(_087_),
    .A(A[0]),
    .X(X[0]));
 sg13g2_a21o_1 _424_ (.A2(_107_),
    .A1(_066_),
    .B1(_106_),
    .X(_108_));
 sg13g2_and2_1 _425_ (.A(_067_),
    .B(_107_),
    .X(_109_));
 sg13g2_a21o_1 _426_ (.A2(_109_),
    .A1(CO[20]),
    .B1(_108_),
    .X(CO[28]));
 sg13g2_xor2_1 _427_ (.B(BI),
    .A(B[29]),
    .X(_110_));
 sg13g2_nand2_1 _428_ (.Y(_111_),
    .A(A[29]),
    .B(_110_));
 sg13g2_a21oi_1 _429_ (.A1(CI),
    .A2(X[0]),
    .Y(_112_),
    .B1(_090_));
 sg13g2_inv_1 _430_ (.Y(X[29]),
    .A(_113_));
 sg13g2_xnor2_1 _431_ (.Y(_113_),
    .A(A[29]),
    .B(_110_));
 sg13g2_nor2_1 _432_ (.A(net6558),
    .B(_113_),
    .Y(_114_));
 sg13g2_inv_1 _433_ (.Y(CO[0]),
    .A(_112_));
 sg13g2_o21ai_1 _434_ (.B1(_111_),
    .Y(_115_),
    .A1(_102_),
    .A2(_113_));
 sg13g2_a21oi_1 _435_ (.A1(_095_),
    .A2(_114_),
    .Y(_116_),
    .B1(_115_));
 sg13g2_and2_1 _436_ (.A(_094_),
    .B(_114_),
    .X(_117_));
 sg13g2_inv_1 _437_ (.Y(_118_),
    .A(_117_));
 sg13g2_o21ai_1 _438_ (.B1(_116_),
    .Y(_119_),
    .A1(_075_),
    .A2(_118_));
 sg13g2_and2_1 _439_ (.A(net6403),
    .B(_117_),
    .X(_120_));
 sg13g2_a21o_1 _440_ (.A2(_120_),
    .A1(CO[21]),
    .B1(_119_),
    .X(CO[29]));
 sg13g2_xor2_1 _441_ (.B(BI),
    .A(B[30]),
    .X(_121_));
 sg13g2_nand2_1 _442_ (.Y(_122_),
    .A(A[30]),
    .B(_121_));
 sg13g2_inv_1 _443_ (.Y(X[30]),
    .A(net6480));
 sg13g2_xnor2_1 _444_ (.Y(_123_),
    .A(A[30]),
    .B(_121_));
 sg13g2_o21ai_1 _445_ (.B1(_122_),
    .Y(_124_),
    .A1(_111_),
    .A2(_123_));
 sg13g2_nor2_1 _446_ (.A(_113_),
    .B(_123_),
    .Y(_125_));
 sg13g2_nand2_1 _447_ (.Y(_126_),
    .A(net6483),
    .B(_125_));
 sg13g2_a21oi_1 _448_ (.A1(net6482),
    .A2(_125_),
    .Y(_127_),
    .B1(_124_));
 sg13g2_o21ai_1 _449_ (.B1(_127_),
    .Y(_128_),
    .A1(_085_),
    .A2(_126_));
 sg13g2_and4_1 _450_ (.A(net6486),
    .B(net6485),
    .C(net6484),
    .D(_125_),
    .X(_129_));
 sg13g2_a21o_1 _451_ (.A2(_129_),
    .A1(CO[22]),
    .B1(_128_),
    .X(CO[30]));
 sg13g2_xor2_1 _452_ (.B(BI),
    .A(B[1]),
    .X(_130_));
 sg13g2_xor2_1 _453_ (.B(BI),
    .A(B[31]),
    .X(_131_));
 sg13g2_nand2_1 _454_ (.Y(_132_),
    .A(A[31]),
    .B(_131_));
 sg13g2_inv_1 _455_ (.Y(X[31]),
    .A(_133_));
 sg13g2_xnor2_1 _456_ (.Y(_133_),
    .A(A[31]),
    .B(_131_));
 sg13g2_nor2_1 _457_ (.A(net6480),
    .B(_133_),
    .Y(_134_));
 sg13g2_nand3_1 _458_ (.B(net6481),
    .C(_134_),
    .A(_097_),
    .Y(_135_));
 sg13g2_nor2_1 _459_ (.A(_060_),
    .B(_135_),
    .Y(_136_));
 sg13g2_nand3b_1 _460_ (.B(net6481),
    .C(_134_),
    .Y(_137_),
    .A_N(_096_));
 sg13g2_nand2_1 _461_ (.Y(_138_),
    .A(A[1]),
    .B(_130_));
 sg13g2_o21ai_1 _462_ (.B1(_132_),
    .Y(_139_),
    .A1(_122_),
    .A2(_133_));
 sg13g2_a21oi_1 _463_ (.A1(_115_),
    .A2(_134_),
    .Y(_140_),
    .B1(_139_));
 sg13g2_and2_1 _464_ (.A(_137_),
    .B(_140_),
    .X(_141_));
 sg13g2_o21ai_1 _465_ (.B1(_141_),
    .Y(_142_),
    .A1(_059_),
    .A2(_135_));
 sg13g2_a21o_1 _466_ (.A2(_136_),
    .A1(CO[15]),
    .B1(_142_),
    .X(CO[31]));
 sg13g2_xor2_1 _467_ (.B(BI),
    .A(B[32]),
    .X(_143_));
 sg13g2_nand2_1 _468_ (.Y(_144_),
    .A(A[32]),
    .B(_143_));
 sg13g2_inv_1 _469_ (.Y(X[32]),
    .A(_145_));
 sg13g2_xnor2_1 _470_ (.Y(_145_),
    .A(A[32]),
    .B(_143_));
 sg13g2_nor2_1 _471_ (.A(_133_),
    .B(_145_),
    .Y(_146_));
 sg13g2_and2_1 _472_ (.A(_125_),
    .B(_146_),
    .X(_147_));
 sg13g2_o21ai_1 _473_ (.B1(_144_),
    .Y(_148_),
    .A1(_132_),
    .A2(_145_));
 sg13g2_a221oi_1 _474_ (.B2(net6402),
    .C1(_148_),
    .B1(_147_),
    .A1(_124_),
    .Y(_149_),
    .A2(_146_));
 sg13g2_nand2_1 _475_ (.Y(_150_),
    .A(net6401),
    .B(_147_));
 sg13g2_and2_1 _476_ (.A(_068_),
    .B(_149_),
    .X(_151_));
 sg13g2_inv_1 _477_ (.Y(X[1]),
    .A(_152_));
 sg13g2_xnor2_1 _478_ (.Y(_152_),
    .A(A[1]),
    .B(_130_));
 sg13g2_a22oi_1 _479_ (.Y(CO[32]),
    .B1(_151_),
    .B2(_069_),
    .A2(_150_),
    .A1(_149_));
 sg13g2_xor2_1 _480_ (.B(BI),
    .A(B[33]),
    .X(_153_));
 sg13g2_inv_1 _481_ (.Y(X[33]),
    .A(_154_));
 sg13g2_xnor2_1 _482_ (.Y(_154_),
    .A(A[33]),
    .B(_153_));
 sg13g2_nor2_1 _483_ (.A(_144_),
    .B(_154_),
    .Y(_155_));
 sg13g2_o21ai_1 _484_ (.B1(_138_),
    .Y(CO[1]),
    .A1(_112_),
    .A2(_152_));
 sg13g2_nor2_1 _485_ (.A(_145_),
    .B(_154_),
    .Y(_156_));
 sg13g2_nand2b_1 _486_ (.Y(_157_),
    .B(_134_),
    .A_N(_116_));
 sg13g2_nand2b_1 _487_ (.Y(_158_),
    .B(_157_),
    .A_N(_139_));
 sg13g2_a221oi_1 _488_ (.B2(_158_),
    .C1(_155_),
    .B1(_156_),
    .A1(A[33]),
    .Y(_159_),
    .A2(_153_));
 sg13g2_nand3_1 _489_ (.B(_134_),
    .C(_156_),
    .A(_117_),
    .Y(_160_));
 sg13g2_o21ai_1 _490_ (.B1(_159_),
    .Y(CO[33]),
    .A1(net5956),
    .A2(_160_));
 sg13g2_xor2_1 _491_ (.B(X[0]),
    .A(CI),
    .X(Y[0]));
 sg13g2_xnor2_1 _492_ (.Y(Y[1]),
    .A(_112_),
    .B(X[1]));
 sg13g2_xnor2_1 _493_ (.Y(Y[2]),
    .A(CO[1]),
    .B(_163_));
 sg13g2_xnor2_1 _494_ (.Y(Y[3]),
    .A(CO[2]),
    .B(_168_));
 sg13g2_xnor2_1 _495_ (.Y(Y[4]),
    .A(CO[3]),
    .B(_173_));
 sg13g2_xor2_1 _496_ (.B(BI),
    .A(B[2]),
    .X(_161_));
 sg13g2_xnor2_1 _497_ (.Y(Y[5]),
    .A(_177_),
    .B(X[5]));
 sg13g2_xnor2_1 _498_ (.Y(Y[6]),
    .A(_185_),
    .B(X[6]));
 sg13g2_nand2_1 _499_ (.Y(_162_),
    .A(A[2]),
    .B(_161_));
 sg13g2_xnor2_1 _500_ (.Y(Y[7]),
    .A(net6597),
    .B(X[7]));
 sg13g2_xnor2_1 _501_ (.Y(Y[8]),
    .A(_201_),
    .B(X[8]));
 sg13g2_xnor2_1 _502_ (.Y(Y[9]),
    .A(CO[8]),
    .B(_211_));
 sg13g2_xnor2_1 _503_ (.Y(Y[10]),
    .A(_217_),
    .B(X[10]));
 sg13g2_xnor2_1 _504_ (.Y(Y[11]),
    .A(CO[10]),
    .B(net6619));
 sg13g2_xnor2_1 _505_ (.Y(Y[12]),
    .A(_233_),
    .B(X[12]));
 sg13g2_xnor2_1 _506_ (.Y(Y[13]),
    .A(_243_),
    .B(X[13]));
 sg13g2_xnor2_1 _507_ (.Y(Y[14]),
    .A(CO[13]),
    .B(net6596));
 sg13g2_inv_1 _508_ (.Y(X[2]),
    .A(_163_));
 sg13g2_xnor2_1 _509_ (.Y(_163_),
    .A(A[2]),
    .B(_161_));
 sg13g2_xnor2_1 _510_ (.Y(Y[15]),
    .A(CO[14]),
    .B(net6595));
 sg13g2_nor2_1 _511_ (.A(_152_),
    .B(_163_),
    .Y(_164_));
 sg13g2_xnor2_1 _512_ (.Y(Y[16]),
    .A(_273_),
    .B(X[16]));
 sg13g2_xnor2_1 _513_ (.Y(Y[17]),
    .A(_284_),
    .B(X[17]));
 sg13g2_xnor2_1 _514_ (.Y(Y[18]),
    .A(CO[17]),
    .B(net6566));
 sg13g2_xnor2_1 _515_ (.Y(Y[19]),
    .A(CO[18]),
    .B(_013_));
 sg13g2_xnor2_1 _516_ (.Y(Y[20]),
    .A(CO[19]),
    .B(net6565));
 sg13g2_xnor2_1 _517_ (.Y(Y[21]),
    .A(CO[20]),
    .B(net6564));
 sg13g2_xnor2_1 _518_ (.Y(Y[22]),
    .A(CO[21]),
    .B(net6563));
 sg13g2_xnor2_1 _519_ (.Y(Y[23]),
    .A(CO[22]),
    .B(net6562));
 sg13g2_xnor2_1 _520_ (.Y(Y[24]),
    .A(CO[23]),
    .B(net6561));
 sg13g2_o21ai_1 _521_ (.B1(_162_),
    .Y(_165_),
    .A1(_138_),
    .A2(_163_));
 sg13g2_xnor2_1 _522_ (.Y(Y[25]),
    .A(CO[24]),
    .B(net6560));
 sg13g2_xnor2_1 _523_ (.Y(Y[26]),
    .A(_079_),
    .B(X[26]));
 sg13g2_a21o_1 _524_ (.A2(_164_),
    .A1(CO[0]),
    .B1(_165_),
    .X(CO[2]));
 sg13g2_xnor2_1 _525_ (.Y(Y[27]),
    .A(CO[26]),
    .B(net6559));
 sg13g2_xnor2_1 _526_ (.Y(Y[28]),
    .A(CO[27]),
    .B(net6558));
 sg13g2_xnor2_1 _527_ (.Y(Y[29]),
    .A(CO[28]),
    .B(_113_));
 sg13g2_xnor2_1 _528_ (.Y(Y[30]),
    .A(CO[29]),
    .B(net6480));
 sg13g2_xnor2_1 _529_ (.Y(Y[31]),
    .A(CO[30]),
    .B(_133_));
 sg13g2_xnor2_1 _530_ (.Y(Y[32]),
    .A(CO[31]),
    .B(_145_));
 sg13g2_xnor2_1 _531_ (.Y(Y[33]),
    .A(CO[32]),
    .B(_154_));
 sg13g2_xor2_1 _532_ (.B(BI),
    .A(B[3]),
    .X(_166_));
 sg13g2_nand2_1 _533_ (.Y(_167_),
    .A(A[3]),
    .B(_166_));
 sg13g2_inv_1 _534_ (.Y(X[3]),
    .A(_168_));
 sg13g2_xnor2_1 _535_ (.Y(_168_),
    .A(A[3]),
    .B(_166_));
 sg13g2_nor2_1 _536_ (.A(_163_),
    .B(_168_),
    .Y(_169_));
 sg13g2_o21ai_1 _537_ (.B1(_167_),
    .Y(_170_),
    .A1(_162_),
    .A2(_168_));
 sg13g2_a21o_1 _538_ (.A2(_169_),
    .A1(CO[1]),
    .B1(_170_),
    .X(CO[3]));
 sg13g2_xor2_1 _539_ (.B(BI),
    .A(B[4]),
    .X(_171_));
 sg13g2_nand2_1 _540_ (.Y(_172_),
    .A(A[4]),
    .B(_171_));
 sg13g2_inv_1 _541_ (.Y(X[4]),
    .A(_173_));
 sg13g2_xnor2_1 _542_ (.Y(_173_),
    .A(A[4]),
    .B(_171_));
 sg13g2_o21ai_1 _543_ (.B1(_172_),
    .Y(_174_),
    .A1(_167_),
    .A2(_173_));
 sg13g2_nor2_1 _544_ (.A(_168_),
    .B(_173_),
    .Y(_175_));
 sg13g2_nor4_1 _545_ (.A(_152_),
    .B(_163_),
    .C(_168_),
    .D(_173_),
    .Y(_176_));
 sg13g2_inv_1 _546_ (.Y(CO[4]),
    .A(_177_));
 sg13g2_a221oi_1 _547_ (.B2(CO[0]),
    .C1(_174_),
    .B1(_176_),
    .A1(_165_),
    .Y(_177_),
    .A2(_175_));
 sg13g2_xor2_1 _548_ (.B(BI),
    .A(B[5]),
    .X(_178_));
 sg13g2_nand2_1 _549_ (.Y(_179_),
    .A(A[5]),
    .B(_178_));
 sg13g2_inv_1 _550_ (.Y(X[5]),
    .A(_180_));
 sg13g2_xnor2_1 _551_ (.Y(_180_),
    .A(A[5]),
    .B(_178_));
 sg13g2_nor2_1 _552_ (.A(_173_),
    .B(_180_),
    .Y(_181_));
 sg13g2_nor4_1 _553_ (.A(_163_),
    .B(_168_),
    .C(_173_),
    .D(_180_),
    .Y(_182_));
 sg13g2_o21ai_1 _554_ (.B1(_179_),
    .Y(_183_),
    .A1(_172_),
    .A2(_180_));
 sg13g2_a21o_1 _555_ (.A2(_181_),
    .A1(_170_),
    .B1(_183_),
    .X(_184_));
 sg13g2_a21oi_1 _556_ (.A1(CO[1]),
    .A2(_182_),
    .Y(_185_),
    .B1(_184_));
 sg13g2_inv_1 _557_ (.Y(CO[5]),
    .A(_185_));
 sg13g2_xor2_1 _558_ (.B(BI),
    .A(B[6]),
    .X(_186_));
 sg13g2_nand2_1 _559_ (.Y(_187_),
    .A(A[6]),
    .B(_186_));
 sg13g2_inv_1 _560_ (.Y(X[6]),
    .A(_188_));
 sg13g2_xnor2_1 _561_ (.Y(_188_),
    .A(A[6]),
    .B(_186_));
 sg13g2_nor2_1 _562_ (.A(_180_),
    .B(_188_),
    .Y(_189_));
 sg13g2_and2_1 _563_ (.A(_175_),
    .B(_189_),
    .X(_190_));
 sg13g2_o21ai_1 _564_ (.B1(_187_),
    .Y(_191_),
    .A1(_179_),
    .A2(_188_));
 sg13g2_a221oi_1 _565_ (.B2(CO[2]),
    .C1(_191_),
    .B1(_190_),
    .A1(_174_),
    .Y(_192_),
    .A2(_189_));
 sg13g2_inv_1 _566_ (.Y(CO[6]),
    .A(net6597));
 sg13g2_xor2_1 _567_ (.B(BI),
    .A(B[7]),
    .X(_193_));
 sg13g2_nand2_1 _568_ (.Y(_194_),
    .A(A[7]),
    .B(_193_));
 sg13g2_inv_1 _569_ (.Y(X[7]),
    .A(_195_));
 sg13g2_xnor2_1 _570_ (.Y(_195_),
    .A(A[7]),
    .B(_193_));
 sg13g2_nor2_1 _571_ (.A(_188_),
    .B(_195_),
    .Y(_196_));
 sg13g2_o21ai_1 _572_ (.B1(_194_),
    .Y(_197_),
    .A1(_187_),
    .A2(_195_));
 sg13g2_a21o_1 _573_ (.A2(_196_),
    .A1(_183_),
    .B1(_197_),
    .X(_198_));
 sg13g2_inv_1 _574_ (.Y(_199_),
    .A(_200_));
 sg13g2_nand2_1 _575_ (.Y(_200_),
    .A(_181_),
    .B(_196_));
 sg13g2_a21oi_1 _576_ (.A1(CO[3]),
    .A2(_199_),
    .Y(_201_),
    .B1(_198_));
 sg13g2_inv_1 _577_ (.Y(CO[7]),
    .A(_201_));
 sg13g2_xor2_1 _578_ (.B(BI),
    .A(B[8]),
    .X(_202_));
 sg13g2_nand2_1 _579_ (.Y(_203_),
    .A(A[8]),
    .B(_202_));
 sg13g2_inv_1 _580_ (.Y(X[8]),
    .A(_204_));
 sg13g2_xnor2_1 _581_ (.Y(_204_),
    .A(A[8]),
    .B(_202_));
 sg13g2_nor2_1 _582_ (.A(_195_),
    .B(_204_),
    .Y(_205_));
 sg13g2_o21ai_1 _583_ (.B1(_203_),
    .Y(_206_),
    .A1(_194_),
    .A2(_204_));
 sg13g2_a21oi_1 _584_ (.A1(_191_),
    .A2(_205_),
    .Y(_207_),
    .B1(_206_));
 sg13g2_nand2_1 _585_ (.Y(_208_),
    .A(_189_),
    .B(_205_));
 sg13g2_o21ai_1 _586_ (.B1(_207_),
    .Y(CO[8]),
    .A1(_177_),
    .A2(_208_));
 sg13g2_xor2_1 _587_ (.B(BI),
    .A(B[9]),
    .X(_209_));
 sg13g2_nand2_1 _588_ (.Y(_210_),
    .A(A[9]),
    .B(_209_));
 sg13g2_inv_1 _589_ (.Y(X[9]),
    .A(_211_));
 sg13g2_xnor2_1 _590_ (.Y(_211_),
    .A(A[9]),
    .B(_209_));
 sg13g2_nor2_1 _591_ (.A(_204_),
    .B(_211_),
    .Y(_212_));
 sg13g2_o21ai_1 _592_ (.B1(_210_),
    .Y(_213_),
    .A1(_203_),
    .A2(_211_));
 sg13g2_a21o_1 _593_ (.A2(_212_),
    .A1(_197_),
    .B1(_213_),
    .X(_214_));
 sg13g2_nor4_1 _594_ (.A(_188_),
    .B(_195_),
    .C(_204_),
    .D(_211_),
    .Y(_215_));
 sg13g2_and2_1 _595_ (.A(_182_),
    .B(_215_),
    .X(_216_));
 sg13g2_a221oi_1 _596_ (.B2(CO[1]),
    .C1(_214_),
    .B1(_216_),
    .A1(_184_),
    .Y(_217_),
    .A2(_215_));
 sg13g2_inv_1 _597_ (.Y(CO[9]),
    .A(_217_));
 sg13g2_xor2_1 _598_ (.B(BI),
    .A(B[10]),
    .X(_218_));
 sg13g2_nand2_1 _599_ (.Y(_219_),
    .A(A[10]),
    .B(_218_));
 sg13g2_inv_1 _600_ (.Y(X[10]),
    .A(_220_));
 sg13g2_xnor2_1 _601_ (.Y(_220_),
    .A(A[10]),
    .B(_218_));
 sg13g2_nor2_1 _602_ (.A(_211_),
    .B(_220_),
    .Y(_221_));
 sg13g2_o21ai_1 _603_ (.B1(_219_),
    .Y(_222_),
    .A1(_210_),
    .A2(_220_));
 sg13g2_a21oi_1 _604_ (.A1(_206_),
    .A2(_221_),
    .Y(_223_),
    .B1(_222_));
 sg13g2_nand2_1 _605_ (.Y(_224_),
    .A(_205_),
    .B(_221_));
 sg13g2_o21ai_1 _606_ (.B1(_223_),
    .Y(CO[10]),
    .A1(net6597),
    .A2(_224_));
 sg13g2_xor2_1 _607_ (.B(BI),
    .A(B[11]),
    .X(_225_));
 sg13g2_nand2_1 _608_ (.Y(_226_),
    .A(A[11]),
    .B(_225_));
 sg13g2_inv_1 _609_ (.Y(X[11]),
    .A(net6619));
 sg13g2_xnor2_1 _610_ (.Y(_227_),
    .A(A[11]),
    .B(_225_));
 sg13g2_nor2_1 _611_ (.A(_220_),
    .B(_227_),
    .Y(_228_));
 sg13g2_and2_1 _612_ (.A(_212_),
    .B(_228_),
    .X(_229_));
 sg13g2_nor2b_1 _613_ (.A(_200_),
    .B_N(_229_),
    .Y(_230_));
 sg13g2_o21ai_1 _614_ (.B1(_226_),
    .Y(_231_),
    .A1(_219_),
    .A2(_227_));
 sg13g2_a21o_1 _615_ (.A2(_228_),
    .A1(_213_),
    .B1(_231_),
    .X(_232_));
 sg13g2_a221oi_1 _616_ (.B2(CO[3]),
    .C1(_232_),
    .B1(_230_),
    .A1(_198_),
    .Y(_233_),
    .A2(_229_));
 sg13g2_inv_1 _617_ (.Y(CO[11]),
    .A(_233_));
 sg13g2_xor2_1 _618_ (.B(BI),
    .A(B[12]),
    .X(_234_));
 sg13g2_nand2_1 _619_ (.Y(_235_),
    .A(A[12]),
    .B(_234_));
 sg13g2_inv_1 _620_ (.Y(X[12]),
    .A(_236_));
 sg13g2_xnor2_1 _621_ (.Y(_236_),
    .A(A[12]),
    .B(_234_));
 sg13g2_nor2_1 _622_ (.A(_227_),
    .B(_236_),
    .Y(_237_));
 sg13g2_o21ai_1 _623_ (.B1(_235_),
    .Y(_238_),
    .A1(_226_),
    .A2(_236_));
 sg13g2_a21oi_1 _624_ (.A1(_222_),
    .A2(_237_),
    .Y(_239_),
    .B1(_238_));
 sg13g2_nand2_1 _625_ (.Y(_240_),
    .A(_221_),
    .B(_237_));
 sg13g2_o21ai_1 _626_ (.B1(_239_),
    .Y(_241_),
    .A1(_207_),
    .A2(_240_));
 sg13g2_nor3_1 _627_ (.A(_177_),
    .B(_208_),
    .C(_240_),
    .Y(_242_));
 sg13g2_inv_1 _628_ (.Y(CO[12]),
    .A(_243_));
 sg13g2_nor2_1 _629_ (.A(_241_),
    .B(_242_),
    .Y(_243_));
 sg13g2_xor2_1 _630_ (.B(BI),
    .A(B[13]),
    .X(_244_));
 sg13g2_nand2_1 _631_ (.Y(_245_),
    .A(A[13]),
    .B(_244_));
 sg13g2_inv_1 _632_ (.Y(X[13]),
    .A(_246_));
 sg13g2_xnor2_1 _633_ (.Y(_246_),
    .A(A[13]),
    .B(_244_));
 sg13g2_nor2_1 _634_ (.A(_236_),
    .B(_246_),
    .Y(_247_));
 sg13g2_and2_1 _635_ (.A(_228_),
    .B(_247_),
    .X(_248_));
 sg13g2_nand2_1 _636_ (.Y(_249_),
    .A(_215_),
    .B(_248_));
 sg13g2_o21ai_1 _637_ (.B1(_245_),
    .Y(_250_),
    .A1(_235_),
    .A2(_246_));
 sg13g2_a21o_1 _638_ (.A2(_247_),
    .A1(_231_),
    .B1(_250_),
    .X(_251_));
 sg13g2_a21oi_1 _639_ (.A1(_214_),
    .A2(_248_),
    .Y(_252_),
    .B1(_251_));
 sg13g2_o21ai_1 _640_ (.B1(_252_),
    .Y(CO[13]),
    .A1(_185_),
    .A2(_249_));
 sg13g2_xor2_1 _641_ (.B(BI),
    .A(B[14]),
    .X(_253_));
 sg13g2_and2_1 _642_ (.A(A[14]),
    .B(_253_),
    .X(_254_));
 sg13g2_nand2_1 _643_ (.Y(_255_),
    .A(A[14]),
    .B(_253_));
 sg13g2_inv_1 _644_ (.Y(X[14]),
    .A(net6596));
 sg13g2_xnor2_1 _645_ (.Y(_256_),
    .A(A[14]),
    .B(_253_));
 sg13g2_nor2_1 _646_ (.A(_246_),
    .B(_256_),
    .Y(_257_));
 sg13g2_and2_1 _647_ (.A(_237_),
    .B(_257_),
    .X(_258_));
 sg13g2_nand2b_1 _648_ (.Y(_259_),
    .B(_258_),
    .A_N(_224_));
 sg13g2_o21ai_1 _649_ (.B1(_255_),
    .Y(_260_),
    .A1(_245_),
    .A2(_256_));
 sg13g2_a21oi_1 _650_ (.A1(_238_),
    .A2(_257_),
    .Y(_261_),
    .B1(_260_));
 sg13g2_nand2b_1 _651_ (.Y(_262_),
    .B(_258_),
    .A_N(_223_));
 sg13g2_and2_1 _652_ (.A(_261_),
    .B(_262_),
    .X(_263_));
 sg13g2_o21ai_1 _653_ (.B1(_263_),
    .Y(CO[14]),
    .A1(_192_),
    .A2(_259_));
 sg13g2_xor2_1 _654_ (.B(BI),
    .A(B[15]),
    .X(_264_));
 sg13g2_and2_1 _655_ (.A(A[15]),
    .B(_264_),
    .X(_265_));
 sg13g2_inv_1 _656_ (.Y(X[15]),
    .A(_266_));
 sg13g2_xnor2_1 _657_ (.Y(_266_),
    .A(A[15]),
    .B(_264_));
 sg13g2_nor2_1 _658_ (.A(_256_),
    .B(_266_),
    .Y(_267_));
 sg13g2_and2_1 _659_ (.A(_247_),
    .B(_267_),
    .X(_268_));
 sg13g2_and2_1 _660_ (.A(_229_),
    .B(_268_),
    .X(_269_));
 sg13g2_nand2_1 _661_ (.Y(_270_),
    .A(_250_),
    .B(_267_));
 sg13g2_a21oi_1 _662_ (.A1(_254_),
    .A2(X[15]),
    .Y(_271_),
    .B1(_265_));
 sg13g2_nand2_1 _663_ (.Y(_272_),
    .A(_270_),
    .B(_271_));
 sg13g2_a221oi_1 _664_ (.B2(CO[7]),
    .C1(_272_),
    .B1(_269_),
    .A1(_232_),
    .Y(_273_),
    .A2(_268_));
 sg13g2_inv_1 _665_ (.Y(CO[15]),
    .A(net6123));
 sg13g2_xor2_1 _666_ (.B(BI),
    .A(net6634),
    .X(_274_));
 sg13g2_and2_1 _667_ (.A(A[16]),
    .B(_274_),
    .X(_275_));
 sg13g2_or2_1 _668_ (.X(_276_),
    .B(_274_),
    .A(A[16]));
 sg13g2_inv_1 _669_ (.Y(X[16]),
    .A(net6594));
 sg13g2_xnor2_1 _670_ (.Y(_277_),
    .A(A[16]),
    .B(_274_));
 sg13g2_nor2_1 _671_ (.A(net6595),
    .B(net6594),
    .Y(_278_));
 sg13g2_a21o_1 _672_ (.A2(_276_),
    .A1(_265_),
    .B1(_275_),
    .X(_279_));
 sg13g2_a21oi_1 _673_ (.A1(_260_),
    .A2(_278_),
    .Y(_280_),
    .B1(_279_));
 sg13g2_nand2_1 _674_ (.Y(_281_),
    .A(net6556),
    .B(_278_));
 sg13g2_o21ai_1 _675_ (.B1(_280_),
    .Y(_282_),
    .A1(_239_),
    .A2(_281_));
 sg13g2_nor2_1 _676_ (.A(_240_),
    .B(_281_),
    .Y(_283_));
 sg13g2_a21oi_1 _677_ (.A1(CO[8]),
    .A2(_283_),
    .Y(_284_),
    .B1(_282_));
 sg13g2_inv_1 _678_ (.Y(CO[16]),
    .A(net6122));
 sg13g2_xor2_1 _679_ (.B(BI),
    .A(net6633),
    .X(_285_));
 sg13g2_and2_1 _680_ (.A(A[17]),
    .B(net6618),
    .X(_286_));
 sg13g2_nor2_1 _681_ (.A(A[17]),
    .B(net6618),
    .Y(_287_));
 sg13g2_xor2_1 _682_ (.B(_285_),
    .A(A[17]),
    .X(X[17]));
 sg13g2_nand2b_1 _683_ (.Y(_288_),
    .B(X[17]),
    .A_N(_277_));
 sg13g2_a21oi_1 _684_ (.A1(_275_),
    .A2(X[17]),
    .Y(_289_),
    .B1(_286_));
 sg13g2_o21ai_1 _685_ (.B1(_289_),
    .Y(_290_),
    .A1(_271_),
    .A2(net6555));
 sg13g2_nor3_1 _686_ (.A(net6596),
    .B(net6595),
    .C(_288_),
    .Y(_291_));
 sg13g2_a21oi_1 _687_ (.A1(_251_),
    .A2(_291_),
    .Y(_292_),
    .B1(_290_));
 sg13g2_nand2_1 _688_ (.Y(_293_),
    .A(net6477),
    .B(_291_));
 sg13g2_o21ai_1 _689_ (.B1(_292_),
    .Y(CO[17]),
    .A1(_217_),
    .A2(_293_));
 sg13g2_buf_1 place5957 (.A(_079_),
    .X(net5956));
 sg13g2_buf_1 place6123 (.A(_284_),
    .X(net6122));
 sg13g2_buf_1 place6124 (.A(_273_),
    .X(net6123));
 sg13g2_buf_1 place6125 (.A(_057_),
    .X(net6124));
 sg13g2_buf_1 place6397 (.A(_262_),
    .X(net6396));
 sg13g2_buf_1 place6402 (.A(_107_),
    .X(net6401));
 sg13g2_buf_1 place6403 (.A(_106_),
    .X(net6402));
 sg13g2_buf_1 place6404 (.A(_076_),
    .X(net6403));
 sg13g2_buf_1 place6405 (.A(_026_),
    .X(net6404));
 sg13g2_buf_1 place6476 (.A(_291_),
    .X(net6475));
 sg13g2_buf_1 place6477 (.A(_261_),
    .X(net6476));
 sg13g2_buf_1 place6478 (.A(_248_),
    .X(net6477));
 sg13g2_buf_1 place6481 (.A(_123_),
    .X(net6480));
 sg13g2_buf_1 place6482 (.A(_114_),
    .X(net6481));
 sg13g2_buf_1 place6483 (.A(_105_),
    .X(net6482));
 sg13g2_buf_1 place6484 (.A(_104_),
    .X(net6483));
 sg13g2_buf_1 place6485 (.A(_104_),
    .X(net6484));
 sg13g2_buf_1 place6486 (.A(_083_),
    .X(net6485));
 sg13g2_buf_1 place6487 (.A(_064_),
    .X(net6486));
 sg13g2_buf_1 place6556 (.A(_288_),
    .X(net6555));
 sg13g2_buf_1 place6557 (.A(_257_),
    .X(net6556));
 sg13g2_buf_1 place6559 (.A(_103_),
    .X(net6558));
 sg13g2_buf_1 place6560 (.A(_093_),
    .X(net6559));
 sg13g2_buf_1 place6561 (.A(_072_),
    .X(net6560));
 sg13g2_buf_1 place6562 (.A(_063_),
    .X(net6561));
 sg13g2_buf_1 place6563 (.A(_053_),
    .X(net6562));
 sg13g2_buf_1 place6564 (.A(_042_),
    .X(net6563));
 sg13g2_buf_1 place6565 (.A(_032_),
    .X(net6564));
 sg13g2_buf_1 place6566 (.A(_022_),
    .X(net6565));
 sg13g2_buf_1 place6567 (.A(_002_),
    .X(net6566));
 sg13g2_buf_2 place6594 (.A(A[27]),
    .X(net6593));
 sg13g2_buf_1 place6595 (.A(_277_),
    .X(net6594));
 sg13g2_buf_1 place6596 (.A(_266_),
    .X(net6595));
 sg13g2_buf_1 place6597 (.A(_256_),
    .X(net6596));
 sg13g2_buf_1 place6598 (.A(_192_),
    .X(net6597));
 sg13g2_buf_1 place6599 (.A(_101_),
    .X(net6598));
 sg13g2_buf_2 place6617 (.A(B[28]),
    .X(net6616));
 sg13g2_buf_1 place6619 (.A(_285_),
    .X(net6618));
 sg13g2_buf_1 place6620 (.A(_227_),
    .X(net6619));
 sg13g2_buf_2 place6634 (.A(B[17]),
    .X(net6633));
 sg13g2_buf_1 place6635 (.A(B[16]),
    .X(net6634));
endmodule
