module I2cGpioExpanderTop (io_address_0_PAD,
    io_address_1_PAD,
    io_address_2_PAD,
    io_clock_PAD,
    io_gpio_0_PAD,
    io_gpio_1_PAD,
    io_gpio_2_PAD,
    io_gpio_3_PAD,
    io_gpio_4_PAD,
    io_gpio_5_PAD,
    io_gpio_6_PAD,
    io_gpio_7_PAD,
    io_i2c_interrupt_PAD,
    io_i2c_scl_PAD,
    io_i2c_sda_PAD,
    io_reset_PAD);
 inout io_address_0_PAD;
 inout io_address_1_PAD;
 inout io_address_2_PAD;
 inout io_clock_PAD;
 inout io_gpio_0_PAD;
 inout io_gpio_1_PAD;
 inout io_gpio_2_PAD;
 inout io_gpio_3_PAD;
 inout io_gpio_4_PAD;
 inout io_gpio_5_PAD;
 inout io_gpio_6_PAD;
 inout io_gpio_7_PAD;
 inout io_i2c_interrupt_PAD;
 inout io_i2c_scl_PAD;
 inout io_i2c_sda_PAD;
 inout io_reset_PAD;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire net324;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire clknet_4_8_0_clock_regs;
 wire _0110_;
 wire net323;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire net322;
 wire _0116_;
 wire _0117_;
 wire clknet_4_10_0_clock_regs;
 wire _0119_;
 wire net299;
 wire net297;
 wire _0122_;
 wire clock_regs;
 wire _0124_;
 wire _0125_;
 wire net298;
 wire _0127_;
 wire net329;
 wire net316;
 wire net315;
 wire _0131_;
 wire net314;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire net313;
 wire _0137_;
 wire net312;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire net311;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire net310;
 wire clknet_4_7_0_clock_regs;
 wire net309;
 wire _0150_;
 wire _0151_;
 wire clknet_4_5_0_clock_regs;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire clknet_0_clock;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire net317;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire net308;
 wire _0169_;
 wire net307;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire net306;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire clknet_4_4_0_clock_regs;
 wire net318;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire net303;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire clknet_0_clock_regs;
 wire clknet_1_0__leaf_clock;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire net302;
 wire clknet_4_2_0_clock_regs;
 wire _0219_;
 wire net305;
 wire net304;
 wire net300;
 wire _0223_;
 wire _0224_;
 wire net320;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire net319;
 wire net295;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire net294;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire net293;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire net301;
 wire net292;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire net296;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire net291;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire net290;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire net289;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire net287;
 wire _0353_;
 wire net288;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire net286;
 wire net284;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire net285;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire net281;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire net283;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire net280;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire net282;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire net152;
 wire net30;
 wire clock;
 wire reset;
 wire sg13g2_IOPad_io_address_0_p2c;
 wire sg13g2_IOPad_io_address_1_p2c;
 wire sg13g2_IOPad_io_address_2_p2c;
 wire sg13g2_IOPad_io_gpio_0_c2p;
 wire sg13g2_IOPad_io_gpio_0_c2p_en;
 wire sg13g2_IOPad_io_gpio_0_p2c;
 wire sg13g2_IOPad_io_gpio_1_c2p;
 wire sg13g2_IOPad_io_gpio_1_c2p_en;
 wire sg13g2_IOPad_io_gpio_1_p2c;
 wire sg13g2_IOPad_io_gpio_2_c2p;
 wire sg13g2_IOPad_io_gpio_2_c2p_en;
 wire sg13g2_IOPad_io_gpio_2_p2c;
 wire sg13g2_IOPad_io_gpio_3_c2p;
 wire sg13g2_IOPad_io_gpio_3_c2p_en;
 wire sg13g2_IOPad_io_gpio_3_p2c;
 wire sg13g2_IOPad_io_gpio_4_c2p;
 wire sg13g2_IOPad_io_gpio_4_c2p_en;
 wire sg13g2_IOPad_io_gpio_4_p2c;
 wire sg13g2_IOPad_io_gpio_5_c2p;
 wire sg13g2_IOPad_io_gpio_5_c2p_en;
 wire sg13g2_IOPad_io_gpio_5_p2c;
 wire sg13g2_IOPad_io_gpio_6_c2p;
 wire sg13g2_IOPad_io_gpio_6_c2p_en;
 wire sg13g2_IOPad_io_gpio_6_p2c;
 wire sg13g2_IOPad_io_gpio_7_c2p;
 wire sg13g2_IOPad_io_gpio_7_c2p_en;
 wire sg13g2_IOPad_io_gpio_7_p2c;
 wire sg13g2_IOPad_io_i2c_scl_p2c;
 wire sg13g2_IOPad_io_i2c_sda_p2c;
 wire \system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[0] ;
 wire \system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[1] ;
 wire \system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[2] ;
 wire \system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[3] ;
 wire \system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[4] ;
 wire \system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[5] ;
 wire \system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[6] ;
 wire \system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[7] ;
 wire \system_expander.gpioCtrl_1.last[0] ;
 wire \system_expander.gpioCtrl_1.last[1] ;
 wire \system_expander.gpioCtrl_1.last[2] ;
 wire \system_expander.gpioCtrl_1.last[3] ;
 wire \system_expander.gpioCtrl_1.last[4] ;
 wire \system_expander.gpioCtrl_1.last[5] ;
 wire \system_expander.gpioCtrl_1.last[6] ;
 wire \system_expander.gpioCtrl_1.last[7] ;
 wire \system_expander.i2cConfig_latch ;
 wire \system_expander.i2cConfig_latchedAddress[0] ;
 wire \system_expander.i2cConfig_latchedAddress[1] ;
 wire \system_expander.i2cConfig_latchedAddress[2] ;
 wire \system_expander.i2cCtrl_io_cmd_payload_data[0] ;
 wire \system_expander.i2cCtrl_io_cmd_payload_data[1] ;
 wire \system_expander.i2cCtrl_io_cmd_payload_data[2] ;
 wire \system_expander.i2cCtrl_io_cmd_payload_data[3] ;
 wire \system_expander.i2cCtrl_io_cmd_payload_data[4] ;
 wire \system_expander.i2cCtrl_io_cmd_payload_data[5] ;
 wire \system_expander.i2cCtrl_io_cmd_payload_data[6] ;
 wire \system_expander.i2cCtrl_io_cmd_payload_data[7] ;
 wire \system_expander.i2cCtrl_io_cmd_payload_read ;
 wire \system_expander.i2cCtrl_io_cmd_payload_reg ;
 wire \system_expander.i2cCtrl_io_cmd_ready ;
 wire \system_expander.i2cCtrl_io_cmd_valid ;
 wire \system_expander.i2cCtrl_io_i2c_interrupts[0] ;
 wire \system_expander.i2cCtrl_io_i2c_scl_write ;
 wire \system_expander.i2cCtrl_io_i2c_sda_write ;
 wire \system_expander.i2cCtrl_io_interrupts[0] ;
 wire \system_expander.i2cCtrl_io_rsp_ready ;
 wire \system_expander.i2cCtrl_io_rsp_valid ;
 wire \system_expander.irq_fall_ctrl.io_masks[0] ;
 wire \system_expander.irq_fall_ctrl.io_masks[1] ;
 wire \system_expander.irq_fall_ctrl.io_masks[2] ;
 wire \system_expander.irq_fall_ctrl.io_masks[3] ;
 wire \system_expander.irq_fall_ctrl.io_masks[4] ;
 wire \system_expander.irq_fall_ctrl.io_masks[5] ;
 wire \system_expander.irq_fall_ctrl.io_masks[6] ;
 wire \system_expander.irq_fall_ctrl.io_masks[7] ;
 wire \system_expander.irq_fall_ctrl.pendings[0] ;
 wire \system_expander.irq_fall_ctrl.pendings[1] ;
 wire \system_expander.irq_fall_ctrl.pendings[2] ;
 wire \system_expander.irq_fall_ctrl.pendings[3] ;
 wire \system_expander.irq_fall_ctrl.pendings[4] ;
 wire \system_expander.irq_fall_ctrl.pendings[5] ;
 wire \system_expander.irq_fall_ctrl.pendings[6] ;
 wire \system_expander.irq_fall_ctrl.pendings[7] ;
 wire \system_expander.irq_high_ctrl.io_masks[0] ;
 wire \system_expander.irq_high_ctrl.io_masks[1] ;
 wire \system_expander.irq_high_ctrl.io_masks[2] ;
 wire \system_expander.irq_high_ctrl.io_masks[3] ;
 wire \system_expander.irq_high_ctrl.io_masks[4] ;
 wire \system_expander.irq_high_ctrl.io_masks[5] ;
 wire \system_expander.irq_high_ctrl.io_masks[6] ;
 wire \system_expander.irq_high_ctrl.io_masks[7] ;
 wire \system_expander.irq_high_ctrl.pendings[0] ;
 wire \system_expander.irq_high_ctrl.pendings[1] ;
 wire \system_expander.irq_high_ctrl.pendings[2] ;
 wire \system_expander.irq_high_ctrl.pendings[3] ;
 wire \system_expander.irq_high_ctrl.pendings[4] ;
 wire \system_expander.irq_high_ctrl.pendings[5] ;
 wire \system_expander.irq_high_ctrl.pendings[6] ;
 wire \system_expander.irq_high_ctrl.pendings[7] ;
 wire \system_expander.irq_low_ctrl.io_masks[0] ;
 wire \system_expander.irq_low_ctrl.io_masks[1] ;
 wire \system_expander.irq_low_ctrl.io_masks[2] ;
 wire \system_expander.irq_low_ctrl.io_masks[3] ;
 wire \system_expander.irq_low_ctrl.io_masks[4] ;
 wire \system_expander.irq_low_ctrl.io_masks[5] ;
 wire \system_expander.irq_low_ctrl.io_masks[6] ;
 wire \system_expander.irq_low_ctrl.io_masks[7] ;
 wire \system_expander.irq_low_ctrl.pendings[0] ;
 wire \system_expander.irq_low_ctrl.pendings[1] ;
 wire \system_expander.irq_low_ctrl.pendings[2] ;
 wire \system_expander.irq_low_ctrl.pendings[3] ;
 wire \system_expander.irq_low_ctrl.pendings[4] ;
 wire \system_expander.irq_low_ctrl.pendings[5] ;
 wire \system_expander.irq_low_ctrl.pendings[6] ;
 wire \system_expander.irq_low_ctrl.pendings[7] ;
 wire \system_expander.irq_rise_ctrl.io_masks[0] ;
 wire \system_expander.irq_rise_ctrl.io_masks[1] ;
 wire \system_expander.irq_rise_ctrl.io_masks[2] ;
 wire \system_expander.irq_rise_ctrl.io_masks[3] ;
 wire \system_expander.irq_rise_ctrl.io_masks[4] ;
 wire \system_expander.irq_rise_ctrl.io_masks[5] ;
 wire \system_expander.irq_rise_ctrl.io_masks[6] ;
 wire \system_expander.irq_rise_ctrl.io_masks[7] ;
 wire \system_expander.irq_rise_ctrl.pendings[0] ;
 wire \system_expander.irq_rise_ctrl.pendings[1] ;
 wire \system_expander.irq_rise_ctrl.pendings[2] ;
 wire \system_expander.irq_rise_ctrl.pendings[3] ;
 wire \system_expander.irq_rise_ctrl.pendings[4] ;
 wire \system_expander.irq_rise_ctrl.pendings[5] ;
 wire \system_expander.irq_rise_ctrl.pendings[6] ;
 wire \system_expander.irq_rise_ctrl.pendings[7] ;
 wire \system_expander.link_data[0] ;
 wire \system_expander.link_data[1] ;
 wire \system_expander.link_data[2] ;
 wire \system_expander.link_data[3] ;
 wire \system_expander.link_data[4] ;
 wire \system_expander.link_data[5] ;
 wire \system_expander.link_data[6] ;
 wire \system_expander.link_data[7] ;
 wire \system_expander.link_error ;
 wire \system_expander.link_regAddr[0] ;
 wire \system_expander.link_regAddr[1] ;
 wire \system_expander.link_regAddr[2] ;
 wire \system_expander.link_regAddr[3] ;
 wire \system_expander.link_regAddr[4] ;
 wire \system_expander.link_regAddr[5] ;
 wire \system_expander.link_regAddr[6] ;
 wire \system_expander.link_regAddr[7] ;
 wire \system_expander.link_state[0] ;
 wire \system_expander.link_state[1] ;
 wire \system_expander.link_state[2] ;
 wire \system_expander.link_state[3] ;
 wire \system_expander.link_state[4] ;
 wire net325;
 wire net;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net326;
 wire net327;
 wire net328;
 wire clknet_4_9_0_clock_regs;
 wire net276;
 wire net278;
 wire net277;
 wire net279;
 wire net321;
 wire clknet_4_1_0_clock_regs;
 wire clknet_4_0_0_clock_regs;
 wire clknet_4_3_0_clock_regs;
 wire clknet_4_6_0_clock_regs;
 wire clknet_4_11_0_clock_regs;
 wire clknet_4_12_0_clock_regs;
 wire clknet_4_13_0_clock_regs;
 wire clknet_4_14_0_clock_regs;
 wire clknet_4_15_0_clock_regs;
 wire clknet_5_0__leaf_clock_regs;
 wire clknet_5_1__leaf_clock_regs;
 wire clknet_5_2__leaf_clock_regs;
 wire clknet_5_3__leaf_clock_regs;
 wire clknet_5_4__leaf_clock_regs;
 wire clknet_5_5__leaf_clock_regs;
 wire clknet_5_6__leaf_clock_regs;
 wire clknet_5_7__leaf_clock_regs;
 wire clknet_5_8__leaf_clock_regs;
 wire clknet_5_9__leaf_clock_regs;
 wire clknet_5_10__leaf_clock_regs;
 wire clknet_5_11__leaf_clock_regs;
 wire clknet_5_12__leaf_clock_regs;
 wire clknet_5_13__leaf_clock_regs;
 wire clknet_5_14__leaf_clock_regs;
 wire clknet_5_15__leaf_clock_regs;
 wire clknet_5_16__leaf_clock_regs;
 wire clknet_5_17__leaf_clock_regs;
 wire clknet_5_18__leaf_clock_regs;
 wire clknet_5_19__leaf_clock_regs;
 wire clknet_5_20__leaf_clock_regs;
 wire clknet_5_21__leaf_clock_regs;
 wire clknet_5_22__leaf_clock_regs;
 wire clknet_5_23__leaf_clock_regs;
 wire clknet_5_24__leaf_clock_regs;
 wire clknet_5_25__leaf_clock_regs;
 wire clknet_5_26__leaf_clock_regs;
 wire clknet_5_27__leaf_clock_regs;
 wire clknet_5_28__leaf_clock_regs;
 wire clknet_5_29__leaf_clock_regs;
 wire clknet_5_30__leaf_clock_regs;
 wire clknet_5_31__leaf_clock_regs;
 wire delaynet_0_clk_core;
 wire delaynet_1_clk_core;
 wire delaynet_2_clk_core;

 I2cDeviceCtrl \system_expander.i2cCtrl  (.clock(clknet_1_0__leaf_clock),
    .io_cmd_payload_read(\system_expander.i2cCtrl_io_cmd_payload_read ),
    .io_cmd_payload_reg(\system_expander.i2cCtrl_io_cmd_payload_reg ),
    .io_cmd_ready(\system_expander.i2cCtrl_io_cmd_ready ),
    .io_cmd_valid(\system_expander.i2cCtrl_io_cmd_valid ),
    .io_i2c_scl_read(sg13g2_IOPad_io_i2c_scl_p2c),
    .io_i2c_scl_write(\system_expander.i2cCtrl_io_i2c_scl_write ),
    .io_i2c_sda_read(sg13g2_IOPad_io_i2c_sda_p2c),
    .io_i2c_sda_write(\system_expander.i2cCtrl_io_i2c_sda_write ),
    .io_rsp_payload_error(\system_expander.link_error ),
    .io_rsp_ready(\system_expander.i2cCtrl_io_rsp_ready ),
    .io_rsp_valid(\system_expander.i2cCtrl_io_rsp_valid ),
    .reset(reset),
    .io_cmd_payload_data({\system_expander.i2cCtrl_io_cmd_payload_data[7] ,
    \system_expander.i2cCtrl_io_cmd_payload_data[6] ,
    \system_expander.i2cCtrl_io_cmd_payload_data[5] ,
    \system_expander.i2cCtrl_io_cmd_payload_data[4] ,
    \system_expander.i2cCtrl_io_cmd_payload_data[3] ,
    \system_expander.i2cCtrl_io_cmd_payload_data[2] ,
    \system_expander.i2cCtrl_io_cmd_payload_data[1] ,
    \system_expander.i2cCtrl_io_cmd_payload_data[0] }),
    .io_config_clockDivider({net7,
    net6,
    net5,
    net4,
    net3,
    net2,
    net16,
    net15,
    net14,
    net13,
    net12,
    net11,
    net10,
    net9,
    net8,
    net58}),
    .io_config_deviceAddr({net18,
    net60,
    net59,
    net17,
    \system_expander.i2cConfig_latchedAddress[2] ,
    \system_expander.i2cConfig_latchedAddress[1] ,
    \system_expander.i2cConfig_latchedAddress[0] }),
    .io_config_timeout({net24,
    net23,
    net22,
    net61,
    net21,
    net20,
    net65,
    net64,
    net63,
    net29,
    net28,
    net27,
    net62,
    net26,
    net25,
    net19}),
    .io_i2c_interrupts({\system_expander.i2cCtrl_io_i2c_interrupts[0] }),
    .io_interrupts({\system_expander.i2cCtrl_io_interrupts[0] }),
    .io_rsp_payload_data({\system_expander.link_data[7] ,
    \system_expander.link_data[6] ,
    \system_expander.link_data[5] ,
    \system_expander.link_data[4] ,
    \system_expander.link_data[3] ,
    \system_expander.link_data[2] ,
    \system_expander.link_data[1] ,
    \system_expander.link_data[0] }));
endmodule
