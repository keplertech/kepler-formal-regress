module I2cGpioExpanderTop (io_address_0_PAD,
    io_address_1_PAD,
    io_address_2_PAD,
    io_clock_PAD,
    io_gpio_0_PAD,
    io_gpio_1_PAD,
    io_gpio_2_PAD,
    io_gpio_3_PAD,
    io_gpio_4_PAD,
    io_gpio_5_PAD,
    io_gpio_6_PAD,
    io_gpio_7_PAD,
    io_i2c_interrupt_PAD,
    io_i2c_scl_PAD,
    io_i2c_sda_PAD,
    io_reset_PAD);
 inout io_address_0_PAD;
 inout io_address_1_PAD;
 inout io_address_2_PAD;
 inout io_clock_PAD;
 inout io_gpio_0_PAD;
 inout io_gpio_1_PAD;
 inout io_gpio_2_PAD;
 inout io_gpio_3_PAD;
 inout io_gpio_4_PAD;
 inout io_gpio_5_PAD;
 inout io_gpio_6_PAD;
 inout io_gpio_7_PAD;
 inout io_i2c_interrupt_PAD;
 inout io_i2c_scl_PAD;
 inout io_i2c_sda_PAD;
 inout io_reset_PAD;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire net324;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire clknet_4_8_0_clock_regs;
 wire _0110_;
 wire net323;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire net322;
 wire _0116_;
 wire _0117_;
 wire clknet_4_10_0_clock_regs;
 wire _0119_;
 wire net299;
 wire net297;
 wire _0122_;
 wire clock_regs;
 wire _0124_;
 wire _0125_;
 wire net298;
 wire _0127_;
 wire net329;
 wire net316;
 wire net315;
 wire _0131_;
 wire net314;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire net313;
 wire _0137_;
 wire net312;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire net311;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire net310;
 wire clknet_4_7_0_clock_regs;
 wire net309;
 wire _0150_;
 wire _0151_;
 wire clknet_4_5_0_clock_regs;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire clknet_0_clock;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire net317;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire net308;
 wire _0169_;
 wire net307;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire net306;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire clknet_4_4_0_clock_regs;
 wire net318;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire net303;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire clknet_0_clock_regs;
 wire clknet_1_0__leaf_clock;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire net302;
 wire clknet_4_2_0_clock_regs;
 wire _0219_;
 wire net305;
 wire net304;
 wire net300;
 wire _0223_;
 wire _0224_;
 wire net320;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire net319;
 wire net295;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire net294;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire net293;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire net301;
 wire net292;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire net296;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire net291;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire net290;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire net289;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire net287;
 wire _0353_;
 wire net288;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire net286;
 wire net284;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire net285;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire net281;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire net283;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire net280;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire net282;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire net152;
 wire net30;
 wire clock;
 wire reset;
 wire sg13g2_IOPad_io_address_0_p2c;
 wire sg13g2_IOPad_io_address_1_p2c;
 wire sg13g2_IOPad_io_address_2_p2c;
 wire sg13g2_IOPad_io_gpio_0_c2p;
 wire sg13g2_IOPad_io_gpio_0_c2p_en;
 wire sg13g2_IOPad_io_gpio_0_p2c;
 wire sg13g2_IOPad_io_gpio_1_c2p;
 wire sg13g2_IOPad_io_gpio_1_c2p_en;
 wire sg13g2_IOPad_io_gpio_1_p2c;
 wire sg13g2_IOPad_io_gpio_2_c2p;
 wire sg13g2_IOPad_io_gpio_2_c2p_en;
 wire sg13g2_IOPad_io_gpio_2_p2c;
 wire sg13g2_IOPad_io_gpio_3_c2p;
 wire sg13g2_IOPad_io_gpio_3_c2p_en;
 wire sg13g2_IOPad_io_gpio_3_p2c;
 wire sg13g2_IOPad_io_gpio_4_c2p;
 wire sg13g2_IOPad_io_gpio_4_c2p_en;
 wire sg13g2_IOPad_io_gpio_4_p2c;
 wire sg13g2_IOPad_io_gpio_5_c2p;
 wire sg13g2_IOPad_io_gpio_5_c2p_en;
 wire sg13g2_IOPad_io_gpio_5_p2c;
 wire sg13g2_IOPad_io_gpio_6_c2p;
 wire sg13g2_IOPad_io_gpio_6_c2p_en;
 wire sg13g2_IOPad_io_gpio_6_p2c;
 wire sg13g2_IOPad_io_gpio_7_c2p;
 wire sg13g2_IOPad_io_gpio_7_c2p_en;
 wire sg13g2_IOPad_io_gpio_7_p2c;
 wire sg13g2_IOPad_io_i2c_scl_p2c;
 wire sg13g2_IOPad_io_i2c_sda_p2c;
 wire \system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[0] ;
 wire \system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[1] ;
 wire \system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[2] ;
 wire \system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[3] ;
 wire \system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[4] ;
 wire \system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[5] ;
 wire \system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[6] ;
 wire \system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[7] ;
 wire \system_expander.gpioCtrl_1.last[0] ;
 wire \system_expander.gpioCtrl_1.last[1] ;
 wire \system_expander.gpioCtrl_1.last[2] ;
 wire \system_expander.gpioCtrl_1.last[3] ;
 wire \system_expander.gpioCtrl_1.last[4] ;
 wire \system_expander.gpioCtrl_1.last[5] ;
 wire \system_expander.gpioCtrl_1.last[6] ;
 wire \system_expander.gpioCtrl_1.last[7] ;
 wire \system_expander.i2cConfig_latch ;
 wire \system_expander.i2cConfig_latchedAddress[0] ;
 wire \system_expander.i2cConfig_latchedAddress[1] ;
 wire \system_expander.i2cConfig_latchedAddress[2] ;
 wire \system_expander.i2cCtrl_io_cmd_payload_data[0] ;
 wire \system_expander.i2cCtrl_io_cmd_payload_data[1] ;
 wire \system_expander.i2cCtrl_io_cmd_payload_data[2] ;
 wire \system_expander.i2cCtrl_io_cmd_payload_data[3] ;
 wire \system_expander.i2cCtrl_io_cmd_payload_data[4] ;
 wire \system_expander.i2cCtrl_io_cmd_payload_data[5] ;
 wire \system_expander.i2cCtrl_io_cmd_payload_data[6] ;
 wire \system_expander.i2cCtrl_io_cmd_payload_data[7] ;
 wire \system_expander.i2cCtrl_io_cmd_payload_read ;
 wire \system_expander.i2cCtrl_io_cmd_payload_reg ;
 wire \system_expander.i2cCtrl_io_cmd_ready ;
 wire \system_expander.i2cCtrl_io_cmd_valid ;
 wire \system_expander.i2cCtrl_io_i2c_interrupts[0] ;
 wire \system_expander.i2cCtrl_io_i2c_scl_write ;
 wire \system_expander.i2cCtrl_io_i2c_sda_write ;
 wire \system_expander.i2cCtrl_io_interrupts[0] ;
 wire \system_expander.i2cCtrl_io_rsp_ready ;
 wire \system_expander.i2cCtrl_io_rsp_valid ;
 wire \system_expander.irq_fall_ctrl.io_masks[0] ;
 wire \system_expander.irq_fall_ctrl.io_masks[1] ;
 wire \system_expander.irq_fall_ctrl.io_masks[2] ;
 wire \system_expander.irq_fall_ctrl.io_masks[3] ;
 wire \system_expander.irq_fall_ctrl.io_masks[4] ;
 wire \system_expander.irq_fall_ctrl.io_masks[5] ;
 wire \system_expander.irq_fall_ctrl.io_masks[6] ;
 wire \system_expander.irq_fall_ctrl.io_masks[7] ;
 wire \system_expander.irq_fall_ctrl.pendings[0] ;
 wire \system_expander.irq_fall_ctrl.pendings[1] ;
 wire \system_expander.irq_fall_ctrl.pendings[2] ;
 wire \system_expander.irq_fall_ctrl.pendings[3] ;
 wire \system_expander.irq_fall_ctrl.pendings[4] ;
 wire \system_expander.irq_fall_ctrl.pendings[5] ;
 wire \system_expander.irq_fall_ctrl.pendings[6] ;
 wire \system_expander.irq_fall_ctrl.pendings[7] ;
 wire \system_expander.irq_high_ctrl.io_masks[0] ;
 wire \system_expander.irq_high_ctrl.io_masks[1] ;
 wire \system_expander.irq_high_ctrl.io_masks[2] ;
 wire \system_expander.irq_high_ctrl.io_masks[3] ;
 wire \system_expander.irq_high_ctrl.io_masks[4] ;
 wire \system_expander.irq_high_ctrl.io_masks[5] ;
 wire \system_expander.irq_high_ctrl.io_masks[6] ;
 wire \system_expander.irq_high_ctrl.io_masks[7] ;
 wire \system_expander.irq_high_ctrl.pendings[0] ;
 wire \system_expander.irq_high_ctrl.pendings[1] ;
 wire \system_expander.irq_high_ctrl.pendings[2] ;
 wire \system_expander.irq_high_ctrl.pendings[3] ;
 wire \system_expander.irq_high_ctrl.pendings[4] ;
 wire \system_expander.irq_high_ctrl.pendings[5] ;
 wire \system_expander.irq_high_ctrl.pendings[6] ;
 wire \system_expander.irq_high_ctrl.pendings[7] ;
 wire \system_expander.irq_low_ctrl.io_masks[0] ;
 wire \system_expander.irq_low_ctrl.io_masks[1] ;
 wire \system_expander.irq_low_ctrl.io_masks[2] ;
 wire \system_expander.irq_low_ctrl.io_masks[3] ;
 wire \system_expander.irq_low_ctrl.io_masks[4] ;
 wire \system_expander.irq_low_ctrl.io_masks[5] ;
 wire \system_expander.irq_low_ctrl.io_masks[6] ;
 wire \system_expander.irq_low_ctrl.io_masks[7] ;
 wire \system_expander.irq_low_ctrl.pendings[0] ;
 wire \system_expander.irq_low_ctrl.pendings[1] ;
 wire \system_expander.irq_low_ctrl.pendings[2] ;
 wire \system_expander.irq_low_ctrl.pendings[3] ;
 wire \system_expander.irq_low_ctrl.pendings[4] ;
 wire \system_expander.irq_low_ctrl.pendings[5] ;
 wire \system_expander.irq_low_ctrl.pendings[6] ;
 wire \system_expander.irq_low_ctrl.pendings[7] ;
 wire \system_expander.irq_rise_ctrl.io_masks[0] ;
 wire \system_expander.irq_rise_ctrl.io_masks[1] ;
 wire \system_expander.irq_rise_ctrl.io_masks[2] ;
 wire \system_expander.irq_rise_ctrl.io_masks[3] ;
 wire \system_expander.irq_rise_ctrl.io_masks[4] ;
 wire \system_expander.irq_rise_ctrl.io_masks[5] ;
 wire \system_expander.irq_rise_ctrl.io_masks[6] ;
 wire \system_expander.irq_rise_ctrl.io_masks[7] ;
 wire \system_expander.irq_rise_ctrl.pendings[0] ;
 wire \system_expander.irq_rise_ctrl.pendings[1] ;
 wire \system_expander.irq_rise_ctrl.pendings[2] ;
 wire \system_expander.irq_rise_ctrl.pendings[3] ;
 wire \system_expander.irq_rise_ctrl.pendings[4] ;
 wire \system_expander.irq_rise_ctrl.pendings[5] ;
 wire \system_expander.irq_rise_ctrl.pendings[6] ;
 wire \system_expander.irq_rise_ctrl.pendings[7] ;
 wire \system_expander.link_data[0] ;
 wire \system_expander.link_data[1] ;
 wire \system_expander.link_data[2] ;
 wire \system_expander.link_data[3] ;
 wire \system_expander.link_data[4] ;
 wire \system_expander.link_data[5] ;
 wire \system_expander.link_data[6] ;
 wire \system_expander.link_data[7] ;
 wire \system_expander.link_error ;
 wire \system_expander.link_regAddr[0] ;
 wire \system_expander.link_regAddr[1] ;
 wire \system_expander.link_regAddr[2] ;
 wire \system_expander.link_regAddr[3] ;
 wire \system_expander.link_regAddr[4] ;
 wire \system_expander.link_regAddr[5] ;
 wire \system_expander.link_regAddr[6] ;
 wire \system_expander.link_regAddr[7] ;
 wire \system_expander.link_state[0] ;
 wire \system_expander.link_state[1] ;
 wire \system_expander.link_state[2] ;
 wire \system_expander.link_state[3] ;
 wire \system_expander.link_state[4] ;
 wire net325;
 wire net;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net326;
 wire net327;
 wire net328;
 wire clknet_4_9_0_clock_regs;
 wire net276;
 wire net278;
 wire net277;
 wire net279;
 wire net321;
 wire clknet_4_1_0_clock_regs;
 wire clknet_4_0_0_clock_regs;
 wire clknet_4_3_0_clock_regs;
 wire clknet_4_6_0_clock_regs;
 wire clknet_4_11_0_clock_regs;
 wire clknet_4_12_0_clock_regs;
 wire clknet_4_13_0_clock_regs;
 wire clknet_4_14_0_clock_regs;
 wire clknet_4_15_0_clock_regs;
 wire clknet_5_0__leaf_clock_regs;
 wire clknet_5_1__leaf_clock_regs;
 wire clknet_5_2__leaf_clock_regs;
 wire clknet_5_3__leaf_clock_regs;
 wire clknet_5_4__leaf_clock_regs;
 wire clknet_5_5__leaf_clock_regs;
 wire clknet_5_6__leaf_clock_regs;
 wire clknet_5_7__leaf_clock_regs;
 wire clknet_5_8__leaf_clock_regs;
 wire clknet_5_9__leaf_clock_regs;
 wire clknet_5_10__leaf_clock_regs;
 wire clknet_5_11__leaf_clock_regs;
 wire clknet_5_12__leaf_clock_regs;
 wire clknet_5_13__leaf_clock_regs;
 wire clknet_5_14__leaf_clock_regs;
 wire clknet_5_15__leaf_clock_regs;
 wire clknet_5_16__leaf_clock_regs;
 wire clknet_5_17__leaf_clock_regs;
 wire clknet_5_18__leaf_clock_regs;
 wire clknet_5_19__leaf_clock_regs;
 wire clknet_5_20__leaf_clock_regs;
 wire clknet_5_21__leaf_clock_regs;
 wire clknet_5_22__leaf_clock_regs;
 wire clknet_5_23__leaf_clock_regs;
 wire clknet_5_24__leaf_clock_regs;
 wire clknet_5_25__leaf_clock_regs;
 wire clknet_5_26__leaf_clock_regs;
 wire clknet_5_27__leaf_clock_regs;
 wire clknet_5_28__leaf_clock_regs;
 wire clknet_5_29__leaf_clock_regs;
 wire clknet_5_30__leaf_clock_regs;
 wire clknet_5_31__leaf_clock_regs;
 wire delaynet_0_clk_core;
 wire delaynet_1_clk_core;
 wire delaynet_2_clk_core;

 bondpad_70x70 IO_BOND_sg13g2_IOPadIOVdd_west_4 (.pad(IOVDD));
 bondpad_70x70 IO_BOND_sg13g2_IOPadIOVss_west_3 (.pad(IOVSS));
 bondpad_70x70 IO_BOND_sg13g2_IOPadVdd_east_0 (.pad(VDD));
 bondpad_70x70 IO_BOND_sg13g2_IOPadVss_east_1 (.pad(VSS));
 bondpad_70x70 IO_BOND_sg13g2_IOPad_io_address_0 (.pad(io_address_0_PAD));
 bondpad_70x70 IO_BOND_sg13g2_IOPad_io_address_1 (.pad(io_address_1_PAD));
 bondpad_70x70 IO_BOND_sg13g2_IOPad_io_address_2 (.pad(io_address_2_PAD));
 bondpad_70x70 IO_BOND_sg13g2_IOPad_io_clock (.pad(io_clock_PAD));
 bondpad_70x70 IO_BOND_sg13g2_IOPad_io_gpio_0 (.pad(io_gpio_0_PAD));
 bondpad_70x70 IO_BOND_sg13g2_IOPad_io_gpio_1 (.pad(io_gpio_1_PAD));
 bondpad_70x70 IO_BOND_sg13g2_IOPad_io_gpio_2 (.pad(io_gpio_2_PAD));
 bondpad_70x70 IO_BOND_sg13g2_IOPad_io_gpio_3 (.pad(io_gpio_3_PAD));
 bondpad_70x70 IO_BOND_sg13g2_IOPad_io_gpio_4 (.pad(io_gpio_4_PAD));
 bondpad_70x70 IO_BOND_sg13g2_IOPad_io_gpio_5 (.pad(io_gpio_5_PAD));
 bondpad_70x70 IO_BOND_sg13g2_IOPad_io_gpio_6 (.pad(io_gpio_6_PAD));
 bondpad_70x70 IO_BOND_sg13g2_IOPad_io_gpio_7 (.pad(io_gpio_7_PAD));
 bondpad_70x70 IO_BOND_sg13g2_IOPad_io_i2c_interrupt (.pad(io_i2c_interrupt_PAD));
 bondpad_70x70 IO_BOND_sg13g2_IOPad_io_i2c_scl (.pad(io_i2c_scl_PAD));
 bondpad_70x70 IO_BOND_sg13g2_IOPad_io_i2c_sda (.pad(io_i2c_sda_PAD));
 bondpad_70x70 IO_BOND_sg13g2_IOPad_io_reset (.pad(io_reset_PAD));
 sg13g2_Corner IO_CORNER_NORTH_EAST_INST ();
 sg13g2_Corner IO_CORNER_NORTH_WEST_INST ();
 sg13g2_Corner IO_CORNER_SOUTH_EAST_INST ();
 sg13g2_Corner IO_CORNER_SOUTH_WEST_INST ();
 sg13g2_Filler200 IO_FILL_IO_EAST_0_0 ();
 sg13g2_Filler400 IO_FILL_IO_EAST_1_0 ();
 sg13g2_Filler400 IO_FILL_IO_EAST_2_0 ();
 sg13g2_Filler400 IO_FILL_IO_EAST_3_0 ();
 sg13g2_Filler200 IO_FILL_IO_EAST_3_2 ();
 sg13g2_Filler400 IO_FILL_IO_EAST_4_0 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_0_0 ();
 sg13g2_Filler400 IO_FILL_IO_NORTH_1_0 ();
 sg13g2_Filler400 IO_FILL_IO_NORTH_2_0 ();
 sg13g2_Filler400 IO_FILL_IO_NORTH_3_0 ();
 sg13g2_Filler400 IO_FILL_IO_NORTH_4_0 ();
 sg13g2_Filler200 IO_FILL_IO_NORTH_5_0 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_0_0 ();
 sg13g2_Filler400 IO_FILL_IO_SOUTH_1_0 ();
 sg13g2_Filler400 IO_FILL_IO_SOUTH_2_0 ();
 sg13g2_Filler400 IO_FILL_IO_SOUTH_3_0 ();
 sg13g2_Filler400 IO_FILL_IO_SOUTH_4_0 ();
 sg13g2_Filler200 IO_FILL_IO_SOUTH_5_0 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_0_0 ();
 sg13g2_Filler400 IO_FILL_IO_WEST_1_0 ();
 sg13g2_Filler400 IO_FILL_IO_WEST_2_0 ();
 sg13g2_Filler400 IO_FILL_IO_WEST_3_0 ();
 sg13g2_Filler200 IO_FILL_IO_WEST_3_2 ();
 sg13g2_Filler400 IO_FILL_IO_WEST_4_0 ();
 sg13g2_nand3_1 _0579_ (.B(\system_expander.i2cCtrl_io_cmd_valid ),
    .C(\system_expander.link_state[0] ),
    .A(reset),
    .Y(_0106_));
 sg13g2_nor3_1 _0580_ (.A(\system_expander.i2cCtrl_io_cmd_payload_read ),
    .B(\system_expander.i2cCtrl_io_cmd_payload_reg ),
    .C(_0106_),
    .Y(_0002_));
 sg13g2_inv_1 _0581_ (.Y(_0107_),
    .A(\system_expander.i2cCtrl_io_cmd_payload_reg ));
 sg13g2_nor3_1 _0582_ (.A(\system_expander.i2cCtrl_io_cmd_payload_read ),
    .B(_0107_),
    .C(_0106_),
    .Y(_0001_));
 sg13g2_inv_1 _0583_ (.Y(_0108_),
    .A(\system_expander.i2cCtrl_io_cmd_payload_read ));
 sg13g2_nor2_1 _0584_ (.A(_0108_),
    .B(_0106_),
    .Y(_0000_));
 sg13g2_or2_1 _0586_ (.X(_0110_),
    .B(\system_expander.link_state[4] ),
    .A(\system_expander.link_state[2] ));
 sg13g2_nor2_1 _0588_ (.A(\system_expander.link_state[3] ),
    .B(_0110_),
    .Y(_0112_));
 sg13g2_nand2b_1 _0589_ (.Y(_0113_),
    .B(\system_expander.link_state[1] ),
    .A_N(\system_expander.i2cCtrl_io_rsp_ready ));
 sg13g2_inv_1 _0590_ (.Y(_0114_),
    .A(reset));
 sg13g2_a21oi_1 _0592_ (.A1(_0112_),
    .A2(_0113_),
    .Y(_0004_),
    .B1(_0114_));
 sg13g2_inv_1 _0593_ (.Y(_0116_),
    .A(\system_expander.i2cCtrl_io_cmd_valid ));
 sg13g2_a22oi_1 _0594_ (.Y(_0117_),
    .B1(\system_expander.i2cCtrl_io_rsp_ready ),
    .B2(\system_expander.link_state[1] ),
    .A2(\system_expander.link_state[0] ),
    .A1(_0116_));
 sg13g2_nand2_1 _0595_ (.Y(_0003_),
    .A(reset),
    .B(_0117_));
 sg13g2_nor2_1 _0597_ (.A(\system_expander.link_state[2] ),
    .B(\system_expander.link_state[4] ),
    .Y(_0119_));
 sg13g2_inv_1 _0600_ (.Y(_0122_),
    .A(net307));
 sg13g2_nand2_1 _0602_ (.Y(_0124_),
    .A(\system_expander.link_state[3] ),
    .B(\system_expander.i2cCtrl_io_cmd_payload_data[0] ));
 sg13g2_o21ai_1 _0603_ (.B1(_0124_),
    .Y(_0125_),
    .A1(\system_expander.link_state[3] ),
    .A2(_0122_));
 sg13g2_nor2_1 _0605_ (.A(\system_expander.link_regAddr[0] ),
    .B(_0119_),
    .Y(_0127_));
 sg13g2_a21o_1 _0606_ (.A2(_0125_),
    .A1(net294),
    .B1(_0127_),
    .X(_0097_));
 sg13g2_o21ai_1 _0610_ (.B1(\system_expander.link_regAddr[1] ),
    .Y(_0131_),
    .A1(_0112_),
    .A2(_0127_));
 sg13g2_and2_1 _0612_ (.A(\system_expander.link_state[3] ),
    .B(net294),
    .X(_0133_));
 sg13g2_nor2_1 _0613_ (.A(_0122_),
    .B(net305),
    .Y(_0134_));
 sg13g2_a22oi_1 _0614_ (.Y(_0135_),
    .B1(_0134_),
    .B2(_0110_),
    .A2(_0133_),
    .A1(\system_expander.i2cCtrl_io_cmd_payload_data[1] ));
 sg13g2_nand2_1 _0615_ (.Y(_0098_),
    .A(_0131_),
    .B(_0135_));
 sg13g2_and3_1 _0617_ (.X(_0137_),
    .A(\system_expander.link_regAddr[0] ),
    .B(\system_expander.link_regAddr[1] ),
    .C(\system_expander.link_regAddr[2] ));
 sg13g2_and2_1 _0619_ (.A(net307),
    .B(\system_expander.link_regAddr[1] ),
    .X(_0139_));
 sg13g2_inv_1 _0620_ (.Y(\system_expander.i2cCtrl_io_cmd_ready ),
    .A(_0112_));
 sg13g2_o21ai_1 _0621_ (.B1(\system_expander.i2cCtrl_io_cmd_ready ),
    .Y(_0140_),
    .A1(_0119_),
    .A2(_0139_));
 sg13g2_inv_1 _0622_ (.Y(_0141_),
    .A(\system_expander.link_regAddr[2] ));
 sg13g2_nand2_1 _0624_ (.Y(_0143_),
    .A(\system_expander.link_state[3] ),
    .B(net294));
 sg13g2_nor2_1 _0625_ (.A(\system_expander.i2cCtrl_io_cmd_payload_data[2] ),
    .B(_0143_),
    .Y(_0144_));
 sg13g2_a221oi_1 _0626_ (.B2(_0141_),
    .C1(_0144_),
    .B1(_0140_),
    .A1(_0110_),
    .Y(_0099_),
    .A2(_0137_));
 sg13g2_inv_2 _0627_ (.Y(_0145_),
    .A(\system_expander.link_regAddr[3] ));
 sg13g2_o21ai_1 _0628_ (.B1(\system_expander.i2cCtrl_io_cmd_ready ),
    .Y(_0146_),
    .A1(net294),
    .A2(_0137_));
 sg13g2_nand3_1 _0632_ (.B(_0110_),
    .C(_0137_),
    .A(\system_expander.link_regAddr[3] ),
    .Y(_0150_));
 sg13g2_o21ai_1 _0633_ (.B1(_0150_),
    .Y(_0151_),
    .A1(net312),
    .A2(_0143_));
 sg13g2_a21oi_1 _0634_ (.A1(_0145_),
    .A2(_0146_),
    .Y(_0100_),
    .B1(_0151_));
 sg13g2_inv_1 _0636_ (.Y(_0153_),
    .A(\system_expander.i2cCtrl_io_cmd_payload_data[4] ));
 sg13g2_a21oi_1 _0637_ (.A1(\system_expander.link_regAddr[3] ),
    .A2(_0137_),
    .Y(_0154_),
    .B1(net294));
 sg13g2_nor3_1 _0638_ (.A(\system_expander.link_regAddr[4] ),
    .B(_0112_),
    .C(_0154_),
    .Y(_0155_));
 sg13g2_a21oi_1 _0639_ (.A1(\system_expander.link_regAddr[4] ),
    .A2(_0150_),
    .Y(_0156_),
    .B1(_0155_));
 sg13g2_a21oi_1 _0640_ (.A1(_0153_),
    .A2(_0133_),
    .Y(_0101_),
    .B1(_0156_));
 sg13g2_inv_1 _0642_ (.Y(_0158_),
    .A(\system_expander.link_regAddr[5] ));
 sg13g2_and3_1 _0643_ (.X(_0159_),
    .A(\system_expander.link_regAddr[3] ),
    .B(\system_expander.link_regAddr[4] ),
    .C(_0137_));
 sg13g2_o21ai_1 _0644_ (.B1(\system_expander.i2cCtrl_io_cmd_ready ),
    .Y(_0160_),
    .A1(net294),
    .A2(_0159_));
 sg13g2_nand3_1 _0646_ (.B(_0110_),
    .C(_0159_),
    .A(\system_expander.link_regAddr[5] ),
    .Y(_0162_));
 sg13g2_o21ai_1 _0647_ (.B1(_0162_),
    .Y(_0163_),
    .A1(\system_expander.i2cCtrl_io_cmd_payload_data[5] ),
    .A2(_0143_));
 sg13g2_a21oi_1 _0648_ (.A1(_0158_),
    .A2(_0160_),
    .Y(_0102_),
    .B1(_0163_));
 sg13g2_a21o_1 _0649_ (.A2(_0159_),
    .A1(\system_expander.link_regAddr[5] ),
    .B1(net294),
    .X(_0164_));
 sg13g2_a21oi_1 _0650_ (.A1(\system_expander.i2cCtrl_io_cmd_ready ),
    .A2(_0164_),
    .Y(_0165_),
    .B1(\system_expander.link_regAddr[6] ));
 sg13g2_nand3_1 _0651_ (.B(\system_expander.link_regAddr[6] ),
    .C(_0159_),
    .A(\system_expander.link_regAddr[5] ),
    .Y(_0166_));
 sg13g2_nor2_1 _0652_ (.A(net294),
    .B(_0166_),
    .Y(_0167_));
 sg13g2_nor2_1 _0654_ (.A(\system_expander.i2cCtrl_io_cmd_payload_data[6] ),
    .B(_0143_),
    .Y(_0169_));
 sg13g2_nor3_1 _0655_ (.A(_0165_),
    .B(_0167_),
    .C(_0169_),
    .Y(_0103_));
 sg13g2_inv_1 _0657_ (.Y(_0171_),
    .A(\system_expander.i2cCtrl_io_cmd_payload_data[7] ));
 sg13g2_a21oi_1 _0658_ (.A1(_0110_),
    .A2(_0166_),
    .Y(_0172_),
    .B1(_0112_));
 sg13g2_nor2_1 _0659_ (.A(\system_expander.link_regAddr[7] ),
    .B(_0172_),
    .Y(_0173_));
 sg13g2_a221oi_1 _0660_ (.B2(\system_expander.link_regAddr[7] ),
    .C1(_0173_),
    .B1(_0167_),
    .A1(_0171_),
    .Y(_0104_),
    .A2(_0133_));
 sg13g2_mux2_1 _0661_ (.A0(sg13g2_IOPad_io_address_0_p2c),
    .A1(\system_expander.i2cConfig_latchedAddress[0] ),
    .S(\system_expander.i2cConfig_latch ),
    .X(_0021_));
 sg13g2_mux2_1 _0662_ (.A0(sg13g2_IOPad_io_address_1_p2c),
    .A1(\system_expander.i2cConfig_latchedAddress[1] ),
    .S(\system_expander.i2cConfig_latch ),
    .X(_0022_));
 sg13g2_mux2_1 _0663_ (.A0(sg13g2_IOPad_io_address_2_p2c),
    .A1(\system_expander.i2cConfig_latchedAddress[2] ),
    .S(\system_expander.i2cConfig_latch ),
    .X(_0023_));
 sg13g2_or4_2 _0664_ (.A(\system_expander.link_regAddr[5] ),
    .B(\system_expander.link_regAddr[4] ),
    .C(\system_expander.link_regAddr[7] ),
    .D(\system_expander.link_regAddr[6] ),
    .X(_0174_));
 sg13g2_nor3_2 _0666_ (.A(net301),
    .B(net302),
    .C(_0174_),
    .Y(_0176_));
 sg13g2_nor2b_1 _0667_ (.A(net306),
    .B_N(net303),
    .Y(_0177_));
 sg13g2_and3_1 _0668_ (.X(_0178_),
    .A(net299),
    .B(_0176_),
    .C(_0177_));
 sg13g2_nand2_1 _0671_ (.Y(_0181_),
    .A(net315),
    .B(net289));
 sg13g2_nand2b_1 _0672_ (.Y(_0182_),
    .B(sg13g2_IOPad_io_gpio_0_c2p_en),
    .A_N(net289));
 sg13g2_a21oi_1 _0673_ (.A1(_0181_),
    .A2(_0182_),
    .Y(_0005_),
    .B1(net320));
 sg13g2_nand2_1 _0674_ (.Y(_0183_),
    .A(net314),
    .B(net290));
 sg13g2_nand2b_1 _0675_ (.Y(_0184_),
    .B(sg13g2_IOPad_io_gpio_1_c2p_en),
    .A_N(net290));
 sg13g2_a21oi_1 _0676_ (.A1(_0183_),
    .A2(_0184_),
    .Y(_0006_),
    .B1(net323));
 sg13g2_nand2_1 _0677_ (.Y(_0185_),
    .A(net313),
    .B(net290));
 sg13g2_nand2b_1 _0678_ (.Y(_0186_),
    .B(sg13g2_IOPad_io_gpio_2_c2p_en),
    .A_N(net290));
 sg13g2_a21oi_1 _0679_ (.A1(_0185_),
    .A2(_0186_),
    .Y(_0007_),
    .B1(net324));
 sg13g2_nand2_1 _0680_ (.Y(_0187_),
    .A(\system_expander.i2cCtrl_io_cmd_payload_data[3] ),
    .B(net290));
 sg13g2_nand2b_1 _0681_ (.Y(_0188_),
    .B(sg13g2_IOPad_io_gpio_3_c2p_en),
    .A_N(net290));
 sg13g2_a21oi_1 _0682_ (.A1(_0187_),
    .A2(_0188_),
    .Y(_0008_),
    .B1(net324));
 sg13g2_nand2_1 _0683_ (.Y(_0189_),
    .A(net311),
    .B(net290));
 sg13g2_nand2b_1 _0684_ (.Y(_0190_),
    .B(sg13g2_IOPad_io_gpio_4_c2p_en),
    .A_N(net290));
 sg13g2_a21oi_1 _0685_ (.A1(_0189_),
    .A2(_0190_),
    .Y(_0009_),
    .B1(net324));
 sg13g2_nand2_1 _0686_ (.Y(_0191_),
    .A(net310),
    .B(net289));
 sg13g2_nand2b_1 _0687_ (.Y(_0192_),
    .B(sg13g2_IOPad_io_gpio_5_c2p_en),
    .A_N(net289));
 sg13g2_a21oi_1 _0689_ (.A1(_0191_),
    .A2(_0192_),
    .Y(_0010_),
    .B1(net316));
 sg13g2_nand2_1 _0690_ (.Y(_0194_),
    .A(net309),
    .B(net289));
 sg13g2_nand2b_1 _0691_ (.Y(_0195_),
    .B(sg13g2_IOPad_io_gpio_6_c2p_en),
    .A_N(net289));
 sg13g2_a21oi_1 _0692_ (.A1(_0194_),
    .A2(_0195_),
    .Y(_0011_),
    .B1(net316));
 sg13g2_nand2_1 _0693_ (.Y(_0196_),
    .A(net308),
    .B(net289));
 sg13g2_nand2b_1 _0694_ (.Y(_0197_),
    .B(sg13g2_IOPad_io_gpio_7_c2p_en),
    .A_N(net289));
 sg13g2_a21oi_1 _0695_ (.A1(_0196_),
    .A2(_0197_),
    .Y(_0012_),
    .B1(net317));
 sg13g2_and3_1 _0696_ (.X(_0198_),
    .A(net299),
    .B(_0134_),
    .C(_0176_));
 sg13g2_nand2_1 _0699_ (.Y(_0201_),
    .A(net315),
    .B(_0198_));
 sg13g2_nand2b_1 _0700_ (.Y(_0202_),
    .B(sg13g2_IOPad_io_gpio_0_c2p),
    .A_N(_0198_));
 sg13g2_a21oi_1 _0701_ (.A1(_0201_),
    .A2(_0202_),
    .Y(_0013_),
    .B1(net320));
 sg13g2_nand2_1 _0702_ (.Y(_0203_),
    .A(net314),
    .B(_0198_));
 sg13g2_nand2b_1 _0703_ (.Y(_0204_),
    .B(sg13g2_IOPad_io_gpio_1_c2p),
    .A_N(_0198_));
 sg13g2_a21oi_1 _0704_ (.A1(_0203_),
    .A2(_0204_),
    .Y(_0014_),
    .B1(net323));
 sg13g2_nand2_1 _0705_ (.Y(_0205_),
    .A(net313),
    .B(net288));
 sg13g2_nand2b_1 _0706_ (.Y(_0206_),
    .B(sg13g2_IOPad_io_gpio_2_c2p),
    .A_N(net288));
 sg13g2_a21oi_1 _0707_ (.A1(_0205_),
    .A2(_0206_),
    .Y(_0015_),
    .B1(net324));
 sg13g2_nand2_1 _0708_ (.Y(_0207_),
    .A(\system_expander.i2cCtrl_io_cmd_payload_data[3] ),
    .B(net288));
 sg13g2_nand2b_1 _0709_ (.Y(_0208_),
    .B(sg13g2_IOPad_io_gpio_3_c2p),
    .A_N(net288));
 sg13g2_a21oi_1 _0710_ (.A1(_0207_),
    .A2(_0208_),
    .Y(_0016_),
    .B1(net324));
 sg13g2_nand2_1 _0711_ (.Y(_0209_),
    .A(net311),
    .B(net288));
 sg13g2_nand2b_1 _0712_ (.Y(_0210_),
    .B(sg13g2_IOPad_io_gpio_4_c2p),
    .A_N(net288));
 sg13g2_a21oi_1 _0713_ (.A1(_0209_),
    .A2(_0210_),
    .Y(_0017_),
    .B1(net324));
 sg13g2_nand2_1 _0714_ (.Y(_0211_),
    .A(net310),
    .B(net287));
 sg13g2_nand2b_1 _0715_ (.Y(_0212_),
    .B(sg13g2_IOPad_io_gpio_5_c2p),
    .A_N(net287));
 sg13g2_a21oi_1 _0716_ (.A1(_0211_),
    .A2(_0212_),
    .Y(_0018_),
    .B1(net316));
 sg13g2_nand2_1 _0717_ (.Y(_0213_),
    .A(net309),
    .B(net287));
 sg13g2_nand2b_1 _0718_ (.Y(_0214_),
    .B(sg13g2_IOPad_io_gpio_6_c2p),
    .A_N(net287));
 sg13g2_a21oi_1 _0719_ (.A1(_0213_),
    .A2(_0214_),
    .Y(_0019_),
    .B1(net316));
 sg13g2_nand2_1 _0720_ (.Y(_0215_),
    .A(net308),
    .B(net287));
 sg13g2_nand2b_1 _0721_ (.Y(_0216_),
    .B(sg13g2_IOPad_io_gpio_7_c2p),
    .A_N(net287));
 sg13g2_a21oi_1 _0723_ (.A1(_0215_),
    .A2(_0216_),
    .Y(_0020_),
    .B1(net317));
 sg13g2_inv_1 _0725_ (.Y(_0219_),
    .A(\system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[0] ));
 sg13g2_nor3_2 _0729_ (.A(\system_expander.link_regAddr[3] ),
    .B(_0141_),
    .C(_0174_),
    .Y(_0223_));
 sg13g2_and2_1 _0730_ (.A(_0177_),
    .B(_0223_),
    .X(_0224_));
 sg13g2_nand3_1 _0732_ (.B(net315),
    .C(_0224_),
    .A(net299),
    .Y(_0226_));
 sg13g2_a22oi_1 _0733_ (.Y(_0227_),
    .B1(_0226_),
    .B2(\system_expander.irq_fall_ctrl.pendings[0] ),
    .A2(_0219_),
    .A1(\system_expander.gpioCtrl_1.last[0] ));
 sg13g2_nor2_1 _0734_ (.A(net319),
    .B(_0227_),
    .Y(_0024_));
 sg13g2_inv_1 _0735_ (.Y(_0228_),
    .A(\system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[1] ));
 sg13g2_nand3_1 _0736_ (.B(net314),
    .C(_0224_),
    .A(net299),
    .Y(_0229_));
 sg13g2_a22oi_1 _0737_ (.Y(_0230_),
    .B1(_0229_),
    .B2(\system_expander.irq_fall_ctrl.pendings[1] ),
    .A2(_0228_),
    .A1(\system_expander.gpioCtrl_1.last[1] ));
 sg13g2_nor2_1 _0738_ (.A(net323),
    .B(_0230_),
    .Y(_0025_));
 sg13g2_inv_1 _0739_ (.Y(_0231_),
    .A(\system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[2] ));
 sg13g2_nand3_1 _0740_ (.B(net313),
    .C(_0224_),
    .A(net295),
    .Y(_0232_));
 sg13g2_a22oi_1 _0741_ (.Y(_0233_),
    .B1(_0232_),
    .B2(\system_expander.irq_fall_ctrl.pendings[2] ),
    .A2(_0231_),
    .A1(\system_expander.gpioCtrl_1.last[2] ));
 sg13g2_nor2_1 _0742_ (.A(net326),
    .B(_0233_),
    .Y(_0026_));
 sg13g2_inv_1 _0743_ (.Y(_0234_),
    .A(\system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[3] ));
 sg13g2_nand3_1 _0744_ (.B(\system_expander.i2cCtrl_io_cmd_payload_data[3] ),
    .C(_0224_),
    .A(net295),
    .Y(_0235_));
 sg13g2_a22oi_1 _0745_ (.Y(_0236_),
    .B1(_0235_),
    .B2(\system_expander.irq_fall_ctrl.pendings[3] ),
    .A2(_0234_),
    .A1(\system_expander.gpioCtrl_1.last[3] ));
 sg13g2_nor2_1 _0746_ (.A(net326),
    .B(_0236_),
    .Y(_0027_));
 sg13g2_inv_1 _0747_ (.Y(_0237_),
    .A(\system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[4] ));
 sg13g2_nand3_1 _0748_ (.B(net311),
    .C(_0224_),
    .A(net295),
    .Y(_0238_));
 sg13g2_a22oi_1 _0749_ (.Y(_0239_),
    .B1(_0238_),
    .B2(\system_expander.irq_fall_ctrl.pendings[4] ),
    .A2(_0237_),
    .A1(\system_expander.gpioCtrl_1.last[4] ));
 sg13g2_nor2_1 _0750_ (.A(net324),
    .B(_0239_),
    .Y(_0028_));
 sg13g2_inv_1 _0751_ (.Y(_0240_),
    .A(\system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[5] ));
 sg13g2_nand3_1 _0752_ (.B(net310),
    .C(net286),
    .A(net297),
    .Y(_0241_));
 sg13g2_a22oi_1 _0753_ (.Y(_0242_),
    .B1(_0241_),
    .B2(\system_expander.irq_fall_ctrl.pendings[5] ),
    .A2(_0240_),
    .A1(\system_expander.gpioCtrl_1.last[5] ));
 sg13g2_nor2_1 _0754_ (.A(net321),
    .B(_0242_),
    .Y(_0029_));
 sg13g2_inv_1 _0755_ (.Y(_0243_),
    .A(\system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[6] ));
 sg13g2_nand3_1 _0756_ (.B(net309),
    .C(net286),
    .A(net297),
    .Y(_0244_));
 sg13g2_a22oi_1 _0757_ (.Y(_0245_),
    .B1(_0244_),
    .B2(\system_expander.irq_fall_ctrl.pendings[6] ),
    .A2(_0243_),
    .A1(\system_expander.gpioCtrl_1.last[6] ));
 sg13g2_nor2_1 _0758_ (.A(net316),
    .B(_0245_),
    .Y(_0030_));
 sg13g2_inv_1 _0759_ (.Y(_0246_),
    .A(\system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[7] ));
 sg13g2_nand3_1 _0760_ (.B(net308),
    .C(net286),
    .A(net297),
    .Y(_0247_));
 sg13g2_a22oi_1 _0761_ (.Y(_0248_),
    .B1(_0247_),
    .B2(\system_expander.irq_fall_ctrl.pendings[7] ),
    .A2(_0246_),
    .A1(\system_expander.gpioCtrl_1.last[7] ));
 sg13g2_nor2_1 _0762_ (.A(net318),
    .B(_0248_),
    .Y(_0031_));
 sg13g2_nor3_2 _0763_ (.A(_0145_),
    .B(net302),
    .C(_0174_),
    .Y(_0249_));
 sg13g2_and3_1 _0764_ (.X(_0250_),
    .A(net299),
    .B(_0177_),
    .C(_0249_));
 sg13g2_nand2_1 _0767_ (.Y(_0253_),
    .A(net315),
    .B(net284));
 sg13g2_nand2b_1 _0768_ (.Y(_0254_),
    .B(\system_expander.irq_fall_ctrl.io_masks[0] ),
    .A_N(net284));
 sg13g2_a21oi_1 _0769_ (.A1(_0253_),
    .A2(_0254_),
    .Y(_0032_),
    .B1(net320));
 sg13g2_nand2_1 _0770_ (.Y(_0255_),
    .A(net314),
    .B(net285));
 sg13g2_nand2b_1 _0771_ (.Y(_0256_),
    .B(\system_expander.irq_fall_ctrl.io_masks[1] ),
    .A_N(net285));
 sg13g2_a21oi_1 _0772_ (.A1(_0255_),
    .A2(_0256_),
    .Y(_0033_),
    .B1(net327));
 sg13g2_nand2_1 _0773_ (.Y(_0257_),
    .A(net313),
    .B(net285));
 sg13g2_nand2b_1 _0774_ (.Y(_0258_),
    .B(\system_expander.irq_fall_ctrl.io_masks[2] ),
    .A_N(net285));
 sg13g2_a21oi_1 _0775_ (.A1(_0257_),
    .A2(_0258_),
    .Y(_0034_),
    .B1(net325));
 sg13g2_nand2_1 _0776_ (.Y(_0259_),
    .A(net312),
    .B(net285));
 sg13g2_nand2b_1 _0777_ (.Y(_0260_),
    .B(\system_expander.irq_fall_ctrl.io_masks[3] ),
    .A_N(net285));
 sg13g2_a21oi_1 _0778_ (.A1(_0259_),
    .A2(_0260_),
    .Y(_0035_),
    .B1(net326));
 sg13g2_nand2_1 _0779_ (.Y(_0261_),
    .A(net311),
    .B(net285));
 sg13g2_nand2b_1 _0780_ (.Y(_0262_),
    .B(\system_expander.irq_fall_ctrl.io_masks[4] ),
    .A_N(net285));
 sg13g2_a21oi_1 _0781_ (.A1(_0261_),
    .A2(_0262_),
    .Y(_0036_),
    .B1(net325));
 sg13g2_nand2_1 _0782_ (.Y(_0263_),
    .A(net310),
    .B(net284));
 sg13g2_nand2b_1 _0783_ (.Y(_0264_),
    .B(\system_expander.irq_fall_ctrl.io_masks[5] ),
    .A_N(net284));
 sg13g2_a21oi_1 _0784_ (.A1(_0263_),
    .A2(_0264_),
    .Y(_0037_),
    .B1(net316));
 sg13g2_nand2_1 _0785_ (.Y(_0265_),
    .A(net309),
    .B(net284));
 sg13g2_nand2b_1 _0786_ (.Y(_0266_),
    .B(\system_expander.irq_fall_ctrl.io_masks[6] ),
    .A_N(net284));
 sg13g2_a21oi_1 _0787_ (.A1(_0265_),
    .A2(_0266_),
    .Y(_0038_),
    .B1(net316));
 sg13g2_nand2_1 _0788_ (.Y(_0267_),
    .A(net308),
    .B(net284));
 sg13g2_nand2b_1 _0789_ (.Y(_0268_),
    .B(\system_expander.irq_fall_ctrl.io_masks[7] ),
    .A_N(net284));
 sg13g2_a21oi_1 _0790_ (.A1(_0267_),
    .A2(_0268_),
    .Y(_0039_),
    .B1(net317));
 sg13g2_nand2_1 _0791_ (.Y(_0269_),
    .A(net299),
    .B(net315));
 sg13g2_and2_1 _0792_ (.A(_0139_),
    .B(_0176_),
    .X(_0270_));
 sg13g2_nand2b_1 _0794_ (.Y(_0272_),
    .B(_0270_),
    .A_N(_0269_));
 sg13g2_a21oi_1 _0795_ (.A1(\system_expander.irq_high_ctrl.pendings[0] ),
    .A2(_0272_),
    .Y(_0273_),
    .B1(\system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[0] ));
 sg13g2_nor2_1 _0796_ (.A(net319),
    .B(_0273_),
    .Y(_0040_));
 sg13g2_nand2_1 _0797_ (.Y(_0274_),
    .A(net299),
    .B(net314));
 sg13g2_nand2b_1 _0798_ (.Y(_0275_),
    .B(net283),
    .A_N(_0274_));
 sg13g2_a21oi_1 _0799_ (.A1(\system_expander.irq_high_ctrl.pendings[1] ),
    .A2(_0275_),
    .Y(_0276_),
    .B1(\system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[1] ));
 sg13g2_nor2_1 _0800_ (.A(net323),
    .B(_0276_),
    .Y(_0041_));
 sg13g2_nand2_1 _0802_ (.Y(_0278_),
    .A(net295),
    .B(net313));
 sg13g2_nand2b_1 _0803_ (.Y(_0279_),
    .B(net283),
    .A_N(_0278_));
 sg13g2_a21oi_1 _0804_ (.A1(\system_expander.irq_high_ctrl.pendings[2] ),
    .A2(_0279_),
    .Y(_0280_),
    .B1(\system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[2] ));
 sg13g2_nor2_1 _0805_ (.A(net325),
    .B(_0280_),
    .Y(_0042_));
 sg13g2_nand2_1 _0806_ (.Y(_0281_),
    .A(net295),
    .B(\system_expander.i2cCtrl_io_cmd_payload_data[3] ));
 sg13g2_nand2b_1 _0807_ (.Y(_0282_),
    .B(net283),
    .A_N(_0281_));
 sg13g2_a21oi_1 _0808_ (.A1(\system_expander.irq_high_ctrl.pendings[3] ),
    .A2(_0282_),
    .Y(_0283_),
    .B1(\system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[3] ));
 sg13g2_nor2_1 _0809_ (.A(net325),
    .B(_0283_),
    .Y(_0043_));
 sg13g2_nand2_1 _0810_ (.Y(_0284_),
    .A(net295),
    .B(net311));
 sg13g2_nand2b_1 _0811_ (.Y(_0285_),
    .B(net283),
    .A_N(_0284_));
 sg13g2_a21oi_1 _0812_ (.A1(\system_expander.irq_high_ctrl.pendings[4] ),
    .A2(_0285_),
    .Y(_0286_),
    .B1(\system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[4] ));
 sg13g2_nor2_1 _0813_ (.A(net322),
    .B(_0286_),
    .Y(_0044_));
 sg13g2_nand2_1 _0814_ (.Y(_0287_),
    .A(net297),
    .B(net310));
 sg13g2_nand2b_1 _0815_ (.Y(_0288_),
    .B(_0270_),
    .A_N(_0287_));
 sg13g2_a21oi_1 _0816_ (.A1(\system_expander.irq_high_ctrl.pendings[5] ),
    .A2(_0288_),
    .Y(_0289_),
    .B1(\system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[5] ));
 sg13g2_nor2_1 _0817_ (.A(net320),
    .B(_0289_),
    .Y(_0045_));
 sg13g2_nand2_1 _0818_ (.Y(_0290_),
    .A(net297),
    .B(net309));
 sg13g2_nand2b_1 _0819_ (.Y(_0291_),
    .B(_0270_),
    .A_N(_0290_));
 sg13g2_a21oi_1 _0820_ (.A1(\system_expander.irq_high_ctrl.pendings[6] ),
    .A2(_0291_),
    .Y(_0292_),
    .B1(\system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[6] ));
 sg13g2_nor2_1 _0821_ (.A(net317),
    .B(_0292_),
    .Y(_0046_));
 sg13g2_nand2_1 _0822_ (.Y(_0293_),
    .A(net297),
    .B(net308));
 sg13g2_nand2b_1 _0823_ (.Y(_0294_),
    .B(_0270_),
    .A_N(_0293_));
 sg13g2_a21oi_1 _0824_ (.A1(\system_expander.irq_high_ctrl.pendings[7] ),
    .A2(_0294_),
    .Y(_0295_),
    .B1(\system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[7] ));
 sg13g2_nor2_1 _0825_ (.A(net317),
    .B(_0295_),
    .Y(_0047_));
 sg13g2_and3_1 _0826_ (.X(_0296_),
    .A(net299),
    .B(_0139_),
    .C(net292));
 sg13g2_nand2_1 _0829_ (.Y(_0299_),
    .A(net315),
    .B(net281));
 sg13g2_nand2b_1 _0830_ (.Y(_0300_),
    .B(\system_expander.irq_high_ctrl.io_masks[0] ),
    .A_N(net281));
 sg13g2_a21oi_1 _0831_ (.A1(_0299_),
    .A2(_0300_),
    .Y(_0048_),
    .B1(net319));
 sg13g2_nand2_1 _0832_ (.Y(_0301_),
    .A(net314),
    .B(net282));
 sg13g2_nand2b_1 _0833_ (.Y(_0302_),
    .B(\system_expander.irq_high_ctrl.io_masks[1] ),
    .A_N(net282));
 sg13g2_a21oi_1 _0835_ (.A1(_0301_),
    .A2(_0302_),
    .Y(_0049_),
    .B1(net323));
 sg13g2_nand2_1 _0836_ (.Y(_0304_),
    .A(net313),
    .B(net282));
 sg13g2_nand2b_1 _0837_ (.Y(_0305_),
    .B(\system_expander.irq_high_ctrl.io_masks[2] ),
    .A_N(net282));
 sg13g2_a21oi_1 _0838_ (.A1(_0304_),
    .A2(_0305_),
    .Y(_0050_),
    .B1(net325));
 sg13g2_nand2_1 _0839_ (.Y(_0306_),
    .A(net312),
    .B(net282));
 sg13g2_nand2b_1 _0840_ (.Y(_0307_),
    .B(\system_expander.irq_high_ctrl.io_masks[3] ),
    .A_N(net282));
 sg13g2_a21oi_1 _0841_ (.A1(_0306_),
    .A2(_0307_),
    .Y(_0051_),
    .B1(net325));
 sg13g2_nand2_1 _0842_ (.Y(_0308_),
    .A(net311),
    .B(net282));
 sg13g2_nand2b_1 _0843_ (.Y(_0309_),
    .B(\system_expander.irq_high_ctrl.io_masks[4] ),
    .A_N(net282));
 sg13g2_a21oi_1 _0844_ (.A1(_0308_),
    .A2(_0309_),
    .Y(_0052_),
    .B1(net324));
 sg13g2_nand2_1 _0845_ (.Y(_0310_),
    .A(\system_expander.i2cCtrl_io_cmd_payload_data[5] ),
    .B(net281));
 sg13g2_nand2b_1 _0846_ (.Y(_0311_),
    .B(\system_expander.irq_high_ctrl.io_masks[5] ),
    .A_N(net281));
 sg13g2_a21oi_1 _0847_ (.A1(_0310_),
    .A2(_0311_),
    .Y(_0053_),
    .B1(net318));
 sg13g2_nand2_1 _0848_ (.Y(_0312_),
    .A(net309),
    .B(net281));
 sg13g2_nand2b_1 _0849_ (.Y(_0313_),
    .B(\system_expander.irq_high_ctrl.io_masks[6] ),
    .A_N(net281));
 sg13g2_a21oi_1 _0850_ (.A1(_0312_),
    .A2(_0313_),
    .Y(_0054_),
    .B1(net318));
 sg13g2_nand2_1 _0851_ (.Y(_0314_),
    .A(net308),
    .B(net281));
 sg13g2_nand2b_1 _0852_ (.Y(_0315_),
    .B(\system_expander.irq_high_ctrl.io_masks[7] ),
    .A_N(net281));
 sg13g2_a21oi_1 _0853_ (.A1(_0314_),
    .A2(_0315_),
    .Y(_0055_),
    .B1(net318));
 sg13g2_nor2_1 _0854_ (.A(net307),
    .B(\system_expander.link_regAddr[1] ),
    .Y(_0316_));
 sg13g2_nand2_2 _0855_ (.Y(_0317_),
    .A(net292),
    .B(_0316_));
 sg13g2_o21ai_1 _0856_ (.B1(\system_expander.irq_low_ctrl.pendings[0] ),
    .Y(_0318_),
    .A1(_0269_),
    .A2(_0317_));
 sg13g2_a21oi_1 _0857_ (.A1(\system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[0] ),
    .A2(_0318_),
    .Y(_0056_),
    .B1(net319));
 sg13g2_o21ai_1 _0858_ (.B1(\system_expander.irq_low_ctrl.pendings[1] ),
    .Y(_0319_),
    .A1(_0274_),
    .A2(_0317_));
 sg13g2_a21oi_1 _0859_ (.A1(\system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[1] ),
    .A2(_0319_),
    .Y(_0057_),
    .B1(net323));
 sg13g2_o21ai_1 _0860_ (.B1(\system_expander.irq_low_ctrl.pendings[2] ),
    .Y(_0320_),
    .A1(_0278_),
    .A2(_0317_));
 sg13g2_a21oi_1 _0861_ (.A1(\system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[2] ),
    .A2(_0320_),
    .Y(_0058_),
    .B1(net326));
 sg13g2_o21ai_1 _0862_ (.B1(\system_expander.irq_low_ctrl.pendings[3] ),
    .Y(_0321_),
    .A1(_0281_),
    .A2(_0317_));
 sg13g2_a21oi_1 _0864_ (.A1(\system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[3] ),
    .A2(_0321_),
    .Y(_0059_),
    .B1(net322));
 sg13g2_o21ai_1 _0865_ (.B1(\system_expander.irq_low_ctrl.pendings[4] ),
    .Y(_0323_),
    .A1(_0284_),
    .A2(_0317_));
 sg13g2_a21oi_1 _0866_ (.A1(\system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[4] ),
    .A2(_0323_),
    .Y(_0060_),
    .B1(net322));
 sg13g2_o21ai_1 _0867_ (.B1(\system_expander.irq_low_ctrl.pendings[5] ),
    .Y(_0324_),
    .A1(_0287_),
    .A2(_0317_));
 sg13g2_a21oi_1 _0868_ (.A1(\system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[5] ),
    .A2(_0324_),
    .Y(_0061_),
    .B1(net321));
 sg13g2_o21ai_1 _0869_ (.B1(\system_expander.irq_low_ctrl.pendings[6] ),
    .Y(_0325_),
    .A1(_0290_),
    .A2(_0317_));
 sg13g2_a21oi_1 _0870_ (.A1(\system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[6] ),
    .A2(_0325_),
    .Y(_0062_),
    .B1(net317));
 sg13g2_o21ai_1 _0871_ (.B1(\system_expander.irq_low_ctrl.pendings[7] ),
    .Y(_0326_),
    .A1(_0293_),
    .A2(_0317_));
 sg13g2_a21oi_1 _0872_ (.A1(\system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[7] ),
    .A2(_0326_),
    .Y(_0063_),
    .B1(net317));
 sg13g2_nor4_2 _0873_ (.A(\system_expander.link_regAddr[5] ),
    .B(\system_expander.link_regAddr[4] ),
    .C(\system_expander.link_regAddr[7] ),
    .Y(_0327_),
    .D(\system_expander.link_regAddr[6] ));
 sg13g2_nand2_2 _0874_ (.Y(_0328_),
    .A(_0141_),
    .B(_0327_));
 sg13g2_nor4_2 _0875_ (.A(net306),
    .B(\system_expander.link_regAddr[1] ),
    .C(_0145_),
    .Y(_0329_),
    .D(_0328_));
 sg13g2_nand3_1 _0877_ (.B(net315),
    .C(_0329_),
    .A(net298),
    .Y(_0331_));
 sg13g2_nand2_2 _0878_ (.Y(_0332_),
    .A(net296),
    .B(net280));
 sg13g2_nand2_1 _0879_ (.Y(_0333_),
    .A(\system_expander.irq_low_ctrl.io_masks[0] ),
    .B(_0332_));
 sg13g2_a21oi_1 _0880_ (.A1(_0331_),
    .A2(_0333_),
    .Y(_0064_),
    .B1(net328));
 sg13g2_nand3_1 _0881_ (.B(net314),
    .C(net280),
    .A(net298),
    .Y(_0334_));
 sg13g2_nand2_1 _0882_ (.Y(_0335_),
    .A(\system_expander.irq_low_ctrl.io_masks[1] ),
    .B(_0332_));
 sg13g2_a21oi_1 _0883_ (.A1(_0334_),
    .A2(_0335_),
    .Y(_0065_),
    .B1(net322));
 sg13g2_nand3_1 _0884_ (.B(net313),
    .C(net280),
    .A(net296),
    .Y(_0336_));
 sg13g2_nand2_1 _0885_ (.Y(_0337_),
    .A(\system_expander.irq_low_ctrl.io_masks[2] ),
    .B(_0332_));
 sg13g2_a21oi_1 _0886_ (.A1(_0336_),
    .A2(_0337_),
    .Y(_0066_),
    .B1(net322));
 sg13g2_nand3_1 _0887_ (.B(net312),
    .C(net280),
    .A(net296),
    .Y(_0338_));
 sg13g2_nand2_1 _0888_ (.Y(_0339_),
    .A(\system_expander.irq_low_ctrl.io_masks[3] ),
    .B(_0332_));
 sg13g2_a21oi_1 _0889_ (.A1(_0338_),
    .A2(_0339_),
    .Y(_0067_),
    .B1(net322));
 sg13g2_nand3_1 _0890_ (.B(net311),
    .C(net280),
    .A(net296),
    .Y(_0340_));
 sg13g2_nand2_1 _0891_ (.Y(_0341_),
    .A(\system_expander.irq_low_ctrl.io_masks[4] ),
    .B(_0332_));
 sg13g2_a21oi_1 _0892_ (.A1(_0340_),
    .A2(_0341_),
    .Y(_0068_),
    .B1(net322));
 sg13g2_nand3_1 _0893_ (.B(\system_expander.i2cCtrl_io_cmd_payload_data[5] ),
    .C(_0329_),
    .A(net297),
    .Y(_0342_));
 sg13g2_nand2_1 _0894_ (.Y(_0343_),
    .A(\system_expander.irq_low_ctrl.io_masks[5] ),
    .B(_0332_));
 sg13g2_a21oi_1 _0896_ (.A1(_0342_),
    .A2(_0343_),
    .Y(_0069_),
    .B1(net328));
 sg13g2_nand3_1 _0897_ (.B(net309),
    .C(_0329_),
    .A(net298),
    .Y(_0345_));
 sg13g2_nand2_1 _0898_ (.Y(_0346_),
    .A(\system_expander.irq_low_ctrl.io_masks[6] ),
    .B(_0332_));
 sg13g2_a21oi_1 _0899_ (.A1(_0345_),
    .A2(_0346_),
    .Y(_0070_),
    .B1(net328));
 sg13g2_nand3_1 _0900_ (.B(net308),
    .C(_0329_),
    .A(net298),
    .Y(_0347_));
 sg13g2_nand2_1 _0901_ (.Y(_0348_),
    .A(\system_expander.irq_low_ctrl.io_masks[7] ),
    .B(_0332_));
 sg13g2_a21oi_1 _0902_ (.A1(_0347_),
    .A2(_0348_),
    .Y(_0071_),
    .B1(net328));
 sg13g2_inv_1 _0903_ (.Y(_0349_),
    .A(\system_expander.gpioCtrl_1.last[0] ));
 sg13g2_nand2b_1 _0904_ (.Y(_0350_),
    .B(net306),
    .A_N(net305));
 sg13g2_nand3_1 _0905_ (.B(\system_expander.link_regAddr[2] ),
    .C(_0327_),
    .A(_0145_),
    .Y(_0351_));
 sg13g2_nor2_1 _0907_ (.A(_0350_),
    .B(_0351_),
    .Y(_0353_));
 sg13g2_nand2b_1 _0909_ (.Y(_0355_),
    .B(net279),
    .A_N(_0269_));
 sg13g2_a22oi_1 _0910_ (.Y(_0356_),
    .B1(\system_expander.irq_rise_ctrl.pendings[0] ),
    .B2(_0355_),
    .A2(\system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[0] ),
    .A1(_0349_));
 sg13g2_nor2_1 _0911_ (.A(net319),
    .B(_0356_),
    .Y(_0072_));
 sg13g2_inv_1 _0912_ (.Y(_0357_),
    .A(\system_expander.gpioCtrl_1.last[1] ));
 sg13g2_nand2b_1 _0913_ (.Y(_0358_),
    .B(net279),
    .A_N(_0274_));
 sg13g2_a22oi_1 _0914_ (.Y(_0359_),
    .B1(\system_expander.irq_rise_ctrl.pendings[1] ),
    .B2(_0358_),
    .A2(\system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[1] ),
    .A1(_0357_));
 sg13g2_nor2_1 _0915_ (.A(net323),
    .B(_0359_),
    .Y(_0073_));
 sg13g2_inv_1 _0916_ (.Y(_0360_),
    .A(\system_expander.gpioCtrl_1.last[2] ));
 sg13g2_nand2b_1 _0917_ (.Y(_0361_),
    .B(_0353_),
    .A_N(_0278_));
 sg13g2_a22oi_1 _0918_ (.Y(_0362_),
    .B1(\system_expander.irq_rise_ctrl.pendings[2] ),
    .B2(_0361_),
    .A2(\system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[2] ),
    .A1(_0360_));
 sg13g2_nor2_1 _0919_ (.A(net326),
    .B(_0362_),
    .Y(_0074_));
 sg13g2_inv_1 _0920_ (.Y(_0363_),
    .A(\system_expander.gpioCtrl_1.last[3] ));
 sg13g2_nand2b_1 _0921_ (.Y(_0364_),
    .B(_0353_),
    .A_N(_0281_));
 sg13g2_a22oi_1 _0922_ (.Y(_0365_),
    .B1(\system_expander.irq_rise_ctrl.pendings[3] ),
    .B2(_0364_),
    .A2(\system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[3] ),
    .A1(_0363_));
 sg13g2_nor2_1 _0923_ (.A(net326),
    .B(_0365_),
    .Y(_0075_));
 sg13g2_inv_1 _0924_ (.Y(_0366_),
    .A(\system_expander.gpioCtrl_1.last[4] ));
 sg13g2_nand2b_1 _0925_ (.Y(_0367_),
    .B(_0353_),
    .A_N(_0284_));
 sg13g2_a22oi_1 _0926_ (.Y(_0368_),
    .B1(\system_expander.irq_rise_ctrl.pendings[4] ),
    .B2(_0367_),
    .A2(\system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[4] ),
    .A1(_0366_));
 sg13g2_nor2_1 _0927_ (.A(net327),
    .B(_0368_),
    .Y(_0076_));
 sg13g2_inv_1 _0928_ (.Y(_0369_),
    .A(\system_expander.gpioCtrl_1.last[5] ));
 sg13g2_nand2b_1 _0929_ (.Y(_0370_),
    .B(net279),
    .A_N(_0287_));
 sg13g2_a22oi_1 _0930_ (.Y(_0371_),
    .B1(\system_expander.irq_rise_ctrl.pendings[5] ),
    .B2(_0370_),
    .A2(\system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[5] ),
    .A1(_0369_));
 sg13g2_nor2_1 _0931_ (.A(net321),
    .B(_0371_),
    .Y(_0077_));
 sg13g2_inv_1 _0932_ (.Y(_0372_),
    .A(\system_expander.gpioCtrl_1.last[6] ));
 sg13g2_nand2b_1 _0933_ (.Y(_0373_),
    .B(net279),
    .A_N(_0290_));
 sg13g2_a22oi_1 _0934_ (.Y(_0374_),
    .B1(\system_expander.irq_rise_ctrl.pendings[6] ),
    .B2(_0373_),
    .A2(\system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[6] ),
    .A1(_0372_));
 sg13g2_nor2_1 _0935_ (.A(net316),
    .B(_0374_),
    .Y(_0078_));
 sg13g2_inv_1 _0936_ (.Y(_0375_),
    .A(\system_expander.gpioCtrl_1.last[7] ));
 sg13g2_nand2b_1 _0937_ (.Y(_0376_),
    .B(net279),
    .A_N(_0293_));
 sg13g2_a22oi_1 _0938_ (.Y(_0377_),
    .B1(\system_expander.irq_rise_ctrl.pendings[7] ),
    .B2(_0376_),
    .A2(\system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[7] ),
    .A1(_0375_));
 sg13g2_nor2_1 _0939_ (.A(net318),
    .B(_0377_),
    .Y(_0079_));
 sg13g2_and3_1 _0940_ (.X(_0378_),
    .A(\system_expander.link_state[4] ),
    .B(_0134_),
    .C(_0249_));
 sg13g2_nand2_1 _0943_ (.Y(_0381_),
    .A(net315),
    .B(net277));
 sg13g2_nand2b_1 _0944_ (.Y(_0382_),
    .B(\system_expander.irq_rise_ctrl.io_masks[0] ),
    .A_N(net277));
 sg13g2_a21oi_1 _0945_ (.A1(_0381_),
    .A2(_0382_),
    .Y(_0080_),
    .B1(net319));
 sg13g2_nand2_1 _0946_ (.Y(_0383_),
    .A(net314),
    .B(net278));
 sg13g2_nand2b_1 _0947_ (.Y(_0384_),
    .B(\system_expander.irq_rise_ctrl.io_masks[1] ),
    .A_N(net278));
 sg13g2_a21oi_1 _0948_ (.A1(_0383_),
    .A2(_0384_),
    .Y(_0081_),
    .B1(net323));
 sg13g2_nand2_1 _0949_ (.Y(_0385_),
    .A(net313),
    .B(net278));
 sg13g2_nand2b_1 _0950_ (.Y(_0386_),
    .B(\system_expander.irq_rise_ctrl.io_masks[2] ),
    .A_N(net278));
 sg13g2_a21oi_1 _0951_ (.A1(_0385_),
    .A2(_0386_),
    .Y(_0082_),
    .B1(net326));
 sg13g2_nand2_1 _0952_ (.Y(_0387_),
    .A(net312),
    .B(net278));
 sg13g2_nand2b_1 _0953_ (.Y(_0388_),
    .B(\system_expander.irq_rise_ctrl.io_masks[3] ),
    .A_N(net278));
 sg13g2_a21oi_1 _0954_ (.A1(_0387_),
    .A2(_0388_),
    .Y(_0083_),
    .B1(net326));
 sg13g2_nand2_1 _0955_ (.Y(_0389_),
    .A(net311),
    .B(net278));
 sg13g2_nand2b_1 _0956_ (.Y(_0390_),
    .B(\system_expander.irq_rise_ctrl.io_masks[4] ),
    .A_N(net278));
 sg13g2_a21oi_1 _0957_ (.A1(_0389_),
    .A2(_0390_),
    .Y(_0084_),
    .B1(net322));
 sg13g2_nand2_1 _0958_ (.Y(_0391_),
    .A(net310),
    .B(net277));
 sg13g2_nand2b_1 _0959_ (.Y(_0392_),
    .B(\system_expander.irq_rise_ctrl.io_masks[5] ),
    .A_N(net277));
 sg13g2_a21oi_1 _0960_ (.A1(_0391_),
    .A2(_0392_),
    .Y(_0085_),
    .B1(net321));
 sg13g2_nand2_1 _0961_ (.Y(_0393_),
    .A(net309),
    .B(net277));
 sg13g2_nand2b_1 _0962_ (.Y(_0394_),
    .B(\system_expander.irq_rise_ctrl.io_masks[6] ),
    .A_N(net277));
 sg13g2_a21oi_1 _0963_ (.A1(_0393_),
    .A2(_0394_),
    .Y(_0086_),
    .B1(net321));
 sg13g2_nand2_1 _0964_ (.Y(_0395_),
    .A(net308),
    .B(net277));
 sg13g2_nand2b_1 _0965_ (.Y(_0396_),
    .B(\system_expander.irq_rise_ctrl.io_masks[7] ),
    .A_N(net277));
 sg13g2_a21oi_1 _0966_ (.A1(_0395_),
    .A2(_0396_),
    .Y(_0087_),
    .B1(net318));
 sg13g2_inv_1 _0967_ (.Y(_0397_),
    .A(\system_expander.link_data[0] ));
 sg13g2_nand2_1 _0968_ (.Y(_0398_),
    .A(\system_expander.link_state[2] ),
    .B(_0327_));
 sg13g2_o21ai_1 _0969_ (.B1(net300),
    .Y(_0399_),
    .A1(\system_expander.link_regAddr[2] ),
    .A2(_0139_));
 sg13g2_nand2b_1 _0970_ (.Y(_0400_),
    .B(_0399_),
    .A_N(_0398_));
 sg13g2_nand2_1 _0972_ (.Y(_0402_),
    .A(\system_expander.irq_rise_ctrl.pendings[0] ),
    .B(\system_expander.irq_rise_ctrl.io_masks[0] ));
 sg13g2_nand2_1 _0973_ (.Y(_0403_),
    .A(net303),
    .B(\system_expander.irq_high_ctrl.io_masks[0] ));
 sg13g2_o21ai_1 _0974_ (.B1(_0403_),
    .Y(_0404_),
    .A1(net303),
    .A2(_0402_));
 sg13g2_nor2b_1 _0975_ (.A(net303),
    .B_N(sg13g2_IOPad_io_gpio_0_c2p),
    .Y(_0405_));
 sg13g2_a22oi_1 _0976_ (.Y(_0406_),
    .B1(_0405_),
    .B2(_0176_),
    .A2(_0404_),
    .A1(net292));
 sg13g2_nor2_1 _0977_ (.A(_0122_),
    .B(_0406_),
    .Y(_0407_));
 sg13g2_and2_1 _0978_ (.A(\system_expander.irq_fall_ctrl.pendings[0] ),
    .B(\system_expander.irq_fall_ctrl.io_masks[0] ),
    .X(_0408_));
 sg13g2_and2_1 _0979_ (.A(net304),
    .B(net302),
    .X(_0409_));
 sg13g2_nor2_1 _0981_ (.A(net304),
    .B(net302),
    .Y(_0411_));
 sg13g2_a221oi_1 _0982_ (.B2(_0409_),
    .C1(_0411_),
    .B1(_0408_),
    .A1(_0141_),
    .Y(_0412_),
    .A2(sg13g2_IOPad_io_gpio_0_c2p_en));
 sg13g2_nor3_1 _0983_ (.A(net306),
    .B(net301),
    .C(_0412_),
    .Y(_0413_));
 sg13g2_a22oi_1 _0984_ (.Y(_0414_),
    .B1(_0177_),
    .B2(\system_expander.irq_fall_ctrl.io_masks[0] ),
    .A2(_0134_),
    .A1(\system_expander.irq_rise_ctrl.io_masks[0] ));
 sg13g2_nor2b_1 _0985_ (.A(_0414_),
    .B_N(_0249_),
    .Y(_0415_));
 sg13g2_nor4_1 _0986_ (.A(net276),
    .B(_0407_),
    .C(_0413_),
    .D(_0415_),
    .Y(_0416_));
 sg13g2_a21o_1 _0987_ (.A2(net292),
    .A1(\system_expander.irq_low_ctrl.pendings[0] ),
    .B1(_0249_),
    .X(_0417_));
 sg13g2_nand3_1 _0988_ (.B(_0316_),
    .C(_0417_),
    .A(\system_expander.irq_low_ctrl.io_masks[0] ),
    .Y(_0418_));
 sg13g2_nand3_1 _0989_ (.B(\system_expander.irq_high_ctrl.io_masks[0] ),
    .C(_0270_),
    .A(\system_expander.irq_high_ctrl.pendings[0] ),
    .Y(_0419_));
 sg13g2_and2_1 _0990_ (.A(_0418_),
    .B(_0419_),
    .X(_0420_));
 sg13g2_nand3_1 _0991_ (.B(_0141_),
    .C(_0316_),
    .A(_0145_),
    .Y(_0421_));
 sg13g2_or2_1 _0992_ (.X(_0422_),
    .B(_0421_),
    .A(_0398_));
 sg13g2_o21ai_1 _0994_ (.B1(net329),
    .Y(_0424_),
    .A1(\system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[0] ),
    .A2(_0422_));
 sg13g2_a221oi_1 _0995_ (.B2(_0420_),
    .C1(_0424_),
    .B1(_0416_),
    .A1(_0397_),
    .Y(_0088_),
    .A2(net276));
 sg13g2_inv_1 _0996_ (.Y(_0425_),
    .A(\system_expander.link_data[1] ));
 sg13g2_nand2_1 _0997_ (.Y(_0426_),
    .A(\system_expander.irq_fall_ctrl.pendings[1] ),
    .B(\system_expander.irq_fall_ctrl.io_masks[1] ));
 sg13g2_nand2_1 _0998_ (.Y(_0427_),
    .A(sg13g2_IOPad_io_gpio_1_c2p_en),
    .B(_0176_));
 sg13g2_o21ai_1 _0999_ (.B1(_0427_),
    .Y(_0428_),
    .A1(_0351_),
    .A2(_0426_));
 sg13g2_a22oi_1 _1000_ (.Y(_0429_),
    .B1(_0409_),
    .B2(\system_expander.irq_high_ctrl.io_masks[1] ),
    .A2(_0411_),
    .A1(sg13g2_IOPad_io_gpio_1_c2p));
 sg13g2_nor2b_1 _1001_ (.A(net304),
    .B_N(net301),
    .Y(_0430_));
 sg13g2_and2_1 _1003_ (.A(\system_expander.irq_high_ctrl.pendings[1] ),
    .B(\system_expander.irq_high_ctrl.io_masks[1] ),
    .X(_0432_));
 sg13g2_nor2b_1 _1004_ (.A(net301),
    .B_N(net304),
    .Y(_0433_));
 sg13g2_a22oi_1 _1005_ (.Y(_0434_),
    .B1(_0432_),
    .B2(_0433_),
    .A2(_0430_),
    .A1(\system_expander.irq_rise_ctrl.io_masks[1] ));
 sg13g2_or2_1 _1006_ (.X(_0435_),
    .B(_0434_),
    .A(net302));
 sg13g2_o21ai_1 _1007_ (.B1(_0435_),
    .Y(_0436_),
    .A1(net301),
    .A2(_0429_));
 sg13g2_nor2_1 _1008_ (.A(_0122_),
    .B(_0174_),
    .Y(_0437_));
 sg13g2_a22oi_1 _1009_ (.Y(_0438_),
    .B1(_0436_),
    .B2(_0437_),
    .A2(_0428_),
    .A1(net293));
 sg13g2_and2_1 _1010_ (.A(\system_expander.irq_low_ctrl.pendings[1] ),
    .B(\system_expander.irq_low_ctrl.io_masks[1] ),
    .X(_0439_));
 sg13g2_nand3b_1 _1011_ (.B(net292),
    .C(_0439_),
    .Y(_0440_),
    .A_N(net305));
 sg13g2_nand3_1 _1012_ (.B(\system_expander.irq_fall_ctrl.io_masks[1] ),
    .C(_0249_),
    .A(net305),
    .Y(_0441_));
 sg13g2_a21oi_2 _1013_ (.B1(net306),
    .Y(_0442_),
    .A2(_0441_),
    .A1(_0440_));
 sg13g2_and2_1 _1014_ (.A(\system_expander.irq_rise_ctrl.pendings[1] ),
    .B(\system_expander.irq_rise_ctrl.io_masks[1] ),
    .X(_0443_));
 sg13g2_nand4_1 _1015_ (.B(_0327_),
    .C(_0399_),
    .A(\system_expander.link_state[2] ),
    .Y(_0444_),
    .D(_0421_));
 sg13g2_a221oi_1 _1017_ (.B2(_0443_),
    .C1(_0444_),
    .B1(net279),
    .A1(\system_expander.irq_low_ctrl.io_masks[1] ),
    .Y(_0446_),
    .A2(net280));
 sg13g2_nor2b_1 _1018_ (.A(_0442_),
    .B_N(_0446_),
    .Y(_0447_));
 sg13g2_o21ai_1 _1019_ (.B1(net329),
    .Y(_0448_),
    .A1(\system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[1] ),
    .A2(_0422_));
 sg13g2_a221oi_1 _1020_ (.B2(_0447_),
    .C1(_0448_),
    .B1(_0438_),
    .A1(_0425_),
    .Y(_0089_),
    .A2(net276));
 sg13g2_inv_1 _1021_ (.Y(_0449_),
    .A(\system_expander.link_data[2] ));
 sg13g2_nand2_1 _1022_ (.Y(_0450_),
    .A(\system_expander.irq_rise_ctrl.pendings[2] ),
    .B(\system_expander.irq_rise_ctrl.io_masks[2] ));
 sg13g2_nand3_1 _1023_ (.B(\system_expander.irq_fall_ctrl.io_masks[2] ),
    .C(net293),
    .A(\system_expander.irq_fall_ctrl.pendings[2] ),
    .Y(_0451_));
 sg13g2_o21ai_1 _1024_ (.B1(_0451_),
    .Y(_0452_),
    .A1(_0350_),
    .A2(_0450_));
 sg13g2_a21oi_1 _1025_ (.A1(net292),
    .A2(_0452_),
    .Y(_0453_),
    .B1(_0444_));
 sg13g2_nand2_1 _1026_ (.Y(_0454_),
    .A(\system_expander.irq_rise_ctrl.io_masks[2] ),
    .B(_0430_));
 sg13g2_nand3_1 _1027_ (.B(\system_expander.irq_high_ctrl.io_masks[2] ),
    .C(_0433_),
    .A(\system_expander.irq_high_ctrl.pendings[2] ),
    .Y(_0455_));
 sg13g2_a21oi_1 _1028_ (.A1(_0454_),
    .A2(_0455_),
    .Y(_0456_),
    .B1(net291));
 sg13g2_nand2_1 _1029_ (.Y(_0457_),
    .A(_0145_),
    .B(_0327_));
 sg13g2_a22oi_1 _1030_ (.Y(_0458_),
    .B1(_0409_),
    .B2(\system_expander.irq_high_ctrl.io_masks[2] ),
    .A2(_0411_),
    .A1(sg13g2_IOPad_io_gpio_2_c2p));
 sg13g2_o21ai_1 _1031_ (.B1(net306),
    .Y(_0459_),
    .A1(_0457_),
    .A2(_0458_));
 sg13g2_nor2_2 _1032_ (.A(net305),
    .B(_0351_),
    .Y(_0460_));
 sg13g2_and2_1 _1033_ (.A(\system_expander.irq_low_ctrl.pendings[2] ),
    .B(\system_expander.irq_low_ctrl.io_masks[2] ),
    .X(_0461_));
 sg13g2_mux2_1 _1034_ (.A0(sg13g2_IOPad_io_gpio_2_c2p_en),
    .A1(\system_expander.irq_fall_ctrl.io_masks[2] ),
    .S(net301),
    .X(_0462_));
 sg13g2_a22oi_1 _1035_ (.Y(_0463_),
    .B1(_0462_),
    .B2(net304),
    .A2(_0430_),
    .A1(\system_expander.irq_low_ctrl.io_masks[2] ));
 sg13g2_o21ai_1 _1036_ (.B1(_0122_),
    .Y(_0464_),
    .A1(net291),
    .A2(_0463_));
 sg13g2_a21o_1 _1037_ (.A2(_0461_),
    .A1(_0460_),
    .B1(_0464_),
    .X(_0465_));
 sg13g2_o21ai_1 _1038_ (.B1(_0465_),
    .Y(_0466_),
    .A1(_0456_),
    .A2(_0459_));
 sg13g2_o21ai_1 _1039_ (.B1(net329),
    .Y(_0467_),
    .A1(\system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[2] ),
    .A2(_0422_));
 sg13g2_a221oi_1 _1040_ (.B2(_0466_),
    .C1(_0467_),
    .B1(_0453_),
    .A1(_0449_),
    .Y(_0090_),
    .A2(_0400_));
 sg13g2_inv_1 _1041_ (.Y(_0468_),
    .A(\system_expander.link_data[3] ));
 sg13g2_nand3_1 _1042_ (.B(\system_expander.irq_low_ctrl.io_masks[3] ),
    .C(net292),
    .A(\system_expander.irq_low_ctrl.pendings[3] ),
    .Y(_0469_));
 sg13g2_nand3_1 _1043_ (.B(\system_expander.irq_fall_ctrl.io_masks[3] ),
    .C(_0249_),
    .A(net304),
    .Y(_0470_));
 sg13g2_o21ai_1 _1044_ (.B1(_0470_),
    .Y(_0471_),
    .A1(net304),
    .A2(_0469_));
 sg13g2_nand2_1 _1045_ (.Y(_0472_),
    .A(_0122_),
    .B(_0471_));
 sg13g2_and2_1 _1046_ (.A(\system_expander.irq_fall_ctrl.pendings[3] ),
    .B(\system_expander.irq_fall_ctrl.io_masks[3] ),
    .X(_0473_));
 sg13g2_a22oi_1 _1047_ (.Y(_0474_),
    .B1(net292),
    .B2(_0473_),
    .A2(_0176_),
    .A1(sg13g2_IOPad_io_gpio_3_c2p_en));
 sg13g2_nand2b_1 _1048_ (.Y(_0475_),
    .B(net293),
    .A_N(_0474_));
 sg13g2_a22oi_1 _1049_ (.Y(_0476_),
    .B1(_0409_),
    .B2(\system_expander.irq_high_ctrl.io_masks[3] ),
    .A2(_0411_),
    .A1(sg13g2_IOPad_io_gpio_3_c2p));
 sg13g2_nor2_1 _1050_ (.A(net301),
    .B(_0476_),
    .Y(_0477_));
 sg13g2_nand2_1 _1051_ (.Y(_0478_),
    .A(\system_expander.irq_rise_ctrl.io_masks[3] ),
    .B(_0430_));
 sg13g2_nand3_1 _1052_ (.B(\system_expander.irq_high_ctrl.io_masks[3] ),
    .C(_0433_),
    .A(\system_expander.irq_high_ctrl.pendings[3] ),
    .Y(_0479_));
 sg13g2_a21oi_1 _1053_ (.A1(_0478_),
    .A2(_0479_),
    .Y(_0480_),
    .B1(net302));
 sg13g2_o21ai_1 _1054_ (.B1(_0437_),
    .Y(_0481_),
    .A1(_0477_),
    .A2(_0480_));
 sg13g2_and2_1 _1055_ (.A(\system_expander.irq_rise_ctrl.pendings[3] ),
    .B(\system_expander.irq_rise_ctrl.io_masks[3] ),
    .X(_0482_));
 sg13g2_a221oi_1 _1056_ (.B2(_0482_),
    .C1(_0444_),
    .B1(_0353_),
    .A1(\system_expander.irq_low_ctrl.io_masks[3] ),
    .Y(_0483_),
    .A2(net280));
 sg13g2_and3_1 _1057_ (.X(_0484_),
    .A(_0475_),
    .B(_0481_),
    .C(_0483_));
 sg13g2_o21ai_1 _1058_ (.B1(net329),
    .Y(_0485_),
    .A1(\system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[3] ),
    .A2(_0422_));
 sg13g2_a221oi_1 _1059_ (.B2(_0484_),
    .C1(_0485_),
    .B1(_0472_),
    .A1(_0468_),
    .Y(_0091_),
    .A2(_0400_));
 sg13g2_inv_1 _1060_ (.Y(_0486_),
    .A(\system_expander.link_data[4] ));
 sg13g2_and2_1 _1061_ (.A(\system_expander.irq_fall_ctrl.pendings[4] ),
    .B(\system_expander.irq_fall_ctrl.io_masks[4] ),
    .X(_0487_));
 sg13g2_and2_1 _1062_ (.A(\system_expander.irq_rise_ctrl.pendings[4] ),
    .B(\system_expander.irq_rise_ctrl.io_masks[4] ),
    .X(_0488_));
 sg13g2_a22oi_1 _1063_ (.Y(_0489_),
    .B1(_0488_),
    .B2(_0134_),
    .A2(_0487_),
    .A1(net293));
 sg13g2_nor2_1 _1064_ (.A(_0351_),
    .B(_0489_),
    .Y(_0490_));
 sg13g2_nor2_1 _1065_ (.A(_0444_),
    .B(_0490_),
    .Y(_0491_));
 sg13g2_nand2_1 _1066_ (.Y(_0492_),
    .A(\system_expander.irq_rise_ctrl.io_masks[4] ),
    .B(_0430_));
 sg13g2_nand3_1 _1067_ (.B(\system_expander.irq_high_ctrl.io_masks[4] ),
    .C(_0433_),
    .A(\system_expander.irq_high_ctrl.pendings[4] ),
    .Y(_0493_));
 sg13g2_a21oi_1 _1068_ (.A1(_0492_),
    .A2(_0493_),
    .Y(_0494_),
    .B1(net291));
 sg13g2_a22oi_1 _1069_ (.Y(_0495_),
    .B1(_0409_),
    .B2(\system_expander.irq_high_ctrl.io_masks[4] ),
    .A2(_0411_),
    .A1(sg13g2_IOPad_io_gpio_4_c2p));
 sg13g2_o21ai_1 _1070_ (.B1(net306),
    .Y(_0496_),
    .A1(_0457_),
    .A2(_0495_));
 sg13g2_and2_1 _1071_ (.A(\system_expander.irq_low_ctrl.pendings[4] ),
    .B(\system_expander.irq_low_ctrl.io_masks[4] ),
    .X(_0497_));
 sg13g2_mux2_1 _1072_ (.A0(sg13g2_IOPad_io_gpio_4_c2p_en),
    .A1(\system_expander.irq_fall_ctrl.io_masks[4] ),
    .S(net301),
    .X(_0498_));
 sg13g2_a22oi_1 _1073_ (.Y(_0499_),
    .B1(_0498_),
    .B2(net304),
    .A2(_0430_),
    .A1(\system_expander.irq_low_ctrl.io_masks[4] ));
 sg13g2_o21ai_1 _1074_ (.B1(_0122_),
    .Y(_0500_),
    .A1(net291),
    .A2(_0499_));
 sg13g2_a21o_1 _1075_ (.A2(_0497_),
    .A1(_0460_),
    .B1(_0500_),
    .X(_0501_));
 sg13g2_o21ai_1 _1076_ (.B1(_0501_),
    .Y(_0502_),
    .A1(_0494_),
    .A2(_0496_));
 sg13g2_o21ai_1 _1077_ (.B1(net329),
    .Y(_0503_),
    .A1(\system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[4] ),
    .A2(_0422_));
 sg13g2_a221oi_1 _1078_ (.B2(_0502_),
    .C1(_0503_),
    .B1(_0491_),
    .A1(_0486_),
    .Y(_0092_),
    .A2(_0400_));
 sg13g2_inv_1 _1079_ (.Y(_0504_),
    .A(\system_expander.link_data[5] ));
 sg13g2_mux2_1 _1080_ (.A0(sg13g2_IOPad_io_gpio_5_c2p),
    .A1(\system_expander.irq_rise_ctrl.io_masks[5] ),
    .S(net300),
    .X(_0505_));
 sg13g2_mux2_1 _1081_ (.A0(sg13g2_IOPad_io_gpio_5_c2p_en),
    .A1(\system_expander.irq_fall_ctrl.io_masks[5] ),
    .S(net300),
    .X(_0506_));
 sg13g2_a22oi_1 _1082_ (.Y(_0507_),
    .B1(_0506_),
    .B2(net293),
    .A2(_0505_),
    .A1(_0134_));
 sg13g2_nand3_1 _1083_ (.B(\system_expander.irq_low_ctrl.io_masks[5] ),
    .C(_0316_),
    .A(net300),
    .Y(_0508_));
 sg13g2_a21oi_1 _1084_ (.A1(_0507_),
    .A2(_0508_),
    .Y(_0509_),
    .B1(net291));
 sg13g2_nand2_1 _1085_ (.Y(_0510_),
    .A(_0433_),
    .B(_0437_));
 sg13g2_o21ai_1 _1086_ (.B1(\system_expander.irq_high_ctrl.io_masks[5] ),
    .Y(_0511_),
    .A1(\system_expander.link_regAddr[2] ),
    .A2(\system_expander.irq_high_ctrl.pendings[5] ));
 sg13g2_nor2_1 _1087_ (.A(_0510_),
    .B(_0511_),
    .Y(_0512_));
 sg13g2_nor3_1 _1088_ (.A(_0444_),
    .B(_0509_),
    .C(_0512_),
    .Y(_0513_));
 sg13g2_and2_1 _1089_ (.A(\system_expander.irq_fall_ctrl.pendings[5] ),
    .B(\system_expander.irq_fall_ctrl.io_masks[5] ),
    .X(_0514_));
 sg13g2_nand2_1 _1090_ (.Y(_0515_),
    .A(\system_expander.irq_low_ctrl.pendings[5] ),
    .B(\system_expander.irq_low_ctrl.io_masks[5] ));
 sg13g2_nand3_1 _1091_ (.B(\system_expander.irq_rise_ctrl.pendings[5] ),
    .C(\system_expander.irq_rise_ctrl.io_masks[5] ),
    .A(net307),
    .Y(_0516_));
 sg13g2_o21ai_1 _1092_ (.B1(_0516_),
    .Y(_0517_),
    .A1(net307),
    .A2(_0515_));
 sg13g2_a22oi_1 _1093_ (.Y(_0518_),
    .B1(_0517_),
    .B2(_0460_),
    .A2(_0514_),
    .A1(net286));
 sg13g2_o21ai_1 _1094_ (.B1(net329),
    .Y(_0519_),
    .A1(\system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[5] ),
    .A2(_0422_));
 sg13g2_a221oi_1 _1095_ (.B2(_0518_),
    .C1(_0519_),
    .B1(_0513_),
    .A1(_0504_),
    .Y(_0093_),
    .A2(net276));
 sg13g2_inv_1 _1096_ (.Y(_0520_),
    .A(\system_expander.link_data[6] ));
 sg13g2_mux2_1 _1097_ (.A0(sg13g2_IOPad_io_gpio_6_c2p),
    .A1(\system_expander.irq_rise_ctrl.io_masks[6] ),
    .S(net300),
    .X(_0521_));
 sg13g2_mux2_1 _1098_ (.A0(sg13g2_IOPad_io_gpio_6_c2p_en),
    .A1(\system_expander.irq_fall_ctrl.io_masks[6] ),
    .S(net300),
    .X(_0522_));
 sg13g2_a22oi_1 _1099_ (.Y(_0523_),
    .B1(_0522_),
    .B2(net293),
    .A2(_0521_),
    .A1(_0134_));
 sg13g2_nand3_1 _1100_ (.B(\system_expander.irq_low_ctrl.io_masks[6] ),
    .C(_0316_),
    .A(net300),
    .Y(_0524_));
 sg13g2_a21oi_1 _1101_ (.A1(_0523_),
    .A2(_0524_),
    .Y(_0525_),
    .B1(net291));
 sg13g2_o21ai_1 _1102_ (.B1(\system_expander.irq_high_ctrl.io_masks[6] ),
    .Y(_0526_),
    .A1(\system_expander.link_regAddr[2] ),
    .A2(\system_expander.irq_high_ctrl.pendings[6] ));
 sg13g2_nor2_1 _1103_ (.A(_0510_),
    .B(_0526_),
    .Y(_0527_));
 sg13g2_nor3_1 _1104_ (.A(_0444_),
    .B(_0525_),
    .C(_0527_),
    .Y(_0528_));
 sg13g2_and2_1 _1105_ (.A(\system_expander.irq_fall_ctrl.pendings[6] ),
    .B(\system_expander.irq_fall_ctrl.io_masks[6] ),
    .X(_0529_));
 sg13g2_nand2_1 _1106_ (.Y(_0530_),
    .A(\system_expander.irq_low_ctrl.pendings[6] ),
    .B(\system_expander.irq_low_ctrl.io_masks[6] ));
 sg13g2_nand3_1 _1107_ (.B(\system_expander.irq_rise_ctrl.pendings[6] ),
    .C(\system_expander.irq_rise_ctrl.io_masks[6] ),
    .A(net307),
    .Y(_0531_));
 sg13g2_o21ai_1 _1108_ (.B1(_0531_),
    .Y(_0532_),
    .A1(net307),
    .A2(_0530_));
 sg13g2_a22oi_1 _1109_ (.Y(_0533_),
    .B1(_0532_),
    .B2(_0460_),
    .A2(_0529_),
    .A1(net286));
 sg13g2_o21ai_1 _1110_ (.B1(net329),
    .Y(_0534_),
    .A1(\system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[6] ),
    .A2(_0422_));
 sg13g2_a221oi_1 _1111_ (.B2(_0533_),
    .C1(_0534_),
    .B1(_0528_),
    .A1(_0520_),
    .Y(_0094_),
    .A2(net276));
 sg13g2_inv_1 _1112_ (.Y(_0535_),
    .A(\system_expander.link_data[7] ));
 sg13g2_nand3_1 _1113_ (.B(\system_expander.irq_fall_ctrl.io_masks[7] ),
    .C(net293),
    .A(\system_expander.irq_fall_ctrl.pendings[7] ),
    .Y(_0536_));
 sg13g2_nand3_1 _1114_ (.B(\system_expander.irq_rise_ctrl.io_masks[7] ),
    .C(_0134_),
    .A(\system_expander.irq_rise_ctrl.pendings[7] ),
    .Y(_0537_));
 sg13g2_a21oi_1 _1115_ (.A1(_0536_),
    .A2(_0537_),
    .Y(_0538_),
    .B1(_0351_));
 sg13g2_nor2_1 _1116_ (.A(_0444_),
    .B(_0538_),
    .Y(_0539_));
 sg13g2_nand2_1 _1117_ (.Y(_0540_),
    .A(\system_expander.irq_rise_ctrl.io_masks[7] ),
    .B(_0430_));
 sg13g2_nand3_1 _1118_ (.B(\system_expander.irq_high_ctrl.io_masks[7] ),
    .C(_0433_),
    .A(\system_expander.irq_high_ctrl.pendings[7] ),
    .Y(_0541_));
 sg13g2_a21oi_1 _1119_ (.A1(_0540_),
    .A2(_0541_),
    .Y(_0542_),
    .B1(net291));
 sg13g2_a22oi_1 _1120_ (.Y(_0543_),
    .B1(_0409_),
    .B2(\system_expander.irq_high_ctrl.io_masks[7] ),
    .A2(_0411_),
    .A1(sg13g2_IOPad_io_gpio_7_c2p));
 sg13g2_o21ai_1 _1121_ (.B1(net306),
    .Y(_0544_),
    .A1(_0457_),
    .A2(_0543_));
 sg13g2_and2_1 _1122_ (.A(\system_expander.irq_low_ctrl.pendings[7] ),
    .B(\system_expander.irq_low_ctrl.io_masks[7] ),
    .X(_0545_));
 sg13g2_mux2_1 _1123_ (.A0(sg13g2_IOPad_io_gpio_7_c2p_en),
    .A1(\system_expander.irq_fall_ctrl.io_masks[7] ),
    .S(net300),
    .X(_0546_));
 sg13g2_a22oi_1 _1124_ (.Y(_0547_),
    .B1(_0546_),
    .B2(net303),
    .A2(_0430_),
    .A1(\system_expander.irq_low_ctrl.io_masks[7] ));
 sg13g2_o21ai_1 _1125_ (.B1(_0122_),
    .Y(_0548_),
    .A1(net291),
    .A2(_0547_));
 sg13g2_a21o_1 _1126_ (.A2(_0545_),
    .A1(_0460_),
    .B1(_0548_),
    .X(_0549_));
 sg13g2_o21ai_1 _1127_ (.B1(_0549_),
    .Y(_0550_),
    .A1(_0542_),
    .A2(_0544_));
 sg13g2_o21ai_1 _1128_ (.B1(net329),
    .Y(_0551_),
    .A1(\system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[7] ),
    .A2(_0422_));
 sg13g2_a221oi_1 _1129_ (.B2(_0550_),
    .C1(_0551_),
    .B1(_0539_),
    .A1(_0535_),
    .Y(_0095_),
    .A2(net276));
 sg13g2_nand2_1 _1130_ (.Y(_0552_),
    .A(\system_expander.i2cCtrl_io_cmd_valid ),
    .B(_0119_));
 sg13g2_o21ai_1 _1131_ (.B1(_0552_),
    .Y(_0553_),
    .A1(\system_expander.i2cCtrl_io_cmd_valid ),
    .A2(\system_expander.link_error ));
 sg13g2_nand2_1 _1132_ (.Y(_0554_),
    .A(_0327_),
    .B(_0399_));
 sg13g2_a21oi_1 _1133_ (.A1(net298),
    .A2(_0421_),
    .Y(_0555_),
    .B1(\system_expander.link_state[2] ));
 sg13g2_o21ai_1 _1134_ (.B1(_0110_),
    .Y(_0556_),
    .A1(_0554_),
    .A2(_0555_));
 sg13g2_inv_1 _1135_ (.Y(_0557_),
    .A(\system_expander.link_error ));
 sg13g2_a221oi_1 _1136_ (.B2(_0557_),
    .C1(_0114_),
    .B1(_0556_),
    .A1(\system_expander.link_state[0] ),
    .Y(_0096_),
    .A2(_0553_));
 sg13g2_a21oi_1 _1137_ (.A1(\system_expander.irq_rise_ctrl.pendings[6] ),
    .A2(\system_expander.irq_rise_ctrl.io_masks[6] ),
    .Y(_0558_),
    .B1(_0488_));
 sg13g2_a21oi_1 _1138_ (.A1(\system_expander.irq_low_ctrl.pendings[5] ),
    .A2(\system_expander.irq_low_ctrl.io_masks[5] ),
    .Y(_0559_),
    .B1(_0529_));
 sg13g2_a21oi_1 _1139_ (.A1(\system_expander.irq_rise_ctrl.pendings[5] ),
    .A2(\system_expander.irq_rise_ctrl.io_masks[5] ),
    .Y(_0560_),
    .B1(_0514_));
 sg13g2_a21oi_1 _1140_ (.A1(\system_expander.irq_high_ctrl.pendings[4] ),
    .A2(\system_expander.irq_high_ctrl.io_masks[4] ),
    .Y(_0561_),
    .B1(_0497_));
 sg13g2_nand4_1 _1141_ (.B(_0559_),
    .C(_0560_),
    .A(_0558_),
    .Y(_0562_),
    .D(_0561_));
 sg13g2_a22oi_1 _1142_ (.Y(_0563_),
    .B1(\system_expander.irq_low_ctrl.io_masks[6] ),
    .B2(\system_expander.irq_low_ctrl.pendings[6] ),
    .A2(\system_expander.irq_high_ctrl.io_masks[5] ),
    .A1(\system_expander.irq_high_ctrl.pendings[5] ));
 sg13g2_a22oi_1 _1143_ (.Y(_0564_),
    .B1(\system_expander.irq_high_ctrl.io_masks[6] ),
    .B2(\system_expander.irq_high_ctrl.pendings[6] ),
    .A2(\system_expander.irq_low_ctrl.io_masks[0] ),
    .A1(\system_expander.irq_low_ctrl.pendings[0] ));
 sg13g2_a22oi_1 _1144_ (.Y(_0565_),
    .B1(\system_expander.irq_fall_ctrl.io_masks[7] ),
    .B2(\system_expander.irq_fall_ctrl.pendings[7] ),
    .A2(\system_expander.irq_rise_ctrl.io_masks[7] ),
    .A1(\system_expander.irq_rise_ctrl.pendings[7] ));
 sg13g2_a21oi_1 _1145_ (.A1(\system_expander.irq_high_ctrl.pendings[7] ),
    .A2(\system_expander.irq_high_ctrl.io_masks[7] ),
    .Y(_0566_),
    .B1(_0545_));
 sg13g2_nand4_1 _1146_ (.B(_0564_),
    .C(_0565_),
    .A(_0563_),
    .Y(_0567_),
    .D(_0566_));
 sg13g2_nor4_1 _1147_ (.A(_0432_),
    .B(_0443_),
    .C(_0439_),
    .D(_0487_),
    .Y(_0568_));
 sg13g2_a22oi_1 _1148_ (.Y(_0569_),
    .B1(\system_expander.irq_fall_ctrl.io_masks[0] ),
    .B2(\system_expander.irq_fall_ctrl.pendings[0] ),
    .A2(\system_expander.irq_high_ctrl.io_masks[0] ),
    .A1(\system_expander.irq_high_ctrl.pendings[0] ));
 sg13g2_nand4_1 _1149_ (.B(_0426_),
    .C(_0568_),
    .A(_0402_),
    .Y(_0570_),
    .D(_0569_));
 sg13g2_a22oi_1 _1150_ (.Y(_0571_),
    .B1(\system_expander.irq_high_ctrl.io_masks[3] ),
    .B2(\system_expander.irq_high_ctrl.pendings[3] ),
    .A2(\system_expander.irq_fall_ctrl.io_masks[2] ),
    .A1(\system_expander.irq_fall_ctrl.pendings[2] ));
 sg13g2_a21oi_1 _1151_ (.A1(\system_expander.irq_low_ctrl.pendings[3] ),
    .A2(\system_expander.irq_low_ctrl.io_masks[3] ),
    .Y(_0572_),
    .B1(_0482_));
 sg13g2_nor2_1 _1152_ (.A(_0461_),
    .B(_0473_),
    .Y(_0573_));
 sg13g2_a22oi_1 _1153_ (.Y(_0574_),
    .B1(\system_expander.irq_rise_ctrl.io_masks[2] ),
    .B2(\system_expander.irq_rise_ctrl.pendings[2] ),
    .A2(\system_expander.irq_high_ctrl.io_masks[2] ),
    .A1(\system_expander.irq_high_ctrl.pendings[2] ));
 sg13g2_nand4_1 _1154_ (.B(_0572_),
    .C(_0573_),
    .A(_0571_),
    .Y(_0575_),
    .D(_0574_));
 sg13g2_or4_1 _1155_ (.A(_0562_),
    .B(_0567_),
    .C(_0570_),
    .D(_0575_),
    .X(\system_expander.i2cCtrl_io_interrupts[0] ));
 sg13g2_nor2_1 _1156_ (.A(\system_expander.link_state[0] ),
    .B(\system_expander.i2cCtrl_io_cmd_ready ),
    .Y(\system_expander.i2cCtrl_io_rsp_valid ));
 sg13g2_buf_16 clkbuf_0_clock (.X(clknet_0_clock),
    .A(clock));
 sg13g2_buf_16 clkbuf_0_clock_regs (.X(clknet_0_clock_regs),
    .A(clock_regs));
 sg13g2_buf_16 clkbuf_1_0__f_clock (.X(clknet_1_0__leaf_clock),
    .A(clknet_0_clock));
 sg13g2_buf_16 clkbuf_4_0_0_clock_regs (.X(clknet_4_0_0_clock_regs),
    .A(clknet_0_clock_regs));
 sg13g2_buf_16 clkbuf_4_10_0_clock_regs (.X(clknet_4_10_0_clock_regs),
    .A(clknet_0_clock_regs));
 sg13g2_buf_16 clkbuf_4_11_0_clock_regs (.X(clknet_4_11_0_clock_regs),
    .A(clknet_0_clock_regs));
 sg13g2_buf_16 clkbuf_4_12_0_clock_regs (.X(clknet_4_12_0_clock_regs),
    .A(clknet_0_clock_regs));
 sg13g2_buf_16 clkbuf_4_13_0_clock_regs (.X(clknet_4_13_0_clock_regs),
    .A(clknet_0_clock_regs));
 sg13g2_buf_16 clkbuf_4_14_0_clock_regs (.X(clknet_4_14_0_clock_regs),
    .A(clknet_0_clock_regs));
 sg13g2_buf_16 clkbuf_4_15_0_clock_regs (.X(clknet_4_15_0_clock_regs),
    .A(clknet_0_clock_regs));
 sg13g2_buf_16 clkbuf_4_1_0_clock_regs (.X(clknet_4_1_0_clock_regs),
    .A(clknet_0_clock_regs));
 sg13g2_buf_16 clkbuf_4_2_0_clock_regs (.X(clknet_4_2_0_clock_regs),
    .A(clknet_0_clock_regs));
 sg13g2_buf_16 clkbuf_4_3_0_clock_regs (.X(clknet_4_3_0_clock_regs),
    .A(clknet_0_clock_regs));
 sg13g2_buf_16 clkbuf_4_4_0_clock_regs (.X(clknet_4_4_0_clock_regs),
    .A(clknet_0_clock_regs));
 sg13g2_buf_16 clkbuf_4_5_0_clock_regs (.X(clknet_4_5_0_clock_regs),
    .A(clknet_0_clock_regs));
 sg13g2_buf_16 clkbuf_4_6_0_clock_regs (.X(clknet_4_6_0_clock_regs),
    .A(clknet_0_clock_regs));
 sg13g2_buf_16 clkbuf_4_7_0_clock_regs (.X(clknet_4_7_0_clock_regs),
    .A(clknet_0_clock_regs));
 sg13g2_buf_16 clkbuf_4_8_0_clock_regs (.X(clknet_4_8_0_clock_regs),
    .A(clknet_0_clock_regs));
 sg13g2_buf_16 clkbuf_4_9_0_clock_regs (.X(clknet_4_9_0_clock_regs),
    .A(clknet_0_clock_regs));
 sg13g2_buf_16 clkbuf_5_0__f_clock_regs (.X(clknet_5_0__leaf_clock_regs),
    .A(clknet_4_0_0_clock_regs));
 sg13g2_buf_16 clkbuf_5_10__f_clock_regs (.X(clknet_5_10__leaf_clock_regs),
    .A(clknet_4_5_0_clock_regs));
 sg13g2_buf_16 clkbuf_5_11__f_clock_regs (.X(clknet_5_11__leaf_clock_regs),
    .A(clknet_4_5_0_clock_regs));
 sg13g2_buf_16 clkbuf_5_12__f_clock_regs (.X(clknet_5_12__leaf_clock_regs),
    .A(clknet_4_6_0_clock_regs));
 sg13g2_buf_16 clkbuf_5_13__f_clock_regs (.X(clknet_5_13__leaf_clock_regs),
    .A(clknet_4_6_0_clock_regs));
 sg13g2_buf_16 clkbuf_5_14__f_clock_regs (.X(clknet_5_14__leaf_clock_regs),
    .A(clknet_4_7_0_clock_regs));
 sg13g2_buf_16 clkbuf_5_15__f_clock_regs (.X(clknet_5_15__leaf_clock_regs),
    .A(clknet_4_7_0_clock_regs));
 sg13g2_buf_16 clkbuf_5_16__f_clock_regs (.X(clknet_5_16__leaf_clock_regs),
    .A(clknet_4_8_0_clock_regs));
 sg13g2_buf_16 clkbuf_5_17__f_clock_regs (.X(clknet_5_17__leaf_clock_regs),
    .A(clknet_4_8_0_clock_regs));
 sg13g2_buf_16 clkbuf_5_18__f_clock_regs (.X(clknet_5_18__leaf_clock_regs),
    .A(clknet_4_9_0_clock_regs));
 sg13g2_buf_16 clkbuf_5_19__f_clock_regs (.X(clknet_5_19__leaf_clock_regs),
    .A(clknet_4_9_0_clock_regs));
 sg13g2_buf_16 clkbuf_5_1__f_clock_regs (.X(clknet_5_1__leaf_clock_regs),
    .A(clknet_4_0_0_clock_regs));
 sg13g2_buf_16 clkbuf_5_20__f_clock_regs (.X(clknet_5_20__leaf_clock_regs),
    .A(clknet_4_10_0_clock_regs));
 sg13g2_buf_16 clkbuf_5_21__f_clock_regs (.X(clknet_5_21__leaf_clock_regs),
    .A(clknet_4_10_0_clock_regs));
 sg13g2_buf_16 clkbuf_5_22__f_clock_regs (.X(clknet_5_22__leaf_clock_regs),
    .A(clknet_4_11_0_clock_regs));
 sg13g2_buf_16 clkbuf_5_23__f_clock_regs (.X(clknet_5_23__leaf_clock_regs),
    .A(clknet_4_11_0_clock_regs));
 sg13g2_buf_16 clkbuf_5_24__f_clock_regs (.X(clknet_5_24__leaf_clock_regs),
    .A(clknet_4_12_0_clock_regs));
 sg13g2_buf_16 clkbuf_5_25__f_clock_regs (.X(clknet_5_25__leaf_clock_regs),
    .A(clknet_4_12_0_clock_regs));
 sg13g2_buf_16 clkbuf_5_26__f_clock_regs (.X(clknet_5_26__leaf_clock_regs),
    .A(clknet_4_13_0_clock_regs));
 sg13g2_buf_16 clkbuf_5_27__f_clock_regs (.X(clknet_5_27__leaf_clock_regs),
    .A(clknet_4_13_0_clock_regs));
 sg13g2_buf_16 clkbuf_5_28__f_clock_regs (.X(clknet_5_28__leaf_clock_regs),
    .A(clknet_4_14_0_clock_regs));
 sg13g2_buf_16 clkbuf_5_29__f_clock_regs (.X(clknet_5_29__leaf_clock_regs),
    .A(clknet_4_14_0_clock_regs));
 sg13g2_buf_16 clkbuf_5_2__f_clock_regs (.X(clknet_5_2__leaf_clock_regs),
    .A(clknet_4_1_0_clock_regs));
 sg13g2_buf_16 clkbuf_5_30__f_clock_regs (.X(clknet_5_30__leaf_clock_regs),
    .A(clknet_4_15_0_clock_regs));
 sg13g2_buf_16 clkbuf_5_31__f_clock_regs (.X(clknet_5_31__leaf_clock_regs),
    .A(clknet_4_15_0_clock_regs));
 sg13g2_buf_16 clkbuf_5_3__f_clock_regs (.X(clknet_5_3__leaf_clock_regs),
    .A(clknet_4_1_0_clock_regs));
 sg13g2_buf_16 clkbuf_5_4__f_clock_regs (.X(clknet_5_4__leaf_clock_regs),
    .A(clknet_4_2_0_clock_regs));
 sg13g2_buf_16 clkbuf_5_5__f_clock_regs (.X(clknet_5_5__leaf_clock_regs),
    .A(clknet_4_2_0_clock_regs));
 sg13g2_buf_16 clkbuf_5_6__f_clock_regs (.X(clknet_5_6__leaf_clock_regs),
    .A(clknet_4_3_0_clock_regs));
 sg13g2_buf_16 clkbuf_5_7__f_clock_regs (.X(clknet_5_7__leaf_clock_regs),
    .A(clknet_4_3_0_clock_regs));
 sg13g2_buf_16 clkbuf_5_8__f_clock_regs (.X(clknet_5_8__leaf_clock_regs),
    .A(clknet_4_4_0_clock_regs));
 sg13g2_buf_16 clkbuf_5_9__f_clock_regs (.X(clknet_5_9__leaf_clock_regs),
    .A(clknet_4_4_0_clock_regs));
 sg13g2_buf_16 clkbuf_regs_0_clk_core (.X(clock_regs),
    .A(delaynet_2_clk_core));
 sg13g2_inv_1 clkload0 (.A(clknet_5_7__leaf_clock_regs));
 sg13g2_inv_1 clkload1 (.A(clknet_5_11__leaf_clock_regs));
 sg13g2_inv_1 clkload2 (.A(clknet_5_15__leaf_clock_regs));
 sg13g2_inv_1 clkload3 (.A(clknet_5_23__leaf_clock_regs));
 sg13g2_inv_1 clkload4 (.A(clknet_5_27__leaf_clock_regs));
 sg13g2_inv_1 clkload5 (.A(clknet_5_31__leaf_clock_regs));
 sg13g2_buf_16 delaybuf_0_clk_core (.X(delaynet_0_clk_core),
    .A(clock));
 sg13g2_buf_16 delaybuf_1_clk_core (.X(delaynet_1_clk_core),
    .A(delaynet_0_clk_core));
 sg13g2_buf_16 delaybuf_2_clk_core (.X(delaynet_2_clk_core),
    .A(delaynet_1_clk_core));
 sg13g2_buf_1 place277 (.A(_0400_),
    .X(net276));
 sg13g2_buf_1 place278 (.A(_0378_),
    .X(net277));
 sg13g2_buf_1 place279 (.A(_0378_),
    .X(net278));
 sg13g2_buf_1 place280 (.A(_0353_),
    .X(net279));
 sg13g2_buf_1 place281 (.A(_0329_),
    .X(net280));
 sg13g2_buf_1 place282 (.A(_0296_),
    .X(net281));
 sg13g2_buf_1 place283 (.A(_0296_),
    .X(net282));
 sg13g2_buf_1 place284 (.A(_0270_),
    .X(net283));
 sg13g2_buf_1 place285 (.A(_0250_),
    .X(net284));
 sg13g2_buf_1 place286 (.A(_0250_),
    .X(net285));
 sg13g2_buf_1 place287 (.A(_0224_),
    .X(net286));
 sg13g2_buf_1 place288 (.A(_0198_),
    .X(net287));
 sg13g2_buf_1 place289 (.A(_0198_),
    .X(net288));
 sg13g2_buf_1 place290 (.A(_0178_),
    .X(net289));
 sg13g2_buf_1 place291 (.A(_0178_),
    .X(net290));
 sg13g2_buf_1 place292 (.A(_0328_),
    .X(net291));
 sg13g2_buf_1 place293 (.A(_0223_),
    .X(net292));
 sg13g2_buf_1 place294 (.A(_0177_),
    .X(net293));
 sg13g2_buf_1 place295 (.A(_0119_),
    .X(net294));
 sg13g2_buf_1 place296 (.A(net296),
    .X(net295));
 sg13g2_buf_1 place297 (.A(net298),
    .X(net296));
 sg13g2_buf_1 place298 (.A(net298),
    .X(net297));
 sg13g2_buf_1 place299 (.A(\system_expander.link_state[4] ),
    .X(net298));
 sg13g2_buf_1 place300 (.A(\system_expander.link_state[4] ),
    .X(net299));
 sg13g2_buf_1 place301 (.A(\system_expander.link_regAddr[3] ),
    .X(net300));
 sg13g2_buf_1 place302 (.A(\system_expander.link_regAddr[3] ),
    .X(net301));
 sg13g2_buf_1 place303 (.A(\system_expander.link_regAddr[2] ),
    .X(net302));
 sg13g2_buf_1 place304 (.A(net305),
    .X(net303));
 sg13g2_buf_1 place305 (.A(net305),
    .X(net304));
 sg13g2_buf_1 place306 (.A(\system_expander.link_regAddr[1] ),
    .X(net305));
 sg13g2_buf_1 place307 (.A(net307),
    .X(net306));
 sg13g2_buf_1 place308 (.A(\system_expander.link_regAddr[0] ),
    .X(net307));
 sg13g2_buf_1 place309 (.A(\system_expander.i2cCtrl_io_cmd_payload_data[7] ),
    .X(net308));
 sg13g2_buf_1 place310 (.A(\system_expander.i2cCtrl_io_cmd_payload_data[6] ),
    .X(net309));
 sg13g2_buf_1 place311 (.A(\system_expander.i2cCtrl_io_cmd_payload_data[5] ),
    .X(net310));
 sg13g2_buf_1 place312 (.A(\system_expander.i2cCtrl_io_cmd_payload_data[4] ),
    .X(net311));
 sg13g2_buf_1 place313 (.A(\system_expander.i2cCtrl_io_cmd_payload_data[3] ),
    .X(net312));
 sg13g2_buf_1 place314 (.A(\system_expander.i2cCtrl_io_cmd_payload_data[2] ),
    .X(net313));
 sg13g2_buf_1 place315 (.A(\system_expander.i2cCtrl_io_cmd_payload_data[1] ),
    .X(net314));
 sg13g2_buf_1 place316 (.A(\system_expander.i2cCtrl_io_cmd_payload_data[0] ),
    .X(net315));
 sg13g2_buf_1 place317 (.A(net321),
    .X(net316));
 sg13g2_buf_1 place318 (.A(net318),
    .X(net317));
 sg13g2_buf_1 place319 (.A(net320),
    .X(net318));
 sg13g2_buf_1 place320 (.A(net320),
    .X(net319));
 sg13g2_buf_1 place321 (.A(net321),
    .X(net320));
 sg13g2_buf_1 place322 (.A(net328),
    .X(net321));
 sg13g2_buf_1 place323 (.A(net328),
    .X(net322));
 sg13g2_buf_1 place324 (.A(net327),
    .X(net323));
 sg13g2_buf_1 place325 (.A(net325),
    .X(net324));
 sg13g2_buf_1 place326 (.A(net327),
    .X(net325));
 sg13g2_buf_1 place327 (.A(net327),
    .X(net326));
 sg13g2_buf_1 place328 (.A(net328),
    .X(net327));
 sg13g2_buf_1 place329 (.A(_0114_),
    .X(net328));
 sg13g2_buf_1 place330 (.A(reset),
    .X(net329));
 sg13g2_IOPadIOVdd sg13g2_IOPadIOVdd_west_4 ();
 sg13g2_IOPadIOVss sg13g2_IOPadIOVss_west_3 ();
 sg13g2_IOPadVdd sg13g2_IOPadVdd_east_0 ();
 sg13g2_IOPadVss sg13g2_IOPadVss_east_1 ();
 sg13g2_IOPadIn sg13g2_IOPad_io_address_0 (.p2c(sg13g2_IOPad_io_address_0_p2c),
    .pad(io_address_0_PAD));
 sg13g2_IOPadIn sg13g2_IOPad_io_address_1 (.p2c(sg13g2_IOPad_io_address_1_p2c),
    .pad(io_address_1_PAD));
 sg13g2_IOPadIn sg13g2_IOPad_io_address_2 (.p2c(sg13g2_IOPad_io_address_2_p2c),
    .pad(io_address_2_PAD));
 sg13g2_IOPadIn sg13g2_IOPad_io_clock (.p2c(clock),
    .pad(io_clock_PAD));
 sg13g2_IOPadInOut16mA sg13g2_IOPad_io_gpio_0 (.c2p(sg13g2_IOPad_io_gpio_0_c2p),
    .c2p_en(sg13g2_IOPad_io_gpio_0_c2p_en),
    .p2c(sg13g2_IOPad_io_gpio_0_p2c),
    .pad(io_gpio_0_PAD));
 sg13g2_IOPadInOut16mA sg13g2_IOPad_io_gpio_1 (.c2p(sg13g2_IOPad_io_gpio_1_c2p),
    .c2p_en(sg13g2_IOPad_io_gpio_1_c2p_en),
    .p2c(sg13g2_IOPad_io_gpio_1_p2c),
    .pad(io_gpio_1_PAD));
 sg13g2_IOPadInOut16mA sg13g2_IOPad_io_gpio_2 (.c2p(sg13g2_IOPad_io_gpio_2_c2p),
    .c2p_en(sg13g2_IOPad_io_gpio_2_c2p_en),
    .p2c(sg13g2_IOPad_io_gpio_2_p2c),
    .pad(io_gpio_2_PAD));
 sg13g2_IOPadInOut16mA sg13g2_IOPad_io_gpio_3 (.c2p(sg13g2_IOPad_io_gpio_3_c2p),
    .c2p_en(sg13g2_IOPad_io_gpio_3_c2p_en),
    .p2c(sg13g2_IOPad_io_gpio_3_p2c),
    .pad(io_gpio_3_PAD));
 sg13g2_IOPadInOut16mA sg13g2_IOPad_io_gpio_4 (.c2p(sg13g2_IOPad_io_gpio_4_c2p),
    .c2p_en(sg13g2_IOPad_io_gpio_4_c2p_en),
    .p2c(sg13g2_IOPad_io_gpio_4_p2c),
    .pad(io_gpio_4_PAD));
 sg13g2_IOPadInOut16mA sg13g2_IOPad_io_gpio_5 (.c2p(sg13g2_IOPad_io_gpio_5_c2p),
    .c2p_en(sg13g2_IOPad_io_gpio_5_c2p_en),
    .p2c(sg13g2_IOPad_io_gpio_5_p2c),
    .pad(io_gpio_5_PAD));
 sg13g2_IOPadInOut16mA sg13g2_IOPad_io_gpio_6 (.c2p(sg13g2_IOPad_io_gpio_6_c2p),
    .c2p_en(sg13g2_IOPad_io_gpio_6_c2p_en),
    .p2c(sg13g2_IOPad_io_gpio_6_p2c),
    .pad(io_gpio_6_PAD));
 sg13g2_IOPadInOut16mA sg13g2_IOPad_io_gpio_7 (.c2p(sg13g2_IOPad_io_gpio_7_c2p),
    .c2p_en(sg13g2_IOPad_io_gpio_7_c2p_en),
    .p2c(sg13g2_IOPad_io_gpio_7_p2c),
    .pad(io_gpio_7_PAD));
 sg13g2_IOPadOut4mA sg13g2_IOPad_io_i2c_interrupt (.c2p(\system_expander.i2cCtrl_io_i2c_interrupts[0] ),
    .pad(io_i2c_interrupt_PAD));
 sg13g2_IOPadInOut4mA sg13g2_IOPad_io_i2c_scl (.c2p(net),
    .c2p_en(\system_expander.i2cCtrl_io_i2c_scl_write ),
    .p2c(sg13g2_IOPad_io_i2c_scl_p2c),
    .pad(io_i2c_scl_PAD));
 sg13g2_tielo sg13g2_IOPad_io_i2c_scl_1 (.L_LO(net));
 sg13g2_IOPadInOut4mA sg13g2_IOPad_io_i2c_sda (.c2p(net1),
    .c2p_en(\system_expander.i2cCtrl_io_i2c_sda_write ),
    .p2c(sg13g2_IOPad_io_i2c_sda_p2c),
    .pad(io_i2c_sda_PAD));
 sg13g2_tielo sg13g2_IOPad_io_i2c_sda_2 (.L_LO(net1));
 sg13g2_IOPadIn sg13g2_IOPad_io_reset (.p2c(reset),
    .pad(io_reset_PAD));
 sg13g2_dfrbpq_1 \system_expander.gpioConfig_direction[0]$_SDFFE_PN0P_  (.RESET_B(net30),
    .D(_0005_),
    .Q(sg13g2_IOPad_io_gpio_0_c2p_en),
    .CLK(clknet_5_11__leaf_clock_regs));
 sg13g2_tiehi \system_expander.gpioConfig_direction[0]$_SDFFE_PN0P__31  (.L_HI(net30));
 sg13g2_dfrbpq_1 \system_expander.gpioConfig_direction[1]$_SDFFE_PN0P_  (.RESET_B(net31),
    .D(_0006_),
    .Q(sg13g2_IOPad_io_gpio_1_c2p_en),
    .CLK(clknet_5_15__leaf_clock_regs));
 sg13g2_tiehi \system_expander.gpioConfig_direction[1]$_SDFFE_PN0P__32  (.L_HI(net31));
 sg13g2_dfrbpq_1 \system_expander.gpioConfig_direction[2]$_SDFFE_PN0P_  (.RESET_B(net32),
    .D(_0007_),
    .Q(sg13g2_IOPad_io_gpio_2_c2p_en),
    .CLK(clknet_5_30__leaf_clock_regs));
 sg13g2_tiehi \system_expander.gpioConfig_direction[2]$_SDFFE_PN0P__33  (.L_HI(net32));
 sg13g2_dfrbpq_1 \system_expander.gpioConfig_direction[3]$_SDFFE_PN0P_  (.RESET_B(net33),
    .D(_0008_),
    .Q(sg13g2_IOPad_io_gpio_3_c2p_en),
    .CLK(clknet_5_28__leaf_clock_regs));
 sg13g2_tiehi \system_expander.gpioConfig_direction[3]$_SDFFE_PN0P__34  (.L_HI(net33));
 sg13g2_dfrbpq_1 \system_expander.gpioConfig_direction[4]$_SDFFE_PN0P_  (.RESET_B(net34),
    .D(_0009_),
    .Q(sg13g2_IOPad_io_gpio_4_c2p_en),
    .CLK(clknet_5_27__leaf_clock_regs));
 sg13g2_tiehi \system_expander.gpioConfig_direction[4]$_SDFFE_PN0P__35  (.L_HI(net34));
 sg13g2_dfrbpq_1 \system_expander.gpioConfig_direction[5]$_SDFFE_PN0P_  (.RESET_B(net35),
    .D(_0010_),
    .Q(sg13g2_IOPad_io_gpio_5_c2p_en),
    .CLK(clknet_5_1__leaf_clock_regs));
 sg13g2_tiehi \system_expander.gpioConfig_direction[5]$_SDFFE_PN0P__36  (.L_HI(net35));
 sg13g2_dfrbpq_1 \system_expander.gpioConfig_direction[6]$_SDFFE_PN0P_  (.RESET_B(net36),
    .D(_0011_),
    .Q(sg13g2_IOPad_io_gpio_6_c2p_en),
    .CLK(clknet_5_0__leaf_clock_regs));
 sg13g2_tiehi \system_expander.gpioConfig_direction[6]$_SDFFE_PN0P__37  (.L_HI(net36));
 sg13g2_dfrbpq_1 \system_expander.gpioConfig_direction[7]$_SDFFE_PN0P_  (.RESET_B(net37),
    .D(_0012_),
    .Q(sg13g2_IOPad_io_gpio_7_c2p_en),
    .CLK(clknet_5_2__leaf_clock_regs));
 sg13g2_tiehi \system_expander.gpioConfig_direction[7]$_SDFFE_PN0P__38  (.L_HI(net37));
 sg13g2_dfrbpq_1 \system_expander.gpioConfig_write[0]$_SDFFE_PN0P_  (.RESET_B(net38),
    .D(_0013_),
    .Q(sg13g2_IOPad_io_gpio_0_c2p),
    .CLK(clknet_5_11__leaf_clock_regs));
 sg13g2_tiehi \system_expander.gpioConfig_write[0]$_SDFFE_PN0P__39  (.L_HI(net38));
 sg13g2_dfrbpq_1 \system_expander.gpioConfig_write[1]$_SDFFE_PN0P_  (.RESET_B(net39),
    .D(_0014_),
    .Q(sg13g2_IOPad_io_gpio_1_c2p),
    .CLK(clknet_5_15__leaf_clock_regs));
 sg13g2_tiehi \system_expander.gpioConfig_write[1]$_SDFFE_PN0P__40  (.L_HI(net39));
 sg13g2_dfrbpq_1 \system_expander.gpioConfig_write[2]$_SDFFE_PN0P_  (.RESET_B(net40),
    .D(_0015_),
    .Q(sg13g2_IOPad_io_gpio_2_c2p),
    .CLK(clknet_5_30__leaf_clock_regs));
 sg13g2_tiehi \system_expander.gpioConfig_write[2]$_SDFFE_PN0P__41  (.L_HI(net40));
 sg13g2_dfrbpq_1 \system_expander.gpioConfig_write[3]$_SDFFE_PN0P_  (.RESET_B(net41),
    .D(_0016_),
    .Q(sg13g2_IOPad_io_gpio_3_c2p),
    .CLK(clknet_5_30__leaf_clock_regs));
 sg13g2_tiehi \system_expander.gpioConfig_write[3]$_SDFFE_PN0P__42  (.L_HI(net41));
 sg13g2_dfrbpq_1 \system_expander.gpioConfig_write[4]$_SDFFE_PN0P_  (.RESET_B(net42),
    .D(_0017_),
    .Q(sg13g2_IOPad_io_gpio_4_c2p),
    .CLK(clknet_5_27__leaf_clock_regs));
 sg13g2_tiehi \system_expander.gpioConfig_write[4]$_SDFFE_PN0P__43  (.L_HI(net42));
 sg13g2_dfrbpq_1 \system_expander.gpioConfig_write[5]$_SDFFE_PN0P_  (.RESET_B(net43),
    .D(_0018_),
    .Q(sg13g2_IOPad_io_gpio_5_c2p),
    .CLK(clknet_5_0__leaf_clock_regs));
 sg13g2_tiehi \system_expander.gpioConfig_write[5]$_SDFFE_PN0P__44  (.L_HI(net43));
 sg13g2_dfrbpq_1 \system_expander.gpioConfig_write[6]$_SDFFE_PN0P_  (.RESET_B(net44),
    .D(_0019_),
    .Q(sg13g2_IOPad_io_gpio_6_c2p),
    .CLK(clknet_5_0__leaf_clock_regs));
 sg13g2_tiehi \system_expander.gpioConfig_write[6]$_SDFFE_PN0P__45  (.L_HI(net44));
 sg13g2_dfrbpq_1 \system_expander.gpioConfig_write[7]$_SDFFE_PN0P_  (.RESET_B(net45),
    .D(_0020_),
    .Q(sg13g2_IOPad_io_gpio_7_c2p),
    .CLK(clknet_5_8__leaf_clock_regs));
 sg13g2_tiehi \system_expander.gpioConfig_write[7]$_SDFFE_PN0P__46  (.L_HI(net45));
 sg13g2_dfrbpq_1 \system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc/buffers_0[0]$_DFF_P_  (.RESET_B(net152),
    .D(sg13g2_IOPad_io_gpio_0_p2c),
    .Q(\system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[0] ),
    .CLK(clknet_5_11__leaf_clock_regs));
 sg13g2_tiehi \system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc/buffers_0[0]$_DFF_P__153  (.L_HI(net152));
 sg13g2_dfrbpq_1 \system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc/buffers_0[1]$_DFF_P_  (.RESET_B(net153),
    .D(sg13g2_IOPad_io_gpio_1_p2c),
    .Q(\system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[1] ),
    .CLK(clknet_5_24__leaf_clock_regs));
 sg13g2_tiehi \system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc/buffers_0[1]$_DFF_P__154  (.L_HI(net153));
 sg13g2_dfrbpq_1 \system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc/buffers_0[2]$_DFF_P_  (.RESET_B(net154),
    .D(sg13g2_IOPad_io_gpio_2_p2c),
    .Q(\system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[2] ),
    .CLK(clknet_5_31__leaf_clock_regs));
 sg13g2_tiehi \system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc/buffers_0[2]$_DFF_P__155  (.L_HI(net154));
 sg13g2_dfrbpq_1 \system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc/buffers_0[3]$_DFF_P_  (.RESET_B(net155),
    .D(sg13g2_IOPad_io_gpio_3_p2c),
    .Q(\system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[3] ),
    .CLK(clknet_5_31__leaf_clock_regs));
 sg13g2_tiehi \system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc/buffers_0[3]$_DFF_P__156  (.L_HI(net155));
 sg13g2_dfrbpq_1 \system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc/buffers_0[4]$_DFF_P_  (.RESET_B(net156),
    .D(sg13g2_IOPad_io_gpio_4_p2c),
    .Q(\system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[4] ),
    .CLK(clknet_5_31__leaf_clock_regs));
 sg13g2_tiehi \system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc/buffers_0[4]$_DFF_P__157  (.L_HI(net156));
 sg13g2_dfrbpq_1 \system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc/buffers_0[5]$_DFF_P_  (.RESET_B(net157),
    .D(sg13g2_IOPad_io_gpio_5_p2c),
    .Q(\system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[5] ),
    .CLK(clknet_5_0__leaf_clock_regs));
 sg13g2_tiehi \system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc/buffers_0[5]$_DFF_P__158  (.L_HI(net157));
 sg13g2_dfrbpq_1 \system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc/buffers_0[6]$_DFF_P_  (.RESET_B(net158),
    .D(sg13g2_IOPad_io_gpio_6_p2c),
    .Q(\system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[6] ),
    .CLK(clknet_5_3__leaf_clock_regs));
 sg13g2_tiehi \system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc/buffers_0[6]$_DFF_P__159  (.L_HI(net158));
 sg13g2_dfrbpq_1 \system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc/buffers_0[7]$_DFF_P_  (.RESET_B(net159),
    .D(sg13g2_IOPad_io_gpio_7_p2c),
    .Q(\system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[7] ),
    .CLK(clknet_5_8__leaf_clock_regs));
 sg13g2_tiehi \system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc/buffers_0[7]$_DFF_P__160  (.L_HI(net159));
 sg13g2_dfrbpq_1 \system_expander.gpioCtrl_1.last[0]$_DFF_P_  (.RESET_B(net46),
    .D(\system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[0] ),
    .Q(\system_expander.gpioCtrl_1.last[0] ),
    .CLK(clknet_5_14__leaf_clock_regs));
 sg13g2_tiehi \system_expander.gpioCtrl_1.last[0]$_DFF_P__47  (.L_HI(net46));
 sg13g2_dfrbpq_1 \system_expander.gpioCtrl_1.last[1]$_DFF_P_  (.RESET_B(net47),
    .D(\system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[1] ),
    .Q(\system_expander.gpioCtrl_1.last[1] ),
    .CLK(clknet_5_26__leaf_clock_regs));
 sg13g2_tiehi \system_expander.gpioCtrl_1.last[1]$_DFF_P__48  (.L_HI(net47));
 sg13g2_dfrbpq_1 \system_expander.gpioCtrl_1.last[2]$_DFF_P_  (.RESET_B(net48),
    .D(\system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[2] ),
    .Q(\system_expander.gpioCtrl_1.last[2] ),
    .CLK(clknet_5_29__leaf_clock_regs));
 sg13g2_tiehi \system_expander.gpioCtrl_1.last[2]$_DFF_P__49  (.L_HI(net48));
 sg13g2_dfrbpq_1 \system_expander.gpioCtrl_1.last[3]$_DFF_P_  (.RESET_B(net49),
    .D(\system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[3] ),
    .Q(\system_expander.gpioCtrl_1.last[3] ),
    .CLK(clknet_5_23__leaf_clock_regs));
 sg13g2_tiehi \system_expander.gpioCtrl_1.last[3]$_DFF_P__50  (.L_HI(net49));
 sg13g2_dfrbpq_1 \system_expander.gpioCtrl_1.last[4]$_DFF_P_  (.RESET_B(net50),
    .D(\system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[4] ),
    .Q(\system_expander.gpioCtrl_1.last[4] ),
    .CLK(clknet_5_26__leaf_clock_regs));
 sg13g2_tiehi \system_expander.gpioCtrl_1.last[4]$_DFF_P__51  (.L_HI(net50));
 sg13g2_dfrbpq_1 \system_expander.gpioCtrl_1.last[5]$_DFF_P_  (.RESET_B(net51),
    .D(\system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[5] ),
    .Q(\system_expander.gpioCtrl_1.last[5] ),
    .CLK(clknet_5_1__leaf_clock_regs));
 sg13g2_tiehi \system_expander.gpioCtrl_1.last[5]$_DFF_P__52  (.L_HI(net51));
 sg13g2_dfrbpq_1 \system_expander.gpioCtrl_1.last[6]$_DFF_P_  (.RESET_B(net52),
    .D(\system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[6] ),
    .Q(\system_expander.gpioCtrl_1.last[6] ),
    .CLK(clknet_5_3__leaf_clock_regs));
 sg13g2_tiehi \system_expander.gpioCtrl_1.last[6]$_DFF_P__53  (.L_HI(net52));
 sg13g2_dfrbpq_1 \system_expander.gpioCtrl_1.last[7]$_DFF_P_  (.RESET_B(net53),
    .D(\system_expander.gpioCtrl_1.io_gpio_pins_read_buffercc_io_dataOut[7] ),
    .Q(\system_expander.gpioCtrl_1.last[7] ),
    .CLK(clknet_5_8__leaf_clock_regs));
 sg13g2_tiehi \system_expander.gpioCtrl_1.last[7]$_DFF_P__54  (.L_HI(net53));
 sg13g2_dfrbpq_1 \system_expander.i2cConfig_latch$_DFF_P_  (.RESET_B(net54),
    .D(reset),
    .Q(\system_expander.i2cConfig_latch ),
    .CLK(clknet_5_21__leaf_clock_regs));
 sg13g2_tiehi \system_expander.i2cConfig_latch$_DFF_P__55  (.L_HI(net54));
 sg13g2_dfrbpq_1 \system_expander.i2cConfig_latchedAddress[0]$_DFFE_PN_  (.RESET_B(net55),
    .D(_0021_),
    .Q(\system_expander.i2cConfig_latchedAddress[0] ),
    .CLK(clknet_5_21__leaf_clock_regs));
 sg13g2_tiehi \system_expander.i2cConfig_latchedAddress[0]$_DFFE_PN__56  (.L_HI(net55));
 sg13g2_dfrbpq_1 \system_expander.i2cConfig_latchedAddress[1]$_DFFE_PN_  (.RESET_B(net56),
    .D(_0022_),
    .Q(\system_expander.i2cConfig_latchedAddress[1] ),
    .CLK(clknet_5_21__leaf_clock_regs));
 sg13g2_tiehi \system_expander.i2cConfig_latchedAddress[1]$_DFFE_PN__57  (.L_HI(net56));
 sg13g2_dfrbpq_1 \system_expander.i2cConfig_latchedAddress[2]$_DFFE_PN_  (.RESET_B(net57),
    .D(_0023_),
    .Q(\system_expander.i2cConfig_latchedAddress[2] ),
    .CLK(clknet_5_21__leaf_clock_regs));
 sg13g2_tiehi \system_expander.i2cConfig_latchedAddress[2]$_DFFE_PN__58  (.L_HI(net57));
 I2cDeviceCtrl \system_expander.i2cCtrl  (.clock(clknet_1_0__leaf_clock),
    .io_cmd_payload_read(\system_expander.i2cCtrl_io_cmd_payload_read ),
    .io_cmd_payload_reg(\system_expander.i2cCtrl_io_cmd_payload_reg ),
    .io_cmd_ready(\system_expander.i2cCtrl_io_cmd_ready ),
    .io_cmd_valid(\system_expander.i2cCtrl_io_cmd_valid ),
    .io_i2c_scl_read(sg13g2_IOPad_io_i2c_scl_p2c),
    .io_i2c_scl_write(\system_expander.i2cCtrl_io_i2c_scl_write ),
    .io_i2c_sda_read(sg13g2_IOPad_io_i2c_sda_p2c),
    .io_i2c_sda_write(\system_expander.i2cCtrl_io_i2c_sda_write ),
    .io_rsp_payload_error(\system_expander.link_error ),
    .io_rsp_ready(\system_expander.i2cCtrl_io_rsp_ready ),
    .io_rsp_valid(\system_expander.i2cCtrl_io_rsp_valid ),
    .reset(reset),
    .io_cmd_payload_data({\system_expander.i2cCtrl_io_cmd_payload_data[7] ,
    \system_expander.i2cCtrl_io_cmd_payload_data[6] ,
    \system_expander.i2cCtrl_io_cmd_payload_data[5] ,
    \system_expander.i2cCtrl_io_cmd_payload_data[4] ,
    \system_expander.i2cCtrl_io_cmd_payload_data[3] ,
    \system_expander.i2cCtrl_io_cmd_payload_data[2] ,
    \system_expander.i2cCtrl_io_cmd_payload_data[1] ,
    \system_expander.i2cCtrl_io_cmd_payload_data[0] }),
    .io_config_clockDivider({net7,
    net6,
    net5,
    net4,
    net3,
    net2,
    net16,
    net15,
    net14,
    net13,
    net12,
    net11,
    net10,
    net9,
    net8,
    net58}),
    .io_config_deviceAddr({net18,
    net60,
    net59,
    net17,
    \system_expander.i2cConfig_latchedAddress[2] ,
    \system_expander.i2cConfig_latchedAddress[1] ,
    \system_expander.i2cConfig_latchedAddress[0] }),
    .io_config_timeout({net24,
    net23,
    net22,
    net61,
    net21,
    net20,
    net65,
    net64,
    net63,
    net29,
    net28,
    net27,
    net62,
    net26,
    net25,
    net19}),
    .io_i2c_interrupts({\system_expander.i2cCtrl_io_i2c_interrupts[0] }),
    .io_interrupts({\system_expander.i2cCtrl_io_interrupts[0] }),
    .io_rsp_payload_data({\system_expander.link_data[7] ,
    \system_expander.link_data[6] ,
    \system_expander.link_data[5] ,
    \system_expander.link_data[4] ,
    \system_expander.link_data[3] ,
    \system_expander.link_data[2] ,
    \system_expander.link_data[1] ,
    \system_expander.link_data[0] }));
 sg13g2_tielo \system_expander.i2cCtrl_10  (.L_LO(net9));
 sg13g2_tielo \system_expander.i2cCtrl_11  (.L_LO(net10));
 sg13g2_tielo \system_expander.i2cCtrl_12  (.L_LO(net11));
 sg13g2_tielo \system_expander.i2cCtrl_13  (.L_LO(net12));
 sg13g2_tielo \system_expander.i2cCtrl_14  (.L_LO(net13));
 sg13g2_tielo \system_expander.i2cCtrl_15  (.L_LO(net14));
 sg13g2_tielo \system_expander.i2cCtrl_16  (.L_LO(net15));
 sg13g2_tielo \system_expander.i2cCtrl_17  (.L_LO(net16));
 sg13g2_tielo \system_expander.i2cCtrl_18  (.L_LO(net17));
 sg13g2_tielo \system_expander.i2cCtrl_19  (.L_LO(net18));
 sg13g2_tielo \system_expander.i2cCtrl_20  (.L_LO(net19));
 sg13g2_tielo \system_expander.i2cCtrl_21  (.L_LO(net20));
 sg13g2_tielo \system_expander.i2cCtrl_22  (.L_LO(net21));
 sg13g2_tielo \system_expander.i2cCtrl_23  (.L_LO(net22));
 sg13g2_tielo \system_expander.i2cCtrl_24  (.L_LO(net23));
 sg13g2_tielo \system_expander.i2cCtrl_25  (.L_LO(net24));
 sg13g2_tielo \system_expander.i2cCtrl_26  (.L_LO(net25));
 sg13g2_tielo \system_expander.i2cCtrl_27  (.L_LO(net26));
 sg13g2_tielo \system_expander.i2cCtrl_28  (.L_LO(net27));
 sg13g2_tielo \system_expander.i2cCtrl_29  (.L_LO(net28));
 sg13g2_tielo \system_expander.i2cCtrl_3  (.L_LO(net2));
 sg13g2_tielo \system_expander.i2cCtrl_30  (.L_LO(net29));
 sg13g2_tielo \system_expander.i2cCtrl_4  (.L_LO(net3));
 sg13g2_tielo \system_expander.i2cCtrl_5  (.L_LO(net4));
 sg13g2_tiehi \system_expander.i2cCtrl_59  (.L_HI(net58));
 sg13g2_tielo \system_expander.i2cCtrl_6  (.L_LO(net5));
 sg13g2_tiehi \system_expander.i2cCtrl_60  (.L_HI(net59));
 sg13g2_tiehi \system_expander.i2cCtrl_61  (.L_HI(net60));
 sg13g2_tiehi \system_expander.i2cCtrl_62  (.L_HI(net61));
 sg13g2_tiehi \system_expander.i2cCtrl_63  (.L_HI(net62));
 sg13g2_tiehi \system_expander.i2cCtrl_64  (.L_HI(net63));
 sg13g2_tiehi \system_expander.i2cCtrl_65  (.L_HI(net64));
 sg13g2_tiehi \system_expander.i2cCtrl_66  (.L_HI(net65));
 sg13g2_tielo \system_expander.i2cCtrl_7  (.L_LO(net6));
 sg13g2_tielo \system_expander.i2cCtrl_8  (.L_LO(net7));
 sg13g2_tielo \system_expander.i2cCtrl_9  (.L_LO(net8));
 sg13g2_dfrbpq_1 \system_expander.irq_fall_ctrl.pendings[0]$_SDFF_PN0_  (.RESET_B(net66),
    .D(_0024_),
    .Q(\system_expander.irq_fall_ctrl.pendings[0] ),
    .CLK(clknet_5_15__leaf_clock_regs));
 sg13g2_tiehi \system_expander.irq_fall_ctrl.pendings[0]$_SDFF_PN0__67  (.L_HI(net66));
 sg13g2_dfrbpq_1 \system_expander.irq_fall_ctrl.pendings[1]$_SDFF_PN0_  (.RESET_B(net67),
    .D(_0025_),
    .Q(\system_expander.irq_fall_ctrl.pendings[1] ),
    .CLK(clknet_5_24__leaf_clock_regs));
 sg13g2_tiehi \system_expander.irq_fall_ctrl.pendings[1]$_SDFF_PN0__68  (.L_HI(net67));
 sg13g2_dfrbpq_1 \system_expander.irq_fall_ctrl.pendings[2]$_SDFF_PN0_  (.RESET_B(net68),
    .D(_0026_),
    .Q(\system_expander.irq_fall_ctrl.pendings[2] ),
    .CLK(clknet_5_29__leaf_clock_regs));
 sg13g2_tiehi \system_expander.irq_fall_ctrl.pendings[2]$_SDFF_PN0__69  (.L_HI(net68));
 sg13g2_dfrbpq_1 \system_expander.irq_fall_ctrl.pendings[3]$_SDFF_PN0_  (.RESET_B(net69),
    .D(_0027_),
    .Q(\system_expander.irq_fall_ctrl.pendings[3] ),
    .CLK(clknet_5_23__leaf_clock_regs));
 sg13g2_tiehi \system_expander.irq_fall_ctrl.pendings[3]$_SDFF_PN0__70  (.L_HI(net69));
 sg13g2_dfrbpq_1 \system_expander.irq_fall_ctrl.pendings[4]$_SDFF_PN0_  (.RESET_B(net70),
    .D(_0028_),
    .Q(\system_expander.irq_fall_ctrl.pendings[4] ),
    .CLK(clknet_5_26__leaf_clock_regs));
 sg13g2_tiehi \system_expander.irq_fall_ctrl.pendings[4]$_SDFF_PN0__71  (.L_HI(net70));
 sg13g2_dfrbpq_1 \system_expander.irq_fall_ctrl.pendings[5]$_SDFF_PN0_  (.RESET_B(net71),
    .D(_0029_),
    .Q(\system_expander.irq_fall_ctrl.pendings[5] ),
    .CLK(clknet_5_1__leaf_clock_regs));
 sg13g2_tiehi \system_expander.irq_fall_ctrl.pendings[5]$_SDFF_PN0__72  (.L_HI(net71));
 sg13g2_dfrbpq_1 \system_expander.irq_fall_ctrl.pendings[6]$_SDFF_PN0_  (.RESET_B(net72),
    .D(_0030_),
    .Q(\system_expander.irq_fall_ctrl.pendings[6] ),
    .CLK(clknet_5_3__leaf_clock_regs));
 sg13g2_tiehi \system_expander.irq_fall_ctrl.pendings[6]$_SDFF_PN0__73  (.L_HI(net72));
 sg13g2_dfrbpq_1 \system_expander.irq_fall_ctrl.pendings[7]$_SDFF_PN0_  (.RESET_B(net73),
    .D(_0031_),
    .Q(\system_expander.irq_fall_ctrl.pendings[7] ),
    .CLK(clknet_5_2__leaf_clock_regs));
 sg13g2_tiehi \system_expander.irq_fall_ctrl.pendings[7]$_SDFF_PN0__74  (.L_HI(net73));
 sg13g2_dfrbpq_1 \system_expander.irq_fall_masks[0]$_SDFFE_PN0P_  (.RESET_B(net74),
    .D(_0032_),
    .Q(\system_expander.irq_fall_ctrl.io_masks[0] ),
    .CLK(clknet_5_10__leaf_clock_regs));
 sg13g2_tiehi \system_expander.irq_fall_masks[0]$_SDFFE_PN0P__75  (.L_HI(net74));
 sg13g2_dfrbpq_1 \system_expander.irq_fall_masks[1]$_SDFFE_PN0P_  (.RESET_B(net75),
    .D(_0033_),
    .Q(\system_expander.irq_fall_ctrl.io_masks[1] ),
    .CLK(clknet_5_25__leaf_clock_regs));
 sg13g2_tiehi \system_expander.irq_fall_masks[1]$_SDFFE_PN0P__76  (.L_HI(net75));
 sg13g2_dfrbpq_1 \system_expander.irq_fall_masks[2]$_SDFFE_PN0P_  (.RESET_B(net76),
    .D(_0034_),
    .Q(\system_expander.irq_fall_ctrl.io_masks[2] ),
    .CLK(clknet_5_30__leaf_clock_regs));
 sg13g2_tiehi \system_expander.irq_fall_masks[2]$_SDFFE_PN0P__77  (.L_HI(net76));
 sg13g2_dfrbpq_1 \system_expander.irq_fall_masks[3]$_SDFFE_PN0P_  (.RESET_B(net77),
    .D(_0035_),
    .Q(\system_expander.irq_fall_ctrl.io_masks[3] ),
    .CLK(clknet_5_19__leaf_clock_regs));
 sg13g2_tiehi \system_expander.irq_fall_masks[3]$_SDFFE_PN0P__78  (.L_HI(net77));
 sg13g2_dfrbpq_1 \system_expander.irq_fall_masks[4]$_SDFFE_PN0P_  (.RESET_B(net78),
    .D(_0036_),
    .Q(\system_expander.irq_fall_ctrl.io_masks[4] ),
    .CLK(clknet_5_25__leaf_clock_regs));
 sg13g2_tiehi \system_expander.irq_fall_masks[4]$_SDFFE_PN0P__79  (.L_HI(net78));
 sg13g2_dfrbpq_1 \system_expander.irq_fall_masks[5]$_SDFFE_PN0P_  (.RESET_B(net79),
    .D(_0037_),
    .Q(\system_expander.irq_fall_ctrl.io_masks[5] ),
    .CLK(clknet_5_1__leaf_clock_regs));
 sg13g2_tiehi \system_expander.irq_fall_masks[5]$_SDFFE_PN0P__80  (.L_HI(net79));
 sg13g2_dfrbpq_1 \system_expander.irq_fall_masks[6]$_SDFFE_PN0P_  (.RESET_B(net80),
    .D(_0038_),
    .Q(\system_expander.irq_fall_ctrl.io_masks[6] ),
    .CLK(clknet_5_3__leaf_clock_regs));
 sg13g2_tiehi \system_expander.irq_fall_masks[6]$_SDFFE_PN0P__81  (.L_HI(net80));
 sg13g2_dfrbpq_1 \system_expander.irq_fall_masks[7]$_SDFFE_PN0P_  (.RESET_B(net81),
    .D(_0039_),
    .Q(\system_expander.irq_fall_ctrl.io_masks[7] ),
    .CLK(clknet_5_2__leaf_clock_regs));
 sg13g2_tiehi \system_expander.irq_fall_masks[7]$_SDFFE_PN0P__82  (.L_HI(net81));
 sg13g2_dfrbpq_1 \system_expander.irq_high_ctrl.pendings[0]$_SDFF_PN0_  (.RESET_B(net82),
    .D(_0040_),
    .Q(\system_expander.irq_high_ctrl.pendings[0] ),
    .CLK(clknet_5_14__leaf_clock_regs));
 sg13g2_tiehi \system_expander.irq_high_ctrl.pendings[0]$_SDFF_PN0__83  (.L_HI(net82));
 sg13g2_dfrbpq_1 \system_expander.irq_high_ctrl.pendings[1]$_SDFF_PN0_  (.RESET_B(net83),
    .D(_0041_),
    .Q(\system_expander.irq_high_ctrl.pendings[1] ),
    .CLK(clknet_5_12__leaf_clock_regs));
 sg13g2_tiehi \system_expander.irq_high_ctrl.pendings[1]$_SDFF_PN0__84  (.L_HI(net83));
 sg13g2_dfrbpq_1 \system_expander.irq_high_ctrl.pendings[2]$_SDFF_PN0_  (.RESET_B(net84),
    .D(_0042_),
    .Q(\system_expander.irq_high_ctrl.pendings[2] ),
    .CLK(clknet_5_28__leaf_clock_regs));
 sg13g2_tiehi \system_expander.irq_high_ctrl.pendings[2]$_SDFF_PN0__85  (.L_HI(net84));
 sg13g2_dfrbpq_1 \system_expander.irq_high_ctrl.pendings[3]$_SDFF_PN0_  (.RESET_B(net85),
    .D(_0043_),
    .Q(\system_expander.irq_high_ctrl.pendings[3] ),
    .CLK(clknet_5_28__leaf_clock_regs));
 sg13g2_tiehi \system_expander.irq_high_ctrl.pendings[3]$_SDFF_PN0__86  (.L_HI(net85));
 sg13g2_dfrbpq_1 \system_expander.irq_high_ctrl.pendings[4]$_SDFF_PN0_  (.RESET_B(net86),
    .D(_0044_),
    .Q(\system_expander.irq_high_ctrl.pendings[4] ),
    .CLK(clknet_5_18__leaf_clock_regs));
 sg13g2_tiehi \system_expander.irq_high_ctrl.pendings[4]$_SDFF_PN0__87  (.L_HI(net86));
 sg13g2_dfrbpq_1 \system_expander.irq_high_ctrl.pendings[5]$_SDFF_PN0_  (.RESET_B(net87),
    .D(_0045_),
    .Q(\system_expander.irq_high_ctrl.pendings[5] ),
    .CLK(clknet_5_6__leaf_clock_regs));
 sg13g2_tiehi \system_expander.irq_high_ctrl.pendings[5]$_SDFF_PN0__88  (.L_HI(net87));
 sg13g2_dfrbpq_1 \system_expander.irq_high_ctrl.pendings[6]$_SDFF_PN0_  (.RESET_B(net88),
    .D(_0046_),
    .Q(\system_expander.irq_high_ctrl.pendings[6] ),
    .CLK(clknet_5_6__leaf_clock_regs));
 sg13g2_tiehi \system_expander.irq_high_ctrl.pendings[6]$_SDFF_PN0__89  (.L_HI(net88));
 sg13g2_dfrbpq_1 \system_expander.irq_high_ctrl.pendings[7]$_SDFF_PN0_  (.RESET_B(net89),
    .D(_0047_),
    .Q(\system_expander.irq_high_ctrl.pendings[7] ),
    .CLK(clknet_5_10__leaf_clock_regs));
 sg13g2_tiehi \system_expander.irq_high_ctrl.pendings[7]$_SDFF_PN0__90  (.L_HI(net89));
 sg13g2_dfrbpq_1 \system_expander.irq_high_masks[0]$_SDFFE_PN0P_  (.RESET_B(net90),
    .D(_0048_),
    .Q(\system_expander.irq_high_ctrl.io_masks[0] ),
    .CLK(clknet_5_14__leaf_clock_regs));
 sg13g2_tiehi \system_expander.irq_high_masks[0]$_SDFFE_PN0P__91  (.L_HI(net90));
 sg13g2_dfrbpq_1 \system_expander.irq_high_masks[1]$_SDFFE_PN0P_  (.RESET_B(net91),
    .D(_0049_),
    .Q(\system_expander.irq_high_ctrl.io_masks[1] ),
    .CLK(clknet_5_12__leaf_clock_regs));
 sg13g2_tiehi \system_expander.irq_high_masks[1]$_SDFFE_PN0P__92  (.L_HI(net91));
 sg13g2_dfrbpq_1 \system_expander.irq_high_masks[2]$_SDFFE_PN0P_  (.RESET_B(net92),
    .D(_0050_),
    .Q(\system_expander.irq_high_ctrl.io_masks[2] ),
    .CLK(clknet_5_27__leaf_clock_regs));
 sg13g2_tiehi \system_expander.irq_high_masks[2]$_SDFFE_PN0P__93  (.L_HI(net92));
 sg13g2_dfrbpq_1 \system_expander.irq_high_masks[3]$_SDFFE_PN0P_  (.RESET_B(net93),
    .D(_0051_),
    .Q(\system_expander.irq_high_ctrl.io_masks[3] ),
    .CLK(clknet_5_25__leaf_clock_regs));
 sg13g2_tiehi \system_expander.irq_high_masks[3]$_SDFFE_PN0P__94  (.L_HI(net93));
 sg13g2_dfrbpq_1 \system_expander.irq_high_masks[4]$_SDFFE_PN0P_  (.RESET_B(net94),
    .D(_0052_),
    .Q(\system_expander.irq_high_ctrl.io_masks[4] ),
    .CLK(clknet_5_24__leaf_clock_regs));
 sg13g2_tiehi \system_expander.irq_high_masks[4]$_SDFFE_PN0P__95  (.L_HI(net94));
 sg13g2_dfrbpq_1 \system_expander.irq_high_masks[5]$_SDFFE_PN0P_  (.RESET_B(net95),
    .D(_0053_),
    .Q(\system_expander.irq_high_ctrl.io_masks[5] ),
    .CLK(clknet_5_9__leaf_clock_regs));
 sg13g2_tiehi \system_expander.irq_high_masks[5]$_SDFFE_PN0P__96  (.L_HI(net95));
 sg13g2_dfrbpq_1 \system_expander.irq_high_masks[6]$_SDFFE_PN0P_  (.RESET_B(net96),
    .D(_0054_),
    .Q(\system_expander.irq_high_ctrl.io_masks[6] ),
    .CLK(clknet_5_9__leaf_clock_regs));
 sg13g2_tiehi \system_expander.irq_high_masks[6]$_SDFFE_PN0P__97  (.L_HI(net96));
 sg13g2_dfrbpq_1 \system_expander.irq_high_masks[7]$_SDFFE_PN0P_  (.RESET_B(net97),
    .D(_0055_),
    .Q(\system_expander.irq_high_ctrl.io_masks[7] ),
    .CLK(clknet_5_9__leaf_clock_regs));
 sg13g2_tiehi \system_expander.irq_high_masks[7]$_SDFFE_PN0P__98  (.L_HI(net97));
 sg13g2_dfrbpq_1 \system_expander.irq_low_ctrl.pendings[0]$_SDFF_PN0_  (.RESET_B(net98),
    .D(_0056_),
    .Q(\system_expander.irq_low_ctrl.pendings[0] ),
    .CLK(clknet_5_12__leaf_clock_regs));
 sg13g2_tiehi \system_expander.irq_low_ctrl.pendings[0]$_SDFF_PN0__99  (.L_HI(net98));
 sg13g2_dfrbpq_1 \system_expander.irq_low_ctrl.pendings[1]$_SDFF_PN0_  (.RESET_B(net99),
    .D(_0057_),
    .Q(\system_expander.irq_low_ctrl.pendings[1] ),
    .CLK(clknet_5_24__leaf_clock_regs));
 sg13g2_tiehi \system_expander.irq_low_ctrl.pendings[1]$_SDFF_PN0__100  (.L_HI(net99));
 sg13g2_dfrbpq_1 \system_expander.irq_low_ctrl.pendings[2]$_SDFF_PN0_  (.RESET_B(net100),
    .D(_0058_),
    .Q(\system_expander.irq_low_ctrl.pendings[2] ),
    .CLK(clknet_5_29__leaf_clock_regs));
 sg13g2_tiehi \system_expander.irq_low_ctrl.pendings[2]$_SDFF_PN0__101  (.L_HI(net100));
 sg13g2_dfrbpq_1 \system_expander.irq_low_ctrl.pendings[3]$_SDFF_PN0_  (.RESET_B(net101),
    .D(_0059_),
    .Q(\system_expander.irq_low_ctrl.pendings[3] ),
    .CLK(clknet_5_22__leaf_clock_regs));
 sg13g2_tiehi \system_expander.irq_low_ctrl.pendings[3]$_SDFF_PN0__102  (.L_HI(net101));
 sg13g2_dfrbpq_1 \system_expander.irq_low_ctrl.pendings[4]$_SDFF_PN0_  (.RESET_B(net102),
    .D(_0060_),
    .Q(\system_expander.irq_low_ctrl.pendings[4] ),
    .CLK(clknet_5_19__leaf_clock_regs));
 sg13g2_tiehi \system_expander.irq_low_ctrl.pendings[4]$_SDFF_PN0__103  (.L_HI(net102));
 sg13g2_dfrbpq_1 \system_expander.irq_low_ctrl.pendings[5]$_SDFF_PN0_  (.RESET_B(net103),
    .D(_0061_),
    .Q(\system_expander.irq_low_ctrl.pendings[5] ),
    .CLK(clknet_5_6__leaf_clock_regs));
 sg13g2_tiehi \system_expander.irq_low_ctrl.pendings[5]$_SDFF_PN0__104  (.L_HI(net103));
 sg13g2_dfrbpq_1 \system_expander.irq_low_ctrl.pendings[6]$_SDFF_PN0_  (.RESET_B(net104),
    .D(_0062_),
    .Q(\system_expander.irq_low_ctrl.pendings[6] ),
    .CLK(clknet_5_6__leaf_clock_regs));
 sg13g2_tiehi \system_expander.irq_low_ctrl.pendings[6]$_SDFF_PN0__105  (.L_HI(net104));
 sg13g2_dfrbpq_1 \system_expander.irq_low_ctrl.pendings[7]$_SDFF_PN0_  (.RESET_B(net105),
    .D(_0063_),
    .Q(\system_expander.irq_low_ctrl.pendings[7] ),
    .CLK(clknet_5_8__leaf_clock_regs));
 sg13g2_tiehi \system_expander.irq_low_ctrl.pendings[7]$_SDFF_PN0__106  (.L_HI(net105));
 sg13g2_dfrbpq_1 \system_expander.irq_low_masks[0]$_SDFFE_PN0P_  (.RESET_B(net106),
    .D(_0064_),
    .Q(\system_expander.irq_low_ctrl.io_masks[0] ),
    .CLK(clknet_5_5__leaf_clock_regs));
 sg13g2_tiehi \system_expander.irq_low_masks[0]$_SDFFE_PN0P__107  (.L_HI(net106));
 sg13g2_dfrbpq_1 \system_expander.irq_low_masks[1]$_SDFFE_PN0P_  (.RESET_B(net107),
    .D(_0065_),
    .Q(\system_expander.irq_low_ctrl.io_masks[1] ),
    .CLK(clknet_5_13__leaf_clock_regs));
 sg13g2_tiehi \system_expander.irq_low_masks[1]$_SDFFE_PN0P__108  (.L_HI(net107));
 sg13g2_dfrbpq_1 \system_expander.irq_low_masks[2]$_SDFFE_PN0P_  (.RESET_B(net108),
    .D(_0066_),
    .Q(\system_expander.irq_low_ctrl.io_masks[2] ),
    .CLK(clknet_5_22__leaf_clock_regs));
 sg13g2_tiehi \system_expander.irq_low_masks[2]$_SDFFE_PN0P__109  (.L_HI(net108));
 sg13g2_dfrbpq_1 \system_expander.irq_low_masks[3]$_SDFFE_PN0P_  (.RESET_B(net109),
    .D(_0067_),
    .Q(\system_expander.irq_low_ctrl.io_masks[3] ),
    .CLK(clknet_5_22__leaf_clock_regs));
 sg13g2_tiehi \system_expander.irq_low_masks[3]$_SDFFE_PN0P__110  (.L_HI(net109));
 sg13g2_dfrbpq_1 \system_expander.irq_low_masks[4]$_SDFFE_PN0P_  (.RESET_B(net110),
    .D(_0068_),
    .Q(\system_expander.irq_low_ctrl.io_masks[4] ),
    .CLK(clknet_5_18__leaf_clock_regs));
 sg13g2_tiehi \system_expander.irq_low_masks[4]$_SDFFE_PN0P__111  (.L_HI(net110));
 sg13g2_dfrbpq_1 \system_expander.irq_low_masks[5]$_SDFFE_PN0P_  (.RESET_B(net111),
    .D(_0069_),
    .Q(\system_expander.irq_low_ctrl.io_masks[5] ),
    .CLK(clknet_5_5__leaf_clock_regs));
 sg13g2_tiehi \system_expander.irq_low_masks[5]$_SDFFE_PN0P__112  (.L_HI(net111));
 sg13g2_dfrbpq_1 \system_expander.irq_low_masks[6]$_SDFFE_PN0P_  (.RESET_B(net112),
    .D(_0070_),
    .Q(\system_expander.irq_low_ctrl.io_masks[6] ),
    .CLK(clknet_5_5__leaf_clock_regs));
 sg13g2_tiehi \system_expander.irq_low_masks[6]$_SDFFE_PN0P__113  (.L_HI(net112));
 sg13g2_dfrbpq_1 \system_expander.irq_low_masks[7]$_SDFFE_PN0P_  (.RESET_B(net113),
    .D(_0071_),
    .Q(\system_expander.irq_low_ctrl.io_masks[7] ),
    .CLK(clknet_5_13__leaf_clock_regs));
 sg13g2_tiehi \system_expander.irq_low_masks[7]$_SDFFE_PN0P__114  (.L_HI(net113));
 sg13g2_dfrbpq_1 \system_expander.irq_rise_ctrl.pendings[0]$_SDFF_PN0_  (.RESET_B(net114),
    .D(_0072_),
    .Q(\system_expander.irq_rise_ctrl.pendings[0] ),
    .CLK(clknet_5_14__leaf_clock_regs));
 sg13g2_tiehi \system_expander.irq_rise_ctrl.pendings[0]$_SDFF_PN0__115  (.L_HI(net114));
 sg13g2_dfrbpq_1 \system_expander.irq_rise_ctrl.pendings[1]$_SDFF_PN0_  (.RESET_B(net115),
    .D(_0073_),
    .Q(\system_expander.irq_rise_ctrl.pendings[1] ),
    .CLK(clknet_5_26__leaf_clock_regs));
 sg13g2_tiehi \system_expander.irq_rise_ctrl.pendings[1]$_SDFF_PN0__116  (.L_HI(net115));
 sg13g2_dfrbpq_1 \system_expander.irq_rise_ctrl.pendings[2]$_SDFF_PN0_  (.RESET_B(net116),
    .D(_0074_),
    .Q(\system_expander.irq_rise_ctrl.pendings[2] ),
    .CLK(clknet_5_29__leaf_clock_regs));
 sg13g2_tiehi \system_expander.irq_rise_ctrl.pendings[2]$_SDFF_PN0__117  (.L_HI(net116));
 sg13g2_dfrbpq_1 \system_expander.irq_rise_ctrl.pendings[3]$_SDFF_PN0_  (.RESET_B(net117),
    .D(_0075_),
    .Q(\system_expander.irq_rise_ctrl.pendings[3] ),
    .CLK(clknet_5_23__leaf_clock_regs));
 sg13g2_tiehi \system_expander.irq_rise_ctrl.pendings[3]$_SDFF_PN0__118  (.L_HI(net117));
 sg13g2_dfrbpq_1 \system_expander.irq_rise_ctrl.pendings[4]$_SDFF_PN0_  (.RESET_B(net118),
    .D(_0076_),
    .Q(\system_expander.irq_rise_ctrl.pendings[4] ),
    .CLK(clknet_5_25__leaf_clock_regs));
 sg13g2_tiehi \system_expander.irq_rise_ctrl.pendings[4]$_SDFF_PN0__119  (.L_HI(net118));
 sg13g2_dfrbpq_1 \system_expander.irq_rise_ctrl.pendings[5]$_SDFF_PN0_  (.RESET_B(net119),
    .D(_0077_),
    .Q(\system_expander.irq_rise_ctrl.pendings[5] ),
    .CLK(clknet_5_7__leaf_clock_regs));
 sg13g2_tiehi \system_expander.irq_rise_ctrl.pendings[5]$_SDFF_PN0__120  (.L_HI(net119));
 sg13g2_dfrbpq_1 \system_expander.irq_rise_ctrl.pendings[6]$_SDFF_PN0_  (.RESET_B(net120),
    .D(_0078_),
    .Q(\system_expander.irq_rise_ctrl.pendings[6] ),
    .CLK(clknet_5_2__leaf_clock_regs));
 sg13g2_tiehi \system_expander.irq_rise_ctrl.pendings[6]$_SDFF_PN0__121  (.L_HI(net120));
 sg13g2_dfrbpq_1 \system_expander.irq_rise_ctrl.pendings[7]$_SDFF_PN0_  (.RESET_B(net121),
    .D(_0079_),
    .Q(\system_expander.irq_rise_ctrl.pendings[7] ),
    .CLK(clknet_5_10__leaf_clock_regs));
 sg13g2_tiehi \system_expander.irq_rise_ctrl.pendings[7]$_SDFF_PN0__122  (.L_HI(net121));
 sg13g2_dfrbpq_1 \system_expander.irq_rise_masks[0]$_SDFFE_PN0P_  (.RESET_B(net122),
    .D(_0080_),
    .Q(\system_expander.irq_rise_ctrl.io_masks[0] ),
    .CLK(clknet_5_10__leaf_clock_regs));
 sg13g2_tiehi \system_expander.irq_rise_masks[0]$_SDFFE_PN0P__123  (.L_HI(net122));
 sg13g2_dfrbpq_1 \system_expander.irq_rise_masks[1]$_SDFFE_PN0P_  (.RESET_B(net123),
    .D(_0081_),
    .Q(\system_expander.irq_rise_ctrl.io_masks[1] ),
    .CLK(clknet_5_13__leaf_clock_regs));
 sg13g2_tiehi \system_expander.irq_rise_masks[1]$_SDFFE_PN0P__124  (.L_HI(net123));
 sg13g2_dfrbpq_1 \system_expander.irq_rise_masks[2]$_SDFFE_PN0P_  (.RESET_B(net124),
    .D(_0082_),
    .Q(\system_expander.irq_rise_ctrl.io_masks[2] ),
    .CLK(clknet_5_28__leaf_clock_regs));
 sg13g2_tiehi \system_expander.irq_rise_masks[2]$_SDFFE_PN0P__125  (.L_HI(net124));
 sg13g2_dfrbpq_1 \system_expander.irq_rise_masks[3]$_SDFFE_PN0P_  (.RESET_B(net125),
    .D(_0083_),
    .Q(\system_expander.irq_rise_ctrl.io_masks[3] ),
    .CLK(clknet_5_22__leaf_clock_regs));
 sg13g2_tiehi \system_expander.irq_rise_masks[3]$_SDFFE_PN0P__126  (.L_HI(net125));
 sg13g2_dfrbpq_1 \system_expander.irq_rise_masks[4]$_SDFFE_PN0P_  (.RESET_B(net126),
    .D(_0084_),
    .Q(\system_expander.irq_rise_ctrl.io_masks[4] ),
    .CLK(clknet_5_18__leaf_clock_regs));
 sg13g2_tiehi \system_expander.irq_rise_masks[4]$_SDFFE_PN0P__127  (.L_HI(net126));
 sg13g2_dfrbpq_1 \system_expander.irq_rise_masks[5]$_SDFFE_PN0P_  (.RESET_B(net127),
    .D(_0085_),
    .Q(\system_expander.irq_rise_ctrl.io_masks[5] ),
    .CLK(clknet_5_7__leaf_clock_regs));
 sg13g2_tiehi \system_expander.irq_rise_masks[5]$_SDFFE_PN0P__128  (.L_HI(net127));
 sg13g2_dfrbpq_1 \system_expander.irq_rise_masks[6]$_SDFFE_PN0P_  (.RESET_B(net128),
    .D(_0086_),
    .Q(\system_expander.irq_rise_ctrl.io_masks[6] ),
    .CLK(clknet_5_5__leaf_clock_regs));
 sg13g2_tiehi \system_expander.irq_rise_masks[6]$_SDFFE_PN0P__129  (.L_HI(net128));
 sg13g2_dfrbpq_1 \system_expander.irq_rise_masks[7]$_SDFFE_PN0P_  (.RESET_B(net129),
    .D(_0087_),
    .Q(\system_expander.irq_rise_ctrl.io_masks[7] ),
    .CLK(clknet_5_9__leaf_clock_regs));
 sg13g2_tiehi \system_expander.irq_rise_masks[7]$_SDFFE_PN0P__130  (.L_HI(net129));
 sg13g2_dfrbpq_1 \system_expander.link_data[0]$_SDFFE_PN0P_  (.RESET_B(net130),
    .D(_0088_),
    .Q(\system_expander.link_data[0] ),
    .CLK(clknet_5_12__leaf_clock_regs));
 sg13g2_tiehi \system_expander.link_data[0]$_SDFFE_PN0P__131  (.L_HI(net130));
 sg13g2_dfrbpq_1 \system_expander.link_data[1]$_SDFFE_PN0P_  (.RESET_B(net131),
    .D(_0089_),
    .Q(\system_expander.link_data[1] ),
    .CLK(clknet_5_18__leaf_clock_regs));
 sg13g2_tiehi \system_expander.link_data[1]$_SDFFE_PN0P__132  (.L_HI(net131));
 sg13g2_dfrbpq_1 \system_expander.link_data[2]$_SDFFE_PN0P_  (.RESET_B(net132),
    .D(_0090_),
    .Q(\system_expander.link_data[2] ),
    .CLK(clknet_5_19__leaf_clock_regs));
 sg13g2_tiehi \system_expander.link_data[2]$_SDFFE_PN0P__133  (.L_HI(net132));
 sg13g2_dfrbpq_1 \system_expander.link_data[3]$_SDFFE_PN0P_  (.RESET_B(net133),
    .D(_0091_),
    .Q(\system_expander.link_data[3] ),
    .CLK(clknet_5_17__leaf_clock_regs));
 sg13g2_tiehi \system_expander.link_data[3]$_SDFFE_PN0P__134  (.L_HI(net133));
 sg13g2_dfrbpq_1 \system_expander.link_data[4]$_SDFFE_PN0P_  (.RESET_B(net134),
    .D(_0092_),
    .Q(\system_expander.link_data[4] ),
    .CLK(clknet_5_19__leaf_clock_regs));
 sg13g2_tiehi \system_expander.link_data[4]$_SDFFE_PN0P__135  (.L_HI(net134));
 sg13g2_dfrbpq_1 \system_expander.link_data[5]$_SDFFE_PN0P_  (.RESET_B(net135),
    .D(_0093_),
    .Q(\system_expander.link_data[5] ),
    .CLK(clknet_5_7__leaf_clock_regs));
 sg13g2_tiehi \system_expander.link_data[5]$_SDFFE_PN0P__136  (.L_HI(net135));
 sg13g2_dfrbpq_1 \system_expander.link_data[6]$_SDFFE_PN0P_  (.RESET_B(net136),
    .D(_0094_),
    .Q(\system_expander.link_data[6] ),
    .CLK(clknet_5_4__leaf_clock_regs));
 sg13g2_tiehi \system_expander.link_data[6]$_SDFFE_PN0P__137  (.L_HI(net136));
 sg13g2_dfrbpq_1 \system_expander.link_data[7]$_SDFFE_PN0P_  (.RESET_B(net137),
    .D(_0095_),
    .Q(\system_expander.link_data[7] ),
    .CLK(clknet_5_13__leaf_clock_regs));
 sg13g2_tiehi \system_expander.link_data[7]$_SDFFE_PN0P__138  (.L_HI(net137));
 sg13g2_dfrbpq_1 \system_expander.link_error$_SDFFE_PN0P_  (.RESET_B(net138),
    .D(_0096_),
    .Q(\system_expander.link_error ),
    .CLK(clknet_5_4__leaf_clock_regs));
 sg13g2_tiehi \system_expander.link_error$_SDFFE_PN0P__139  (.L_HI(net138));
 sg13g2_dfrbpq_1 \system_expander.link_regAddr[0]$_DFFE_PP_  (.RESET_B(net139),
    .D(_0097_),
    .Q(\system_expander.link_regAddr[0] ),
    .CLK(clknet_5_17__leaf_clock_regs));
 sg13g2_tiehi \system_expander.link_regAddr[0]$_DFFE_PP__140  (.L_HI(net139));
 sg13g2_dfrbpq_1 \system_expander.link_regAddr[1]$_DFFE_PP_  (.RESET_B(net140),
    .D(_0098_),
    .Q(\system_expander.link_regAddr[1] ),
    .CLK(clknet_5_16__leaf_clock_regs));
 sg13g2_tiehi \system_expander.link_regAddr[1]$_DFFE_PP__141  (.L_HI(net140));
 sg13g2_dfrbpq_1 \system_expander.link_regAddr[2]$_DFFE_PP_  (.RESET_B(net141),
    .D(_0099_),
    .Q(\system_expander.link_regAddr[2] ),
    .CLK(clknet_5_17__leaf_clock_regs));
 sg13g2_tiehi \system_expander.link_regAddr[2]$_DFFE_PP__142  (.L_HI(net141));
 sg13g2_dfrbpq_1 \system_expander.link_regAddr[3]$_DFFE_PP_  (.RESET_B(net142),
    .D(_0100_),
    .Q(\system_expander.link_regAddr[3] ),
    .CLK(clknet_5_17__leaf_clock_regs));
 sg13g2_tiehi \system_expander.link_regAddr[3]$_DFFE_PP__143  (.L_HI(net142));
 sg13g2_dfrbpq_1 \system_expander.link_regAddr[4]$_DFFE_PP_  (.RESET_B(net143),
    .D(_0101_),
    .Q(\system_expander.link_regAddr[4] ),
    .CLK(clknet_5_20__leaf_clock_regs));
 sg13g2_tiehi \system_expander.link_regAddr[4]$_DFFE_PP__144  (.L_HI(net143));
 sg13g2_dfrbpq_1 \system_expander.link_regAddr[5]$_DFFE_PP_  (.RESET_B(net144),
    .D(_0102_),
    .Q(\system_expander.link_regAddr[5] ),
    .CLK(clknet_5_20__leaf_clock_regs));
 sg13g2_tiehi \system_expander.link_regAddr[5]$_DFFE_PP__145  (.L_HI(net144));
 sg13g2_dfrbpq_1 \system_expander.link_regAddr[6]$_DFFE_PP_  (.RESET_B(net145),
    .D(_0103_),
    .Q(\system_expander.link_regAddr[6] ),
    .CLK(clknet_5_20__leaf_clock_regs));
 sg13g2_tiehi \system_expander.link_regAddr[6]$_DFFE_PP__146  (.L_HI(net145));
 sg13g2_dfrbpq_1 \system_expander.link_regAddr[7]$_DFFE_PP_  (.RESET_B(net146),
    .D(_0104_),
    .Q(\system_expander.link_regAddr[7] ),
    .CLK(clknet_5_20__leaf_clock_regs));
 sg13g2_tiehi \system_expander.link_regAddr[7]$_DFFE_PP__147  (.L_HI(net146));
 sg13g2_dfrbpq_1 \system_expander.link_state[0]$_DFF_P_  (.RESET_B(net147),
    .D(_0003_),
    .Q(\system_expander.link_state[0] ),
    .CLK(clknet_5_4__leaf_clock_regs));
 sg13g2_tiehi \system_expander.link_state[0]$_DFF_P__148  (.L_HI(net147));
 sg13g2_dfrbpq_1 \system_expander.link_state[1]$_DFF_P_  (.RESET_B(net148),
    .D(_0004_),
    .Q(\system_expander.link_state[1] ),
    .CLK(clknet_5_4__leaf_clock_regs));
 sg13g2_tiehi \system_expander.link_state[1]$_DFF_P__149  (.L_HI(net148));
 sg13g2_dfrbpq_1 \system_expander.link_state[2]$_DFF_P_  (.RESET_B(net149),
    .D(_0000_),
    .Q(\system_expander.link_state[2] ),
    .CLK(clknet_5_16__leaf_clock_regs));
 sg13g2_tiehi \system_expander.link_state[2]$_DFF_P__150  (.L_HI(net149));
 sg13g2_dfrbpq_1 \system_expander.link_state[3]$_DFF_P_  (.RESET_B(net150),
    .D(_0001_),
    .Q(\system_expander.link_state[3] ),
    .CLK(clknet_5_16__leaf_clock_regs));
 sg13g2_tiehi \system_expander.link_state[3]$_DFF_P__151  (.L_HI(net150));
 sg13g2_dfrbpq_1 \system_expander.link_state[4]$_DFF_P_  (.RESET_B(net151),
    .D(_0002_),
    .Q(\system_expander.link_state[4] ),
    .CLK(clknet_5_16__leaf_clock_regs));
 sg13g2_tiehi \system_expander.link_state[4]$_DFF_P__152  (.L_HI(net151));
endmodule
