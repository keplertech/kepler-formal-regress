module I2cDeviceCtrl (clock,
    io_cmd_payload_read,
    io_cmd_payload_reg,
    io_cmd_ready,
    io_cmd_valid,
    io_i2c_scl_read,
    io_i2c_scl_write,
    io_i2c_sda_read,
    io_i2c_sda_write,
    io_rsp_payload_error,
    io_rsp_ready,
    io_rsp_valid,
    reset,
    io_cmd_payload_data,
    io_config_clockDivider,
    io_config_deviceAddr,
    io_config_timeout,
    io_i2c_interrupts,
    io_interrupts,
    io_rsp_payload_data);
 input clock;
 output io_cmd_payload_read;
 output io_cmd_payload_reg;
 input io_cmd_ready;
 output io_cmd_valid;
 input io_i2c_scl_read;
 output io_i2c_scl_write;
 input io_i2c_sda_read;
 output io_i2c_sda_write;
 input io_rsp_payload_error;
 output io_rsp_ready;
 input io_rsp_valid;
 input reset;
 output [7:0] io_cmd_payload_data;
 input [15:0] io_config_clockDivider;
 input [6:0] io_config_deviceAddr;
 input [15:0] io_config_timeout;
 output [0:0] io_i2c_interrupts;
 input [0:0] io_interrupts;
 input [7:0] io_rsp_payload_data;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _076_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _083_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _089_;
 wire _091_;
 wire _093_;
 wire _094_;
 wire _096_;
 wire _097_;
 wire _099_;
 wire _101_;
 wire _102_;
 wire _104_;
 wire _105_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _112_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _137_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _205_;
 wire _206_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _297_;
 wire _298_;
 wire _300_;
 wire _301_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire net75;
 wire net1;
 wire \_zz_ctrl_sdaWrite[0] ;
 wire \_zz_ctrl_sdaWrite[1] ;
 wire \_zz_ctrl_sdaWrite[2] ;
 wire \_zz_ctrl_sdaWrite[3] ;
 wire \_zz_ctrl_sdaWrite[4] ;
 wire \_zz_ctrl_sdaWrite[5] ;
 wire \_zz_ctrl_sdaWrite[6] ;
 wire \_zz_ctrl_sdaWrite[7] ;
 wire \_zz_ctrl_sdaWrite_1[0] ;
 wire \_zz_ctrl_sdaWrite_1[1] ;
 wire \_zz_ctrl_sdaWrite_1[2] ;
 wire _zz_filter_sampler_sclSamples_0;
 wire _zz_filter_sampler_sclSamples_1;
 wire _zz_filter_sampler_sclSamples_2;
 wire _zz_filter_sampler_sdaSamples_0;
 wire _zz_filter_sampler_sdaSamples_1;
 wire _zz_filter_sampler_sdaSamples_2;
 wire \ctrl_bitCounter[3] ;
 wire \ctrl_bitCounter[4] ;
 wire ctrl_cmdLock;
 wire \ctrl_frameCounter[0] ;
 wire \ctrl_frameCounter[1] ;
 wire \ctrl_frameCounter[2] ;
 wire \ctrl_frameCounter[3] ;
 wire ctrl_response_error;
 wire \ctrl_state[0] ;
 wire \ctrl_state[1] ;
 wire ctrl_transmission;
 wire filter_scl;
 wire filter_scl_regNext;
 wire filter_sda;
 wire filter_sda_regNext;
 wire \filter_timer_counter[0] ;
 wire \filter_timer_counter[10] ;
 wire \filter_timer_counter[11] ;
 wire \filter_timer_counter[12] ;
 wire \filter_timer_counter[13] ;
 wire \filter_timer_counter[14] ;
 wire \filter_timer_counter[15] ;
 wire \filter_timer_counter[1] ;
 wire \filter_timer_counter[2] ;
 wire \filter_timer_counter[3] ;
 wire \filter_timer_counter[4] ;
 wire \filter_timer_counter[5] ;
 wire \filter_timer_counter[6] ;
 wire \filter_timer_counter[7] ;
 wire \filter_timer_counter[8] ;
 wire \filter_timer_counter[9] ;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net79;
 wire net142;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net143;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net144;
 wire net130;
 wire net131;
 wire timeout_transmission;
 wire \timeout_value[0] ;
 wire \timeout_value[10] ;
 wire \timeout_value[11] ;
 wire \timeout_value[12] ;
 wire \timeout_value[13] ;
 wire \timeout_value[14] ;
 wire \timeout_value[15] ;
 wire \timeout_value[1] ;
 wire \timeout_value[2] ;
 wire \timeout_value[3] ;
 wire \timeout_value[4] ;
 wire \timeout_value[5] ;
 wire \timeout_value[6] ;
 wire \timeout_value[7] ;
 wire \timeout_value[8] ;
 wire \timeout_value[9] ;
 wire \io_i2c_scl_read_buffercc/_0_ ;
 wire \io_i2c_scl_read_buffercc/_1_ ;
 wire net77;
 wire \io_i2c_scl_read_buffercc/buffers_0 ;
 wire \io_i2c_sda_read_buffercc/_0_ ;
 wire \io_i2c_sda_read_buffercc/_1_ ;
 wire \io_i2c_sda_read_buffercc/buffers_0 ;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net76;
 wire net78;
 wire net188;
 wire clknet_4_1_0_clock;
 wire clknet_4_6_0_clock;
 wire net198;
 wire net189;
 wire net190;
 wire net192;
 wire net191;
 wire net193;
 wire net200;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net199;
 wire clknet_0_clock;
 wire clknet_4_0_0_clock;
 wire clknet_4_5_0_clock;
 wire net186;
 wire net185;
 wire clknet_4_3_0_clock;
 wire clknet_4_4_0_clock;
 wire net187;
 wire clknet_4_2_0_clock;
 wire clknet_4_7_0_clock;
 wire clknet_4_8_0_clock;
 wire clknet_4_9_0_clock;
 wire clknet_4_10_0_clock;
 wire clknet_4_11_0_clock;
 wire clknet_4_12_0_clock;
 wire clknet_4_13_0_clock;
 wire clknet_4_14_0_clock;
 wire clknet_4_15_0_clock;

 sg13g2_nor3_1 _366_ (.A(\ctrl_frameCounter[1] ),
    .B(\ctrl_frameCounter[3] ),
    .C(\ctrl_frameCounter[2] ),
    .Y(_076_));
 sg13g2_and2_1 _367_ (.A(\ctrl_frameCounter[0] ),
    .B(_076_),
    .X(net141));
 sg13g2_xor2_1 _369_ (.B(filter_sda_regNext),
    .A(filter_sda),
    .X(_078_));
 sg13g2_nand2_1 _370_ (.Y(_079_),
    .A(filter_scl),
    .B(_078_));
 sg13g2_xor2_1 _371_ (.B(\timeout_value[11] ),
    .A(net105),
    .X(_080_));
 sg13g2_xor2_1 _372_ (.B(\timeout_value[10] ),
    .A(net104),
    .X(_081_));
 sg13g2_xor2_1 _374_ (.B(\timeout_value[0] ),
    .A(net103),
    .X(_083_));
 sg13g2_xor2_1 _376_ (.B(\timeout_value[8] ),
    .A(net117),
    .X(_085_));
 sg13g2_nor4_1 _377_ (.A(_080_),
    .B(_081_),
    .C(_083_),
    .D(_085_),
    .Y(_086_));
 sg13g2_xor2_1 _378_ (.B(\timeout_value[3] ),
    .A(net112),
    .X(_087_));
 sg13g2_xor2_1 _380_ (.B(\timeout_value[5] ),
    .A(net114),
    .X(_089_));
 sg13g2_xor2_1 _382_ (.B(\timeout_value[7] ),
    .A(net116),
    .X(_091_));
 sg13g2_xor2_1 _384_ (.B(\timeout_value[6] ),
    .A(net115),
    .X(_093_));
 sg13g2_nor4_1 _385_ (.A(_087_),
    .B(_089_),
    .C(_091_),
    .D(_093_),
    .Y(_094_));
 sg13g2_xor2_1 _387_ (.B(\timeout_value[13] ),
    .A(net107),
    .X(_096_));
 sg13g2_xor2_1 _388_ (.B(\timeout_value[15] ),
    .A(net109),
    .X(_097_));
 sg13g2_xor2_1 _390_ (.B(\timeout_value[1] ),
    .A(net110),
    .X(_099_));
 sg13g2_xor2_1 _392_ (.B(\timeout_value[12] ),
    .A(net106),
    .X(_101_));
 sg13g2_nor4_1 _393_ (.A(_096_),
    .B(_097_),
    .C(_099_),
    .D(_101_),
    .Y(_102_));
 sg13g2_xor2_1 _395_ (.B(\timeout_value[4] ),
    .A(net113),
    .X(_104_));
 sg13g2_xor2_1 _396_ (.B(\timeout_value[2] ),
    .A(net111),
    .X(_105_));
 sg13g2_xor2_1 _398_ (.B(\timeout_value[9] ),
    .A(net118),
    .X(_107_));
 sg13g2_xor2_1 _399_ (.B(\timeout_value[14] ),
    .A(net108),
    .X(_108_));
 sg13g2_nor4_1 _400_ (.A(_104_),
    .B(_105_),
    .C(_107_),
    .D(_108_),
    .Y(_109_));
 sg13g2_nand4_1 _401_ (.B(_094_),
    .C(_102_),
    .A(_086_),
    .Y(_110_),
    .D(_109_));
 sg13g2_nand2_1 _403_ (.Y(_112_),
    .A(_079_),
    .B(_110_));
 sg13g2_nor2b_1 _405_ (.A(net79),
    .B_N(net142),
    .Y(_114_));
 sg13g2_nand2_1 _406_ (.Y(_115_),
    .A(net200),
    .B(_114_));
 sg13g2_inv_4 _407_ (.A(net131),
    .Y(_116_));
 sg13g2_nor4_1 _412_ (.A(\ctrl_bitCounter[4] ),
    .B(\_zz_ctrl_sdaWrite_1[1] ),
    .C(\_zz_ctrl_sdaWrite_1[0] ),
    .D(\_zz_ctrl_sdaWrite_1[2] ),
    .Y(_121_));
 sg13g2_nand2_1 _413_ (.Y(_122_),
    .A(\ctrl_bitCounter[3] ),
    .B(_121_));
 sg13g2_nor2_1 _414_ (.A(_116_),
    .B(_122_),
    .Y(_123_));
 sg13g2_nor2_1 _415_ (.A(net195),
    .B(net140),
    .Y(_124_));
 sg13g2_mux2_1 _416_ (.A0(net140),
    .A1(_124_),
    .S(_076_),
    .X(_125_));
 sg13g2_nor2_1 _417_ (.A(ctrl_cmdLock),
    .B(_125_),
    .Y(_126_));
 sg13g2_nand3_1 _418_ (.B(_123_),
    .C(_126_),
    .A(\ctrl_state[0] ),
    .Y(_127_));
 sg13g2_o21ai_1 _419_ (.B1(_127_),
    .Y(_009_),
    .A1(_112_),
    .A2(_115_));
 sg13g2_inv_1 _420_ (.Y(_128_),
    .A(net130));
 sg13g2_nand3_1 _421_ (.B(_128_),
    .C(\ctrl_state[1] ),
    .A(net200),
    .Y(_129_));
 sg13g2_nand3_1 _422_ (.B(net142),
    .C(net79),
    .A(net200),
    .Y(_130_));
 sg13g2_o21ai_1 _423_ (.B1(_130_),
    .Y(_008_),
    .A1(_112_),
    .A2(_129_));
 sg13g2_a22oi_1 _424_ (.Y(_131_),
    .B1(_078_),
    .B2(net194),
    .A2(\ctrl_state[1] ),
    .A1(net130));
 sg13g2_nor2_1 _425_ (.A(\ctrl_state[1] ),
    .B(_114_),
    .Y(_132_));
 sg13g2_a21oi_1 _426_ (.A1(_110_),
    .A2(_131_),
    .Y(_133_),
    .B1(_132_));
 sg13g2_nor3_1 _427_ (.A(ctrl_cmdLock),
    .B(_125_),
    .C(_122_),
    .Y(_134_));
 sg13g2_nand2b_1 _428_ (.Y(_135_),
    .B(\ctrl_state[0] ),
    .A_N(_134_));
 sg13g2_nand3b_1 _430_ (.B(_135_),
    .C(net200),
    .Y(_007_),
    .A_N(_133_));
 sg13g2_nand3b_1 _431_ (.B(filter_scl_regNext),
    .C(ctrl_transmission),
    .Y(_137_),
    .A_N(net194));
 sg13g2_nor3_1 _433_ (.A(\ctrl_state[0] ),
    .B(net142),
    .C(_128_),
    .Y(net144));
 sg13g2_a21o_1 _435_ (.A2(_137_),
    .A1(ctrl_cmdLock),
    .B1(net144),
    .X(_000_));
 sg13g2_inv_1 _436_ (.Y(_140_),
    .A(net129));
 sg13g2_nor2_1 _437_ (.A(ctrl_response_error),
    .B(net144),
    .Y(_141_));
 sg13g2_and2_1 _438_ (.A(_079_),
    .B(_110_),
    .X(_142_));
 sg13g2_a22oi_1 _440_ (.Y(_006_),
    .B1(_141_),
    .B2(_142_),
    .A2(net144),
    .A1(_140_));
 sg13g2_inv_1 _441_ (.Y(_144_),
    .A(filter_sda));
 sg13g2_and3_1 _442_ (.X(_145_),
    .A(\_zz_ctrl_sdaWrite_1[1] ),
    .B(net196),
    .C(\_zz_ctrl_sdaWrite_1[2] ));
 sg13g2_nor4_1 _443_ (.A(net195),
    .B(\ctrl_frameCounter[1] ),
    .C(\ctrl_frameCounter[3] ),
    .D(\ctrl_frameCounter[2] ),
    .Y(_146_));
 sg13g2_nand2_1 _444_ (.Y(_147_),
    .A(net194),
    .B(ctrl_transmission));
 sg13g2_nor4_1 _445_ (.A(filter_scl_regNext),
    .B(\ctrl_bitCounter[3] ),
    .C(\ctrl_bitCounter[4] ),
    .D(_147_),
    .Y(_148_));
 sg13g2_nand3_1 _447_ (.B(_146_),
    .C(_148_),
    .A(_145_),
    .Y(_150_));
 sg13g2_nand4_1 _448_ (.B(_079_),
    .C(_110_),
    .A(net140),
    .Y(_151_),
    .D(_150_));
 sg13g2_o21ai_1 _449_ (.B1(_151_),
    .Y(_005_),
    .A1(_144_),
    .A2(_150_));
 sg13g2_nor2b_1 _450_ (.A(net194),
    .B_N(filter_scl_regNext),
    .Y(_152_));
 sg13g2_nand4_1 _451_ (.B(ctrl_transmission),
    .C(_121_),
    .A(\ctrl_bitCounter[3] ),
    .Y(_153_),
    .D(_152_));
 sg13g2_nand4_1 _453_ (.B(_079_),
    .C(_110_),
    .A(net195),
    .Y(_155_),
    .D(_153_));
 sg13g2_o21ai_1 _454_ (.B1(_155_),
    .Y(_001_),
    .A1(net195),
    .A2(_153_));
 sg13g2_nand2_1 _455_ (.Y(_156_),
    .A(\ctrl_frameCounter[1] ),
    .B(_153_));
 sg13g2_nor2_1 _456_ (.A(net195),
    .B(_153_),
    .Y(_157_));
 sg13g2_nor2b_1 _457_ (.A(\ctrl_frameCounter[1] ),
    .B_N(net195),
    .Y(_158_));
 sg13g2_nor2_1 _458_ (.A(_122_),
    .B(_137_),
    .Y(_159_));
 sg13g2_a22oi_1 _459_ (.Y(_160_),
    .B1(_158_),
    .B2(_159_),
    .A2(_157_),
    .A1(\ctrl_frameCounter[1] ));
 sg13g2_o21ai_1 _460_ (.B1(_160_),
    .Y(_002_),
    .A1(_112_),
    .A2(_156_));
 sg13g2_nand2_1 _461_ (.Y(_161_),
    .A(\ctrl_frameCounter[2] ),
    .B(_153_));
 sg13g2_nand2_1 _462_ (.Y(_162_),
    .A(net195),
    .B(\ctrl_frameCounter[1] ));
 sg13g2_xnor2_1 _463_ (.Y(_163_),
    .A(\ctrl_frameCounter[2] ),
    .B(_162_));
 sg13g2_nand2_1 _464_ (.Y(_164_),
    .A(_159_),
    .B(_163_));
 sg13g2_o21ai_1 _465_ (.B1(_164_),
    .Y(_003_),
    .A1(_112_),
    .A2(_161_));
 sg13g2_nand2_1 _466_ (.Y(_165_),
    .A(\ctrl_frameCounter[3] ),
    .B(_153_));
 sg13g2_nand3_1 _467_ (.B(\ctrl_frameCounter[1] ),
    .C(\ctrl_frameCounter[2] ),
    .A(net195),
    .Y(_166_));
 sg13g2_nor2_1 _468_ (.A(\ctrl_frameCounter[3] ),
    .B(_166_),
    .Y(_167_));
 sg13g2_and2_1 _469_ (.A(\ctrl_frameCounter[3] ),
    .B(_166_),
    .X(_168_));
 sg13g2_o21ai_1 _470_ (.B1(_159_),
    .Y(_169_),
    .A1(_167_),
    .A2(_168_));
 sg13g2_o21ai_1 _471_ (.B1(_169_),
    .Y(_004_),
    .A1(_112_),
    .A2(_165_));
 sg13g2_and2_1 _472_ (.A(ctrl_transmission),
    .B(_152_),
    .X(_170_));
 sg13g2_nor2_1 _474_ (.A(net196),
    .B(_170_),
    .Y(_172_));
 sg13g2_a21o_1 _475_ (.A2(_170_),
    .A1(net196),
    .B1(_159_),
    .X(_173_));
 sg13g2_a21oi_1 _476_ (.A1(_142_),
    .A2(_172_),
    .Y(_014_),
    .B1(_173_));
 sg13g2_nor2_1 _477_ (.A(\_zz_ctrl_sdaWrite_1[1] ),
    .B(_170_),
    .Y(_174_));
 sg13g2_or2_1 _478_ (.X(_175_),
    .B(net196),
    .A(\_zz_ctrl_sdaWrite_1[1] ));
 sg13g2_nand2_1 _479_ (.Y(_176_),
    .A(\_zz_ctrl_sdaWrite_1[1] ),
    .B(net196));
 sg13g2_a21oi_1 _480_ (.A1(_175_),
    .A2(_176_),
    .Y(_177_),
    .B1(_137_));
 sg13g2_a21oi_1 _481_ (.A1(_142_),
    .A2(_174_),
    .Y(_015_),
    .B1(_177_));
 sg13g2_nor2_1 _482_ (.A(\_zz_ctrl_sdaWrite_1[2] ),
    .B(_170_),
    .Y(_178_));
 sg13g2_xor2_1 _483_ (.B(_176_),
    .A(\_zz_ctrl_sdaWrite_1[2] ),
    .X(_179_));
 sg13g2_a22oi_1 _484_ (.Y(_016_),
    .B1(_179_),
    .B2(_170_),
    .A2(_178_),
    .A1(_142_));
 sg13g2_nand2_1 _485_ (.Y(_180_),
    .A(_170_),
    .B(_145_));
 sg13g2_nand3_1 _486_ (.B(net196),
    .C(\_zz_ctrl_sdaWrite_1[2] ),
    .A(\_zz_ctrl_sdaWrite_1[1] ),
    .Y(_181_));
 sg13g2_a21oi_1 _487_ (.A1(_122_),
    .A2(_181_),
    .Y(_182_),
    .B1(_137_));
 sg13g2_mux2_1 _488_ (.A0(_180_),
    .A1(_182_),
    .S(\ctrl_bitCounter[3] ),
    .X(_183_));
 sg13g2_o21ai_1 _489_ (.B1(_183_),
    .Y(_017_),
    .A1(_142_),
    .A2(_170_));
 sg13g2_nor2_1 _490_ (.A(_137_),
    .B(_181_),
    .Y(_184_));
 sg13g2_nand3_1 _491_ (.B(\ctrl_bitCounter[4] ),
    .C(_184_),
    .A(\ctrl_bitCounter[3] ),
    .Y(_185_));
 sg13g2_a221oi_1 _492_ (.B2(\ctrl_bitCounter[3] ),
    .C1(\ctrl_bitCounter[4] ),
    .B1(_184_),
    .A1(net194),
    .Y(_186_),
    .A2(_078_));
 sg13g2_o21ai_1 _493_ (.B1(_186_),
    .Y(_187_),
    .A1(_110_),
    .A2(_170_));
 sg13g2_and2_1 _494_ (.A(_185_),
    .B(_187_),
    .X(_018_));
 sg13g2_mux2_1 _495_ (.A0(\_zz_ctrl_sdaWrite[7] ),
    .A1(net121),
    .S(net192),
    .X(_019_));
 sg13g2_mux2_1 _496_ (.A0(\_zz_ctrl_sdaWrite[6] ),
    .A1(net122),
    .S(net192),
    .X(_020_));
 sg13g2_mux2_1 _497_ (.A0(\_zz_ctrl_sdaWrite[5] ),
    .A1(net123),
    .S(net192),
    .X(_021_));
 sg13g2_mux2_1 _498_ (.A0(\_zz_ctrl_sdaWrite[4] ),
    .A1(net124),
    .S(net192),
    .X(_022_));
 sg13g2_mux2_1 _499_ (.A0(\_zz_ctrl_sdaWrite[3] ),
    .A1(net125),
    .S(net192),
    .X(_023_));
 sg13g2_mux2_1 _500_ (.A0(\_zz_ctrl_sdaWrite[2] ),
    .A1(net126),
    .S(net192),
    .X(_024_));
 sg13g2_mux2_1 _501_ (.A0(\_zz_ctrl_sdaWrite[1] ),
    .A1(net127),
    .S(net192),
    .X(_025_));
 sg13g2_mux2_1 _502_ (.A0(\_zz_ctrl_sdaWrite[0] ),
    .A1(net128),
    .S(net192),
    .X(_026_));
 sg13g2_mux2_1 _503_ (.A0(net132),
    .A1(filter_sda),
    .S(net191),
    .X(_028_));
 sg13g2_mux2_1 _504_ (.A0(net133),
    .A1(net132),
    .S(net191),
    .X(_029_));
 sg13g2_mux2_1 _505_ (.A0(net134),
    .A1(net133),
    .S(net191),
    .X(_030_));
 sg13g2_mux2_1 _506_ (.A0(net135),
    .A1(net134),
    .S(net191),
    .X(_031_));
 sg13g2_mux2_1 _507_ (.A0(net136),
    .A1(net135),
    .S(net191),
    .X(_032_));
 sg13g2_mux2_1 _508_ (.A0(net137),
    .A1(net136),
    .S(net191),
    .X(_033_));
 sg13g2_mux2_1 _509_ (.A0(net138),
    .A1(net137),
    .S(net191),
    .X(_034_));
 sg13g2_mux2_1 _510_ (.A0(net139),
    .A1(net138),
    .S(net191),
    .X(_035_));
 sg13g2_inv_1 _511_ (.Y(_188_),
    .A(filter_scl));
 sg13g2_o21ai_1 _512_ (.B1(timeout_transmission),
    .Y(_189_),
    .A1(filter_sda_regNext),
    .A2(_188_));
 sg13g2_inv_1 _513_ (.Y(_190_),
    .A(timeout_transmission));
 sg13g2_nand2_1 _514_ (.Y(_191_),
    .A(filter_sda_regNext),
    .B(filter_scl));
 sg13g2_a21o_1 _515_ (.A2(_191_),
    .A1(_190_),
    .B1(filter_sda),
    .X(_192_));
 sg13g2_a21oi_1 _517_ (.A1(_189_),
    .A2(_192_),
    .Y(_057_),
    .B1(_116_));
 sg13g2_nor4_2 _518_ (.A(\filter_timer_counter[0] ),
    .B(\filter_timer_counter[1] ),
    .C(\filter_timer_counter[2] ),
    .Y(_194_),
    .D(\filter_timer_counter[3] ));
 sg13g2_nor4_2 _519_ (.A(\filter_timer_counter[4] ),
    .B(\filter_timer_counter[5] ),
    .C(\filter_timer_counter[6] ),
    .Y(_195_),
    .D(\filter_timer_counter[7] ));
 sg13g2_nor2_1 _520_ (.A(\filter_timer_counter[9] ),
    .B(\filter_timer_counter[8] ),
    .Y(_196_));
 sg13g2_and3_1 _521_ (.X(_197_),
    .A(_194_),
    .B(_195_),
    .C(_196_));
 sg13g2_or3_1 _524_ (.A(\filter_timer_counter[13] ),
    .B(\filter_timer_counter[15] ),
    .C(\filter_timer_counter[14] ),
    .X(_200_));
 sg13g2_or2_2 _525_ (.X(_201_),
    .B(\filter_timer_counter[10] ),
    .A(\filter_timer_counter[11] ));
 sg13g2_nor3_2 _526_ (.A(\filter_timer_counter[12] ),
    .B(_200_),
    .C(_201_),
    .Y(_202_));
 sg13g2_nand2_1 _527_ (.Y(_203_),
    .A(_197_),
    .B(_202_));
 sg13g2_nand2_1 _529_ (.Y(_205_),
    .A(_zz_filter_sampler_sclSamples_1),
    .B(_203_));
 sg13g2_nand3_1 _530_ (.B(_195_),
    .C(_196_),
    .A(_194_),
    .Y(_206_));
 sg13g2_or3_2 _532_ (.A(\filter_timer_counter[12] ),
    .B(_200_),
    .C(_201_),
    .X(_208_));
 sg13g2_nor2_2 _533_ (.A(_206_),
    .B(_208_),
    .Y(_209_));
 sg13g2_nand2_1 _534_ (.Y(_210_),
    .A(_zz_filter_sampler_sclSamples_0),
    .B(net188));
 sg13g2_nand3_1 _535_ (.B(_205_),
    .C(_210_),
    .A(net199),
    .Y(_010_));
 sg13g2_nand2_1 _536_ (.Y(_211_),
    .A(_zz_filter_sampler_sclSamples_2),
    .B(_203_));
 sg13g2_nand2_1 _537_ (.Y(_212_),
    .A(_zz_filter_sampler_sclSamples_1),
    .B(net188));
 sg13g2_nand3_1 _538_ (.B(_211_),
    .C(_212_),
    .A(net199),
    .Y(_011_));
 sg13g2_nand2_1 _539_ (.Y(_213_),
    .A(_zz_filter_sampler_sdaSamples_1),
    .B(_203_));
 sg13g2_nand2_1 _540_ (.Y(_214_),
    .A(_zz_filter_sampler_sdaSamples_0),
    .B(_209_));
 sg13g2_nand3_1 _541_ (.B(_213_),
    .C(_214_),
    .A(net199),
    .Y(_012_));
 sg13g2_nand2_1 _542_ (.Y(_215_),
    .A(_zz_filter_sampler_sdaSamples_2),
    .B(_203_));
 sg13g2_nand2_1 _543_ (.Y(_216_),
    .A(_zz_filter_sampler_sdaSamples_1),
    .B(_209_));
 sg13g2_nand3_1 _544_ (.B(_215_),
    .C(_216_),
    .A(net199),
    .Y(_013_));
 sg13g2_nand2_1 _545_ (.Y(_217_),
    .A(net131),
    .B(net140));
 sg13g2_or4_1 _546_ (.A(\ctrl_bitCounter[3] ),
    .B(\ctrl_bitCounter[4] ),
    .C(_146_),
    .D(_217_),
    .X(_218_));
 sg13g2_mux4_1 _547_ (.S0(net196),
    .A0(\_zz_ctrl_sdaWrite[0] ),
    .A1(\_zz_ctrl_sdaWrite[1] ),
    .A2(\_zz_ctrl_sdaWrite[2] ),
    .A3(\_zz_ctrl_sdaWrite[3] ),
    .S1(\_zz_ctrl_sdaWrite_1[1] ),
    .X(_219_));
 sg13g2_mux4_1 _548_ (.S0(net196),
    .A0(\_zz_ctrl_sdaWrite[4] ),
    .A1(\_zz_ctrl_sdaWrite[5] ),
    .A2(\_zz_ctrl_sdaWrite[6] ),
    .A3(\_zz_ctrl_sdaWrite[7] ),
    .S1(\_zz_ctrl_sdaWrite_1[1] ),
    .X(_220_));
 sg13g2_mux2_1 _549_ (.A0(_219_),
    .A1(_220_),
    .S(\_zz_ctrl_sdaWrite_1[2] ),
    .X(_221_));
 sg13g2_xnor2_1 _550_ (.Y(_222_),
    .A(net96),
    .B(net133));
 sg13g2_xnor2_1 _551_ (.Y(_223_),
    .A(net97),
    .B(net134));
 sg13g2_xnor2_1 _552_ (.Y(_224_),
    .A(net102),
    .B(net139));
 sg13g2_nand3_1 _553_ (.B(_223_),
    .C(_224_),
    .A(_222_),
    .Y(_225_));
 sg13g2_xor2_1 _554_ (.B(net136),
    .A(net99),
    .X(_226_));
 sg13g2_xor2_1 _555_ (.B(net137),
    .A(net100),
    .X(_227_));
 sg13g2_xnor2_1 _556_ (.Y(_228_),
    .A(net101),
    .B(net138));
 sg13g2_xnor2_1 _557_ (.Y(_229_),
    .A(net98),
    .B(net135));
 sg13g2_nand3_1 _558_ (.B(_228_),
    .C(_229_),
    .A(_146_),
    .Y(_230_));
 sg13g2_nor4_1 _559_ (.A(_225_),
    .B(_226_),
    .C(_227_),
    .D(_230_),
    .Y(_231_));
 sg13g2_nor3_1 _560_ (.A(net140),
    .B(ctrl_response_error),
    .C(_146_),
    .Y(_232_));
 sg13g2_o21ai_1 _561_ (.B1(_123_),
    .Y(_233_),
    .A1(_231_),
    .A2(_232_));
 sg13g2_o21ai_1 _562_ (.B1(_233_),
    .Y(_027_),
    .A1(_218_),
    .A2(_221_));
 sg13g2_nand2_1 _563_ (.Y(_040_),
    .A(_144_),
    .B(net200));
 sg13g2_nand4_1 _564_ (.B(ctrl_transmission),
    .C(_079_),
    .A(net200),
    .Y(_234_),
    .D(_110_));
 sg13g2_o21ai_1 _565_ (.B1(_234_),
    .Y(_036_),
    .A1(_191_),
    .A2(_040_));
 sg13g2_nor3_1 _566_ (.A(_zz_filter_sampler_sclSamples_2),
    .B(_zz_filter_sampler_sclSamples_1),
    .C(_zz_filter_sampler_sclSamples_0),
    .Y(_235_));
 sg13g2_mux2_1 _567_ (.A0(_188_),
    .A1(_235_),
    .S(_209_),
    .X(_236_));
 sg13g2_and2_1 _568_ (.A(_zz_filter_sampler_sclSamples_1),
    .B(_zz_filter_sampler_sclSamples_0),
    .X(_237_));
 sg13g2_a21oi_1 _569_ (.A1(_zz_filter_sampler_sclSamples_2),
    .A2(_237_),
    .Y(_238_),
    .B1(filter_scl));
 sg13g2_o21ai_1 _570_ (.B1(net199),
    .Y(_037_),
    .A1(_236_),
    .A2(_238_));
 sg13g2_nand2_1 _571_ (.Y(_038_),
    .A(_188_),
    .B(net199));
 sg13g2_nor3_1 _572_ (.A(_zz_filter_sampler_sdaSamples_2),
    .B(_zz_filter_sampler_sdaSamples_1),
    .C(_zz_filter_sampler_sdaSamples_0),
    .Y(_239_));
 sg13g2_mux2_1 _573_ (.A0(_144_),
    .A1(_239_),
    .S(_209_),
    .X(_240_));
 sg13g2_and2_1 _574_ (.A(_zz_filter_sampler_sdaSamples_1),
    .B(_zz_filter_sampler_sdaSamples_0),
    .X(_241_));
 sg13g2_a21oi_1 _575_ (.A1(_zz_filter_sampler_sdaSamples_2),
    .A2(_241_),
    .Y(_242_),
    .B1(filter_sda));
 sg13g2_o21ai_1 _576_ (.B1(net199),
    .Y(_039_),
    .A1(_240_),
    .A2(_242_));
 sg13g2_nor2_1 _577_ (.A(net80),
    .B(net189),
    .Y(_243_));
 sg13g2_nor3_1 _578_ (.A(\filter_timer_counter[0] ),
    .B(net198),
    .C(_243_),
    .Y(_041_));
 sg13g2_xnor2_1 _579_ (.Y(_244_),
    .A(\filter_timer_counter[10] ),
    .B(_206_));
 sg13g2_o21ai_1 _580_ (.B1(_244_),
    .Y(_245_),
    .A1(net81),
    .A2(_203_));
 sg13g2_nor2_1 _581_ (.A(net198),
    .B(_245_),
    .Y(_042_));
 sg13g2_nor2_1 _582_ (.A(\filter_timer_counter[11] ),
    .B(\filter_timer_counter[10] ),
    .Y(_246_));
 sg13g2_nand4_1 _583_ (.B(_195_),
    .C(_196_),
    .A(_194_),
    .Y(_247_),
    .D(_246_));
 sg13g2_o21ai_1 _585_ (.B1(\filter_timer_counter[11] ),
    .Y(_249_),
    .A1(\filter_timer_counter[10] ),
    .A2(_206_));
 sg13g2_o21ai_1 _586_ (.B1(net131),
    .Y(_250_),
    .A1(net82),
    .A2(net189));
 sg13g2_a21oi_1 _587_ (.A1(_247_),
    .A2(_249_),
    .Y(_043_),
    .B1(_250_));
 sg13g2_nor2_1 _588_ (.A(net83),
    .B(_200_),
    .Y(_251_));
 sg13g2_nor3_1 _589_ (.A(net193),
    .B(_247_),
    .C(_251_),
    .Y(_252_));
 sg13g2_a21oi_1 _590_ (.A1(net193),
    .A2(_247_),
    .Y(_253_),
    .B1(_252_));
 sg13g2_nor2_1 _591_ (.A(net197),
    .B(_253_),
    .Y(_044_));
 sg13g2_o21ai_1 _592_ (.B1(\filter_timer_counter[13] ),
    .Y(_254_),
    .A1(net193),
    .A2(_247_));
 sg13g2_nor3_1 _593_ (.A(\filter_timer_counter[15] ),
    .B(\filter_timer_counter[14] ),
    .C(net84),
    .Y(_255_));
 sg13g2_or4_1 _594_ (.A(\filter_timer_counter[13] ),
    .B(net193),
    .C(_247_),
    .D(_255_),
    .X(_256_));
 sg13g2_a21oi_1 _595_ (.A1(_254_),
    .A2(_256_),
    .Y(_045_),
    .B1(net197));
 sg13g2_inv_1 _596_ (.Y(_257_),
    .A(\filter_timer_counter[14] ));
 sg13g2_o21ai_1 _597_ (.B1(_257_),
    .Y(_258_),
    .A1(\filter_timer_counter[15] ),
    .A2(net85));
 sg13g2_nor3_1 _598_ (.A(\filter_timer_counter[13] ),
    .B(net193),
    .C(_247_),
    .Y(_259_));
 sg13g2_mux2_1 _599_ (.A0(_257_),
    .A1(_258_),
    .S(_259_),
    .X(_260_));
 sg13g2_nor2_1 _600_ (.A(net197),
    .B(_260_),
    .Y(_046_));
 sg13g2_nor4_2 _601_ (.A(\filter_timer_counter[13] ),
    .B(net193),
    .C(\filter_timer_counter[14] ),
    .Y(_261_),
    .D(_247_));
 sg13g2_nand3b_1 _602_ (.B(net86),
    .C(_261_),
    .Y(_262_),
    .A_N(\filter_timer_counter[15] ));
 sg13g2_nand2b_1 _603_ (.Y(_263_),
    .B(\filter_timer_counter[15] ),
    .A_N(_261_));
 sg13g2_a21oi_1 _604_ (.A1(_262_),
    .A2(_263_),
    .Y(_047_),
    .B1(net197));
 sg13g2_nor2_1 _605_ (.A(net87),
    .B(net189),
    .Y(_264_));
 sg13g2_xor2_1 _606_ (.B(\filter_timer_counter[1] ),
    .A(\filter_timer_counter[0] ),
    .X(_265_));
 sg13g2_nor3_1 _607_ (.A(net198),
    .B(_264_),
    .C(_265_),
    .Y(_048_));
 sg13g2_nor2_1 _608_ (.A(net88),
    .B(net189),
    .Y(_266_));
 sg13g2_nor2_1 _609_ (.A(\filter_timer_counter[0] ),
    .B(\filter_timer_counter[1] ),
    .Y(_267_));
 sg13g2_xnor2_1 _610_ (.Y(_268_),
    .A(\filter_timer_counter[2] ),
    .B(_267_));
 sg13g2_nor3_1 _611_ (.A(net198),
    .B(_266_),
    .C(_268_),
    .Y(_049_));
 sg13g2_nor2_1 _612_ (.A(net89),
    .B(net189),
    .Y(_269_));
 sg13g2_nor3_1 _613_ (.A(\filter_timer_counter[0] ),
    .B(\filter_timer_counter[1] ),
    .C(\filter_timer_counter[2] ),
    .Y(_270_));
 sg13g2_xnor2_1 _614_ (.Y(_271_),
    .A(\filter_timer_counter[3] ),
    .B(_270_));
 sg13g2_nor3_1 _615_ (.A(net198),
    .B(_269_),
    .C(_271_),
    .Y(_050_));
 sg13g2_inv_1 _616_ (.Y(_272_),
    .A(net90));
 sg13g2_nand2b_1 _617_ (.Y(_273_),
    .B(\filter_timer_counter[4] ),
    .A_N(_194_));
 sg13g2_nand2b_1 _618_ (.Y(_274_),
    .B(_194_),
    .A_N(\filter_timer_counter[4] ));
 sg13g2_a221oi_1 _619_ (.B2(_274_),
    .C1(net197),
    .B1(_273_),
    .A1(_272_),
    .Y(_051_),
    .A2(net188));
 sg13g2_inv_1 _620_ (.Y(_275_),
    .A(net91));
 sg13g2_nand2_1 _621_ (.Y(_276_),
    .A(\filter_timer_counter[5] ),
    .B(_274_));
 sg13g2_or2_1 _622_ (.X(_277_),
    .B(_274_),
    .A(\filter_timer_counter[5] ));
 sg13g2_a221oi_1 _623_ (.B2(_277_),
    .C1(net197),
    .B1(_276_),
    .A1(_275_),
    .Y(_052_),
    .A2(net188));
 sg13g2_nor2_1 _624_ (.A(net92),
    .B(net189),
    .Y(_278_));
 sg13g2_xor2_1 _625_ (.B(_277_),
    .A(\filter_timer_counter[6] ),
    .X(_279_));
 sg13g2_nor3_1 _626_ (.A(net197),
    .B(_278_),
    .C(_279_),
    .Y(_053_));
 sg13g2_inv_1 _627_ (.Y(_280_),
    .A(net93));
 sg13g2_o21ai_1 _628_ (.B1(\filter_timer_counter[7] ),
    .Y(_281_),
    .A1(\filter_timer_counter[6] ),
    .A2(_277_));
 sg13g2_nand2_1 _629_ (.Y(_282_),
    .A(_194_),
    .B(_195_));
 sg13g2_a221oi_1 _630_ (.B2(_282_),
    .C1(net197),
    .B1(_281_),
    .A1(_280_),
    .Y(_054_),
    .A2(net188));
 sg13g2_xnor2_1 _631_ (.Y(_283_),
    .A(\filter_timer_counter[8] ),
    .B(_282_));
 sg13g2_o21ai_1 _632_ (.B1(_283_),
    .Y(_284_),
    .A1(net94),
    .A2(net189));
 sg13g2_nor2_1 _633_ (.A(net198),
    .B(_284_),
    .Y(_055_));
 sg13g2_o21ai_1 _634_ (.B1(\filter_timer_counter[9] ),
    .Y(_285_),
    .A1(\filter_timer_counter[8] ),
    .A2(_282_));
 sg13g2_o21ai_1 _635_ (.B1(net131),
    .Y(_286_),
    .A1(net95),
    .A2(net189));
 sg13g2_a21oi_1 _636_ (.A1(_206_),
    .A2(_285_),
    .Y(_056_),
    .B1(_286_));
 sg13g2_nor2_1 _637_ (.A(_190_),
    .B(_116_),
    .Y(_287_));
 sg13g2_nand3_1 _638_ (.B(_202_),
    .C(_287_),
    .A(_197_),
    .Y(_288_));
 sg13g2_nand2b_1 _640_ (.Y(_290_),
    .B(filter_sda_regNext),
    .A_N(filter_sda));
 sg13g2_nand3_1 _641_ (.B(filter_scl_regNext),
    .C(_290_),
    .A(filter_scl),
    .Y(_291_));
 sg13g2_or2_1 _642_ (.X(_292_),
    .B(filter_scl_regNext),
    .A(filter_scl));
 sg13g2_nor4_1 _643_ (.A(\filter_timer_counter[12] ),
    .B(_190_),
    .C(_200_),
    .D(_201_),
    .Y(_293_));
 sg13g2_a221oi_1 _644_ (.B2(_197_),
    .C1(_116_),
    .B1(_293_),
    .A1(_291_),
    .Y(_294_),
    .A2(_292_));
 sg13g2_nand2_1 _647_ (.Y(_297_),
    .A(\timeout_value[0] ),
    .B(net185));
 sg13g2_o21ai_1 _648_ (.B1(_297_),
    .Y(_058_),
    .A1(\timeout_value[0] ),
    .A2(net187));
 sg13g2_nand4_1 _649_ (.B(\timeout_value[1] ),
    .C(\timeout_value[2] ),
    .A(\timeout_value[0] ),
    .Y(_298_),
    .D(\timeout_value[3] ));
 sg13g2_nand3_1 _651_ (.B(\timeout_value[5] ),
    .C(\timeout_value[6] ),
    .A(\timeout_value[4] ),
    .Y(_300_));
 sg13g2_or2_2 _652_ (.X(_301_),
    .B(_300_),
    .A(_298_));
 sg13g2_nand3_1 _654_ (.B(\timeout_value[8] ),
    .C(\timeout_value[9] ),
    .A(\timeout_value[7] ),
    .Y(_303_));
 sg13g2_o21ai_1 _655_ (.B1(\timeout_value[10] ),
    .Y(_304_),
    .A1(net190),
    .A2(_303_));
 sg13g2_or3_1 _656_ (.A(\timeout_value[10] ),
    .B(net190),
    .C(_303_),
    .X(_305_));
 sg13g2_a21oi_2 _657_ (.B1(net187),
    .Y(_306_),
    .A2(_305_),
    .A1(_304_));
 sg13g2_a21o_1 _658_ (.A2(net185),
    .A1(\timeout_value[10] ),
    .B1(_306_),
    .X(_059_));
 sg13g2_nand4_1 _659_ (.B(\timeout_value[8] ),
    .C(\timeout_value[9] ),
    .A(\timeout_value[7] ),
    .Y(_307_),
    .D(\timeout_value[10] ));
 sg13g2_o21ai_1 _660_ (.B1(\timeout_value[11] ),
    .Y(_308_),
    .A1(net190),
    .A2(_307_));
 sg13g2_or3_1 _661_ (.A(\timeout_value[11] ),
    .B(_301_),
    .C(_307_),
    .X(_309_));
 sg13g2_a21oi_2 _662_ (.B1(net187),
    .Y(_310_),
    .A2(_309_),
    .A1(_308_));
 sg13g2_a21o_1 _663_ (.A2(net186),
    .A1(\timeout_value[11] ),
    .B1(_310_),
    .X(_060_));
 sg13g2_nand2_1 _664_ (.Y(_311_),
    .A(\timeout_value[4] ),
    .B(\timeout_value[5] ));
 sg13g2_nand2_1 _665_ (.Y(_312_),
    .A(\timeout_value[6] ),
    .B(\timeout_value[11] ));
 sg13g2_nor4_2 _666_ (.A(_298_),
    .B(_311_),
    .C(_307_),
    .Y(_313_),
    .D(_312_));
 sg13g2_nand2b_1 _667_ (.Y(_314_),
    .B(\timeout_value[12] ),
    .A_N(_313_));
 sg13g2_nand2b_1 _668_ (.Y(_315_),
    .B(_313_),
    .A_N(\timeout_value[12] ));
 sg13g2_a21oi_2 _669_ (.B1(_288_),
    .Y(_316_),
    .A2(_315_),
    .A1(_314_));
 sg13g2_a21o_1 _670_ (.A2(_294_),
    .A1(\timeout_value[12] ),
    .B1(_316_),
    .X(_061_));
 sg13g2_nand2_1 _671_ (.Y(_317_),
    .A(\timeout_value[13] ),
    .B(_294_));
 sg13g2_nor4_2 _672_ (.A(_190_),
    .B(_116_),
    .C(_206_),
    .Y(_318_),
    .D(_208_));
 sg13g2_nand2_1 _673_ (.Y(_319_),
    .A(\timeout_value[12] ),
    .B(_313_));
 sg13g2_nand3_1 _674_ (.B(_318_),
    .C(_319_),
    .A(\timeout_value[13] ),
    .Y(_320_));
 sg13g2_or3_1 _675_ (.A(\timeout_value[13] ),
    .B(_288_),
    .C(_319_),
    .X(_321_));
 sg13g2_nand3_1 _676_ (.B(_320_),
    .C(_321_),
    .A(_317_),
    .Y(_062_));
 sg13g2_nand2_1 _677_ (.Y(_322_),
    .A(\timeout_value[14] ),
    .B(_294_));
 sg13g2_nand3_1 _678_ (.B(\timeout_value[13] ),
    .C(_313_),
    .A(\timeout_value[12] ),
    .Y(_323_));
 sg13g2_nand3_1 _679_ (.B(_318_),
    .C(_323_),
    .A(\timeout_value[14] ),
    .Y(_324_));
 sg13g2_inv_1 _680_ (.Y(_325_),
    .A(\timeout_value[14] ));
 sg13g2_nand3b_1 _681_ (.B(_325_),
    .C(_318_),
    .Y(_326_),
    .A_N(_323_));
 sg13g2_nand3_1 _682_ (.B(_324_),
    .C(_326_),
    .A(_322_),
    .Y(_063_));
 sg13g2_nand2_1 _683_ (.Y(_327_),
    .A(\timeout_value[15] ),
    .B(_294_));
 sg13g2_nand4_1 _684_ (.B(\timeout_value[13] ),
    .C(\timeout_value[14] ),
    .A(\timeout_value[12] ),
    .Y(_328_),
    .D(_313_));
 sg13g2_nand3_1 _685_ (.B(_318_),
    .C(_328_),
    .A(\timeout_value[15] ),
    .Y(_329_));
 sg13g2_or4_1 _686_ (.A(_325_),
    .B(\timeout_value[15] ),
    .C(_288_),
    .D(_323_),
    .X(_330_));
 sg13g2_nand3_1 _687_ (.B(_329_),
    .C(_330_),
    .A(_327_),
    .Y(_064_));
 sg13g2_nand2b_1 _688_ (.Y(_331_),
    .B(\timeout_value[1] ),
    .A_N(\timeout_value[0] ));
 sg13g2_nand2b_1 _689_ (.Y(_332_),
    .B(\timeout_value[0] ),
    .A_N(\timeout_value[1] ));
 sg13g2_a21oi_2 _690_ (.B1(net187),
    .Y(_333_),
    .A2(_332_),
    .A1(_331_));
 sg13g2_a21o_1 _691_ (.A2(net185),
    .A1(\timeout_value[1] ),
    .B1(_333_),
    .X(_065_));
 sg13g2_nand2_1 _692_ (.Y(_334_),
    .A(\timeout_value[0] ),
    .B(\timeout_value[1] ));
 sg13g2_xor2_1 _693_ (.B(_334_),
    .A(\timeout_value[2] ),
    .X(_335_));
 sg13g2_nand2_1 _694_ (.Y(_336_),
    .A(\timeout_value[2] ),
    .B(net185));
 sg13g2_o21ai_1 _695_ (.B1(_336_),
    .Y(_066_),
    .A1(net187),
    .A2(_335_));
 sg13g2_nand3_1 _696_ (.B(\timeout_value[1] ),
    .C(\timeout_value[2] ),
    .A(\timeout_value[0] ),
    .Y(_337_));
 sg13g2_xor2_1 _697_ (.B(_337_),
    .A(\timeout_value[3] ),
    .X(_338_));
 sg13g2_nand2_1 _698_ (.Y(_339_),
    .A(\timeout_value[3] ),
    .B(net185));
 sg13g2_o21ai_1 _699_ (.B1(_339_),
    .Y(_067_),
    .A1(net187),
    .A2(_338_));
 sg13g2_nand2_1 _700_ (.Y(_340_),
    .A(\timeout_value[4] ),
    .B(_298_));
 sg13g2_inv_1 _701_ (.Y(_341_),
    .A(\timeout_value[4] ));
 sg13g2_nand2b_1 _702_ (.Y(_342_),
    .B(_341_),
    .A_N(_298_));
 sg13g2_a21oi_2 _703_ (.B1(_288_),
    .Y(_343_),
    .A2(_342_),
    .A1(_340_));
 sg13g2_a21o_1 _704_ (.A2(net186),
    .A1(\timeout_value[4] ),
    .B1(_343_),
    .X(_068_));
 sg13g2_o21ai_1 _705_ (.B1(\timeout_value[5] ),
    .Y(_344_),
    .A1(_341_),
    .A2(_298_));
 sg13g2_or3_1 _706_ (.A(_341_),
    .B(\timeout_value[5] ),
    .C(_298_),
    .X(_345_));
 sg13g2_a21oi_2 _707_ (.B1(_288_),
    .Y(_346_),
    .A2(_345_),
    .A1(_344_));
 sg13g2_a21o_1 _708_ (.A2(net186),
    .A1(\timeout_value[5] ),
    .B1(_346_),
    .X(_069_));
 sg13g2_o21ai_1 _709_ (.B1(\timeout_value[6] ),
    .Y(_347_),
    .A1(_298_),
    .A2(_311_));
 sg13g2_or3_1 _710_ (.A(\timeout_value[6] ),
    .B(_298_),
    .C(_311_),
    .X(_348_));
 sg13g2_a21oi_2 _711_ (.B1(_288_),
    .Y(_349_),
    .A2(_348_),
    .A1(_347_));
 sg13g2_a21o_1 _712_ (.A2(net186),
    .A1(\timeout_value[6] ),
    .B1(_349_),
    .X(_070_));
 sg13g2_nand2_1 _713_ (.Y(_350_),
    .A(\timeout_value[7] ),
    .B(net186));
 sg13g2_nand3_1 _714_ (.B(_318_),
    .C(net190),
    .A(\timeout_value[7] ),
    .Y(_351_));
 sg13g2_inv_1 _715_ (.Y(_352_),
    .A(\timeout_value[7] ));
 sg13g2_nand3b_1 _716_ (.B(_352_),
    .C(_318_),
    .Y(_353_),
    .A_N(net190));
 sg13g2_nand3_1 _717_ (.B(_351_),
    .C(_353_),
    .A(_350_),
    .Y(_071_));
 sg13g2_nand3_1 _718_ (.B(_202_),
    .C(_287_),
    .A(_197_),
    .Y(_354_));
 sg13g2_nor2_1 _719_ (.A(_352_),
    .B(net190),
    .Y(_355_));
 sg13g2_xnor2_1 _720_ (.Y(_356_),
    .A(\timeout_value[8] ),
    .B(_355_));
 sg13g2_nand2_1 _721_ (.Y(_357_),
    .A(\timeout_value[8] ),
    .B(net186));
 sg13g2_o21ai_1 _722_ (.B1(_357_),
    .Y(_072_),
    .A1(_354_),
    .A2(_356_));
 sg13g2_nand2_1 _723_ (.Y(_358_),
    .A(\timeout_value[7] ),
    .B(\timeout_value[8] ));
 sg13g2_o21ai_1 _724_ (.B1(\timeout_value[9] ),
    .Y(_359_),
    .A1(net190),
    .A2(_358_));
 sg13g2_or3_1 _725_ (.A(\timeout_value[9] ),
    .B(net190),
    .C(_358_),
    .X(_360_));
 sg13g2_a21oi_1 _726_ (.A1(_359_),
    .A2(_360_),
    .Y(_361_),
    .B1(net187));
 sg13g2_a21o_1 _727_ (.A2(net185),
    .A1(\timeout_value[9] ),
    .B1(_361_),
    .X(_073_));
 sg13g2_tielo _731__1 (.L_LO(io_i2c_scl_write));
 sg13g2_dfrbpq_1 \_zz_filter_sampler_sclSamples_1$_SDFFE_PN1P_  (.RESET_B(net1),
    .D(_010_),
    .Q(_zz_filter_sampler_sclSamples_1),
    .CLK(clknet_4_9_0_clock));
 sg13g2_tiehi \_zz_filter_sampler_sclSamples_1$_SDFFE_PN1P__2  (.L_HI(net1));
 sg13g2_dfrbpq_1 \_zz_filter_sampler_sclSamples_2$_SDFFE_PN1P_  (.RESET_B(net2),
    .D(_011_),
    .Q(_zz_filter_sampler_sclSamples_2),
    .CLK(clknet_4_8_0_clock));
 sg13g2_tiehi \_zz_filter_sampler_sclSamples_2$_SDFFE_PN1P__3  (.L_HI(net2));
 sg13g2_dfrbpq_1 \_zz_filter_sampler_sdaSamples_1$_SDFFE_PN1P_  (.RESET_B(net3),
    .D(_012_),
    .Q(_zz_filter_sampler_sdaSamples_1),
    .CLK(clknet_4_9_0_clock));
 sg13g2_tiehi \_zz_filter_sampler_sdaSamples_1$_SDFFE_PN1P__4  (.L_HI(net3));
 sg13g2_dfrbpq_1 \_zz_filter_sampler_sdaSamples_2$_SDFFE_PN1P_  (.RESET_B(net4),
    .D(_013_),
    .Q(_zz_filter_sampler_sdaSamples_2),
    .CLK(clknet_4_9_0_clock));
 sg13g2_tiehi \_zz_filter_sampler_sdaSamples_2$_SDFFE_PN1P__5  (.L_HI(net4));
 sg13g2_buf_4 clkbuf_0_clock (.X(clknet_0_clock),
    .A(clock));
 sg13g2_buf_8 clkbuf_4_0_0_clock (.A(clknet_0_clock),
    .X(clknet_4_0_0_clock));
 sg13g2_buf_8 clkbuf_4_10_0_clock (.A(clknet_0_clock),
    .X(clknet_4_10_0_clock));
 sg13g2_buf_8 clkbuf_4_11_0_clock (.A(clknet_0_clock),
    .X(clknet_4_11_0_clock));
 sg13g2_buf_8 clkbuf_4_12_0_clock (.A(clknet_0_clock),
    .X(clknet_4_12_0_clock));
 sg13g2_buf_8 clkbuf_4_13_0_clock (.A(clknet_0_clock),
    .X(clknet_4_13_0_clock));
 sg13g2_buf_8 clkbuf_4_14_0_clock (.A(clknet_0_clock),
    .X(clknet_4_14_0_clock));
 sg13g2_buf_8 clkbuf_4_15_0_clock (.A(clknet_0_clock),
    .X(clknet_4_15_0_clock));
 sg13g2_buf_8 clkbuf_4_1_0_clock (.A(clknet_0_clock),
    .X(clknet_4_1_0_clock));
 sg13g2_buf_8 clkbuf_4_2_0_clock (.A(clknet_0_clock),
    .X(clknet_4_2_0_clock));
 sg13g2_buf_8 clkbuf_4_3_0_clock (.A(clknet_0_clock),
    .X(clknet_4_3_0_clock));
 sg13g2_buf_8 clkbuf_4_4_0_clock (.A(clknet_0_clock),
    .X(clknet_4_4_0_clock));
 sg13g2_buf_8 clkbuf_4_5_0_clock (.A(clknet_0_clock),
    .X(clknet_4_5_0_clock));
 sg13g2_buf_8 clkbuf_4_6_0_clock (.A(clknet_0_clock),
    .X(clknet_4_6_0_clock));
 sg13g2_buf_8 clkbuf_4_7_0_clock (.A(clknet_0_clock),
    .X(clknet_4_7_0_clock));
 sg13g2_buf_8 clkbuf_4_8_0_clock (.A(clknet_0_clock),
    .X(clknet_4_8_0_clock));
 sg13g2_buf_8 clkbuf_4_9_0_clock (.A(clknet_0_clock),
    .X(clknet_4_9_0_clock));
 sg13g2_inv_1 clkload0 (.A(clknet_4_7_0_clock));
 sg13g2_inv_1 clkload1 (.A(clknet_4_15_0_clock));
 sg13g2_dfrbpq_1 \ctrl_bitCounter[0]$_SDFFCE_PN1P_  (.RESET_B(net5),
    .D(_014_),
    .Q(\_zz_ctrl_sdaWrite_1[0] ),
    .CLK(clknet_4_3_0_clock));
 sg13g2_tiehi \ctrl_bitCounter[0]$_SDFFCE_PN1P__6  (.L_HI(net5));
 sg13g2_dfrbpq_1 \ctrl_bitCounter[1]$_SDFFCE_PN1P_  (.RESET_B(net6),
    .D(_015_),
    .Q(\_zz_ctrl_sdaWrite_1[1] ),
    .CLK(clknet_4_3_0_clock));
 sg13g2_tiehi \ctrl_bitCounter[1]$_SDFFCE_PN1P__7  (.L_HI(net6));
 sg13g2_dfrbpq_1 \ctrl_bitCounter[2]$_SDFFCE_PN1P_  (.RESET_B(net7),
    .D(_016_),
    .Q(\_zz_ctrl_sdaWrite_1[2] ),
    .CLK(clknet_4_3_0_clock));
 sg13g2_tiehi \ctrl_bitCounter[2]$_SDFFCE_PN1P__8  (.L_HI(net7));
 sg13g2_dfrbpq_1 \ctrl_bitCounter[3]$_SDFFCE_PN1P_  (.RESET_B(net8),
    .D(_017_),
    .Q(\ctrl_bitCounter[3] ),
    .CLK(clknet_4_9_0_clock));
 sg13g2_tiehi \ctrl_bitCounter[3]$_SDFFCE_PN1P__9  (.L_HI(net8));
 sg13g2_dfrbpq_1 \ctrl_bitCounter[4]$_SDFFCE_PN1P_  (.RESET_B(net9),
    .D(_018_),
    .Q(\ctrl_bitCounter[4] ),
    .CLK(clknet_4_1_0_clock));
 sg13g2_tiehi \ctrl_bitCounter[4]$_SDFFCE_PN1P__10  (.L_HI(net9));
 sg13g2_dfrbpq_1 \ctrl_cmdLock$_DFF_P_  (.RESET_B(net10),
    .D(_000_),
    .Q(ctrl_cmdLock),
    .CLK(clknet_4_1_0_clock));
 sg13g2_tiehi \ctrl_cmdLock$_DFF_P__11  (.L_HI(net10));
 sg13g2_dfrbpq_1 \ctrl_frameCounter[0]$_DFF_P_  (.RESET_B(net11),
    .D(_001_),
    .Q(\ctrl_frameCounter[0] ),
    .CLK(clknet_4_4_0_clock));
 sg13g2_tiehi \ctrl_frameCounter[0]$_DFF_P__12  (.L_HI(net11));
 sg13g2_dfrbpq_1 \ctrl_frameCounter[1]$_DFF_P_  (.RESET_B(net12),
    .D(_002_),
    .Q(\ctrl_frameCounter[1] ),
    .CLK(clknet_4_6_0_clock));
 sg13g2_tiehi \ctrl_frameCounter[1]$_DFF_P__13  (.L_HI(net12));
 sg13g2_dfrbpq_1 \ctrl_frameCounter[2]$_DFF_P_  (.RESET_B(net13),
    .D(_003_),
    .Q(\ctrl_frameCounter[2] ),
    .CLK(clknet_4_5_0_clock));
 sg13g2_tiehi \ctrl_frameCounter[2]$_DFF_P__14  (.L_HI(net13));
 sg13g2_dfrbpq_1 \ctrl_frameCounter[3]$_DFF_P_  (.RESET_B(net14),
    .D(_004_),
    .Q(\ctrl_frameCounter[3] ),
    .CLK(clknet_4_6_0_clock));
 sg13g2_tiehi \ctrl_frameCounter[3]$_DFF_P__15  (.L_HI(net14));
 sg13g2_dfrbpq_1 \ctrl_read$_DFF_P_  (.RESET_B(net15),
    .D(_005_),
    .Q(net140),
    .CLK(clknet_4_6_0_clock));
 sg13g2_tiehi \ctrl_read$_DFF_P__16  (.L_HI(net15));
 sg13g2_dfrbpq_1 \ctrl_response_data[0]$_DFFE_PP_  (.RESET_B(net16),
    .D(_019_),
    .Q(\_zz_ctrl_sdaWrite[7] ),
    .CLK(clknet_4_0_0_clock));
 sg13g2_tiehi \ctrl_response_data[0]$_DFFE_PP__17  (.L_HI(net16));
 sg13g2_dfrbpq_1 \ctrl_response_data[1]$_DFFE_PP_  (.RESET_B(net17),
    .D(_020_),
    .Q(\_zz_ctrl_sdaWrite[6] ),
    .CLK(clknet_4_2_0_clock));
 sg13g2_tiehi \ctrl_response_data[1]$_DFFE_PP__18  (.L_HI(net17));
 sg13g2_dfrbpq_1 \ctrl_response_data[2]$_DFFE_PP_  (.RESET_B(net18),
    .D(_021_),
    .Q(\_zz_ctrl_sdaWrite[5] ),
    .CLK(clknet_4_0_0_clock));
 sg13g2_tiehi \ctrl_response_data[2]$_DFFE_PP__19  (.L_HI(net18));
 sg13g2_dfrbpq_1 \ctrl_response_data[3]$_DFFE_PP_  (.RESET_B(net19),
    .D(_022_),
    .Q(\_zz_ctrl_sdaWrite[4] ),
    .CLK(clknet_4_2_0_clock));
 sg13g2_tiehi \ctrl_response_data[3]$_DFFE_PP__20  (.L_HI(net19));
 sg13g2_dfrbpq_1 \ctrl_response_data[4]$_DFFE_PP_  (.RESET_B(net20),
    .D(_023_),
    .Q(\_zz_ctrl_sdaWrite[3] ),
    .CLK(clknet_4_0_0_clock));
 sg13g2_tiehi \ctrl_response_data[4]$_DFFE_PP__21  (.L_HI(net20));
 sg13g2_dfrbpq_1 \ctrl_response_data[5]$_DFFE_PP_  (.RESET_B(net21),
    .D(_024_),
    .Q(\_zz_ctrl_sdaWrite[2] ),
    .CLK(clknet_4_0_0_clock));
 sg13g2_tiehi \ctrl_response_data[5]$_DFFE_PP__22  (.L_HI(net21));
 sg13g2_dfrbpq_1 \ctrl_response_data[6]$_DFFE_PP_  (.RESET_B(net22),
    .D(_025_),
    .Q(\_zz_ctrl_sdaWrite[1] ),
    .CLK(clknet_4_0_0_clock));
 sg13g2_tiehi \ctrl_response_data[6]$_DFFE_PP__23  (.L_HI(net22));
 sg13g2_dfrbpq_1 \ctrl_response_data[7]$_DFFE_PP_  (.RESET_B(net23),
    .D(_026_),
    .Q(\_zz_ctrl_sdaWrite[0] ),
    .CLK(clknet_4_1_0_clock));
 sg13g2_tiehi \ctrl_response_data[7]$_DFFE_PP__24  (.L_HI(net23));
 sg13g2_dfrbpq_1 \ctrl_response_error$_DFF_P_  (.RESET_B(net24),
    .D(_006_),
    .Q(ctrl_response_error),
    .CLK(clknet_4_1_0_clock));
 sg13g2_tiehi \ctrl_response_error$_DFF_P__25  (.L_HI(net24));
 sg13g2_dfrbpq_1 \ctrl_sdaWrite$_SDFF_PN0_  (.RESET_B(net25),
    .D(_027_),
    .Q(net143),
    .CLK(clknet_4_4_0_clock));
 sg13g2_tiehi \ctrl_sdaWrite$_SDFF_PN0__26  (.L_HI(net25));
 sg13g2_dfrbpq_1 \ctrl_shiftRegister[0]$_DFFE_PP_  (.RESET_B(net26),
    .D(_028_),
    .Q(net132),
    .CLK(clknet_4_7_0_clock));
 sg13g2_tiehi \ctrl_shiftRegister[0]$_DFFE_PP__27  (.L_HI(net26));
 sg13g2_dfrbpq_1 \ctrl_shiftRegister[1]$_DFFE_PP_  (.RESET_B(net27),
    .D(_029_),
    .Q(net133),
    .CLK(clknet_4_7_0_clock));
 sg13g2_tiehi \ctrl_shiftRegister[1]$_DFFE_PP__28  (.L_HI(net27));
 sg13g2_dfrbpq_1 \ctrl_shiftRegister[2]$_DFFE_PP_  (.RESET_B(net28),
    .D(_030_),
    .Q(net134),
    .CLK(clknet_4_7_0_clock));
 sg13g2_tiehi \ctrl_shiftRegister[2]$_DFFE_PP__29  (.L_HI(net28));
 sg13g2_dfrbpq_1 \ctrl_shiftRegister[3]$_DFFE_PP_  (.RESET_B(net29),
    .D(_031_),
    .Q(net135),
    .CLK(clknet_4_5_0_clock));
 sg13g2_tiehi \ctrl_shiftRegister[3]$_DFFE_PP__30  (.L_HI(net29));
 sg13g2_dfrbpq_1 \ctrl_shiftRegister[4]$_DFFE_PP_  (.RESET_B(net30),
    .D(_032_),
    .Q(net136),
    .CLK(clknet_4_4_0_clock));
 sg13g2_tiehi \ctrl_shiftRegister[4]$_DFFE_PP__31  (.L_HI(net30));
 sg13g2_dfrbpq_1 \ctrl_shiftRegister[5]$_DFFE_PP_  (.RESET_B(net31),
    .D(_033_),
    .Q(net137),
    .CLK(clknet_4_5_0_clock));
 sg13g2_tiehi \ctrl_shiftRegister[5]$_DFFE_PP__32  (.L_HI(net31));
 sg13g2_dfrbpq_1 \ctrl_shiftRegister[6]$_DFFE_PP_  (.RESET_B(net32),
    .D(_034_),
    .Q(net138),
    .CLK(clknet_4_5_0_clock));
 sg13g2_tiehi \ctrl_shiftRegister[6]$_DFFE_PP__33  (.L_HI(net32));
 sg13g2_dfrbpq_1 \ctrl_shiftRegister[7]$_DFFE_PP_  (.RESET_B(net33),
    .D(_035_),
    .Q(net139),
    .CLK(clknet_4_5_0_clock));
 sg13g2_tiehi \ctrl_shiftRegister[7]$_DFFE_PP__34  (.L_HI(net33));
 sg13g2_dfrbpq_1 \ctrl_state[0]$_DFF_P_  (.RESET_B(net34),
    .D(_007_),
    .Q(\ctrl_state[0] ),
    .CLK(clknet_4_4_0_clock));
 sg13g2_tiehi \ctrl_state[0]$_DFF_P__35  (.L_HI(net34));
 sg13g2_dfrbpq_1 \ctrl_state[1]$_DFF_P_  (.RESET_B(net35),
    .D(_008_),
    .Q(\ctrl_state[1] ),
    .CLK(clknet_4_1_0_clock));
 sg13g2_tiehi \ctrl_state[1]$_DFF_P__36  (.L_HI(net35));
 sg13g2_dfrbpq_1 \ctrl_state[2]$_DFF_P_  (.RESET_B(net36),
    .D(_009_),
    .Q(net142),
    .CLK(clknet_4_4_0_clock));
 sg13g2_tiehi \ctrl_state[2]$_DFF_P__37  (.L_HI(net36));
 sg13g2_dfrbpq_1 \ctrl_transmission$_SDFFE_PN0P_  (.RESET_B(net37),
    .D(_036_),
    .Q(ctrl_transmission),
    .CLK(clknet_4_12_0_clock));
 sg13g2_tiehi \ctrl_transmission$_SDFFE_PN0P__38  (.L_HI(net37));
 sg13g2_dfrbpq_1 \filter_scl$_SDFFE_PN1P_  (.RESET_B(net38),
    .D(_037_),
    .Q(filter_scl),
    .CLK(clknet_4_9_0_clock));
 sg13g2_tiehi \filter_scl$_SDFFE_PN1P__39  (.L_HI(net38));
 sg13g2_dfrbpq_1 \filter_scl_regNext$_SDFF_PN1_  (.RESET_B(net39),
    .D(_038_),
    .Q(filter_scl_regNext),
    .CLK(clknet_4_12_0_clock));
 sg13g2_tiehi \filter_scl_regNext$_SDFF_PN1__40  (.L_HI(net39));
 sg13g2_dfrbpq_1 \filter_sda$_SDFFE_PN1P_  (.RESET_B(net40),
    .D(_039_),
    .Q(filter_sda),
    .CLK(clknet_4_12_0_clock));
 sg13g2_tiehi \filter_sda$_SDFFE_PN1P__41  (.L_HI(net40));
 sg13g2_dfrbpq_1 \filter_sda_regNext$_SDFF_PN1_  (.RESET_B(net41),
    .D(_040_),
    .Q(filter_sda_regNext),
    .CLK(clknet_4_12_0_clock));
 sg13g2_tiehi \filter_sda_regNext$_SDFF_PN1__42  (.L_HI(net41));
 sg13g2_dfrbpq_1 \filter_timer_counter[0]$_SDFF_PN0_  (.RESET_B(net42),
    .D(_041_),
    .Q(\filter_timer_counter[0] ),
    .CLK(clknet_4_2_0_clock));
 sg13g2_tiehi \filter_timer_counter[0]$_SDFF_PN0__43  (.L_HI(net42));
 sg13g2_dfrbpq_1 \filter_timer_counter[10]$_SDFF_PN0_  (.RESET_B(net43),
    .D(_042_),
    .Q(\filter_timer_counter[10] ),
    .CLK(clknet_4_14_0_clock));
 sg13g2_tiehi \filter_timer_counter[10]$_SDFF_PN0__44  (.L_HI(net43));
 sg13g2_dfrbpq_1 \filter_timer_counter[11]$_SDFF_PN0_  (.RESET_B(net44),
    .D(_043_),
    .Q(\filter_timer_counter[11] ),
    .CLK(clknet_4_11_0_clock));
 sg13g2_tiehi \filter_timer_counter[11]$_SDFF_PN0__45  (.L_HI(net44));
 sg13g2_dfrbpq_1 \filter_timer_counter[12]$_SDFF_PN0_  (.RESET_B(net45),
    .D(_044_),
    .Q(\filter_timer_counter[12] ),
    .CLK(clknet_4_11_0_clock));
 sg13g2_tiehi \filter_timer_counter[12]$_SDFF_PN0__46  (.L_HI(net45));
 sg13g2_dfrbpq_1 \filter_timer_counter[13]$_SDFF_PN0_  (.RESET_B(net46),
    .D(_045_),
    .Q(\filter_timer_counter[13] ),
    .CLK(clknet_4_11_0_clock));
 sg13g2_tiehi \filter_timer_counter[13]$_SDFF_PN0__47  (.L_HI(net46));
 sg13g2_dfrbpq_1 \filter_timer_counter[14]$_SDFF_PN0_  (.RESET_B(net47),
    .D(_046_),
    .Q(\filter_timer_counter[14] ),
    .CLK(clknet_4_11_0_clock));
 sg13g2_tiehi \filter_timer_counter[14]$_SDFF_PN0__48  (.L_HI(net47));
 sg13g2_dfrbpq_1 \filter_timer_counter[15]$_SDFF_PN0_  (.RESET_B(net48),
    .D(_047_),
    .Q(\filter_timer_counter[15] ),
    .CLK(clknet_4_11_0_clock));
 sg13g2_tiehi \filter_timer_counter[15]$_SDFF_PN0__49  (.L_HI(net48));
 sg13g2_dfrbpq_1 \filter_timer_counter[1]$_SDFF_PN0_  (.RESET_B(net49),
    .D(_048_),
    .Q(\filter_timer_counter[1] ),
    .CLK(clknet_4_8_0_clock));
 sg13g2_tiehi \filter_timer_counter[1]$_SDFF_PN0__50  (.L_HI(net49));
 sg13g2_dfrbpq_1 \filter_timer_counter[2]$_SDFF_PN0_  (.RESET_B(net50),
    .D(_049_),
    .Q(\filter_timer_counter[2] ),
    .CLK(clknet_4_8_0_clock));
 sg13g2_tiehi \filter_timer_counter[2]$_SDFF_PN0__51  (.L_HI(net50));
 sg13g2_dfrbpq_1 \filter_timer_counter[3]$_SDFF_PN0_  (.RESET_B(net51),
    .D(_050_),
    .Q(\filter_timer_counter[3] ),
    .CLK(clknet_4_8_0_clock));
 sg13g2_tiehi \filter_timer_counter[3]$_SDFF_PN0__52  (.L_HI(net51));
 sg13g2_dfrbpq_1 \filter_timer_counter[4]$_SDFF_PN0_  (.RESET_B(net52),
    .D(_051_),
    .Q(\filter_timer_counter[4] ),
    .CLK(clknet_4_10_0_clock));
 sg13g2_tiehi \filter_timer_counter[4]$_SDFF_PN0__53  (.L_HI(net52));
 sg13g2_dfrbpq_1 \filter_timer_counter[5]$_SDFF_PN0_  (.RESET_B(net53),
    .D(_052_),
    .Q(\filter_timer_counter[5] ),
    .CLK(clknet_4_10_0_clock));
 sg13g2_tiehi \filter_timer_counter[5]$_SDFF_PN0__54  (.L_HI(net53));
 sg13g2_dfrbpq_1 \filter_timer_counter[6]$_SDFF_PN0_  (.RESET_B(net54),
    .D(_053_),
    .Q(\filter_timer_counter[6] ),
    .CLK(clknet_4_10_0_clock));
 sg13g2_tiehi \filter_timer_counter[6]$_SDFF_PN0__55  (.L_HI(net54));
 sg13g2_dfrbpq_1 \filter_timer_counter[7]$_SDFF_PN0_  (.RESET_B(net55),
    .D(_054_),
    .Q(\filter_timer_counter[7] ),
    .CLK(clknet_4_10_0_clock));
 sg13g2_tiehi \filter_timer_counter[7]$_SDFF_PN0__56  (.L_HI(net55));
 sg13g2_dfrbpq_1 \filter_timer_counter[8]$_SDFF_PN0_  (.RESET_B(net56),
    .D(_055_),
    .Q(\filter_timer_counter[8] ),
    .CLK(clknet_4_10_0_clock));
 sg13g2_tiehi \filter_timer_counter[8]$_SDFF_PN0__57  (.L_HI(net56));
 sg13g2_dfrbpq_1 \filter_timer_counter[9]$_SDFF_PN0_  (.RESET_B(net57),
    .D(_056_),
    .Q(\filter_timer_counter[9] ),
    .CLK(clknet_4_8_0_clock));
 sg13g2_tiehi \filter_timer_counter[9]$_SDFF_PN0__58  (.L_HI(net57));
 sg13g2_buf_1 input100 (.A(io_config_deviceAddr[3]),
    .X(net99));
 sg13g2_buf_1 input101 (.A(io_config_deviceAddr[4]),
    .X(net100));
 sg13g2_buf_1 input102 (.A(io_config_deviceAddr[5]),
    .X(net101));
 sg13g2_buf_1 input103 (.A(io_config_deviceAddr[6]),
    .X(net102));
 sg13g2_buf_1 input104 (.A(io_config_timeout[0]),
    .X(net103));
 sg13g2_buf_1 input105 (.A(io_config_timeout[10]),
    .X(net104));
 sg13g2_buf_1 input106 (.A(io_config_timeout[11]),
    .X(net105));
 sg13g2_buf_1 input107 (.A(io_config_timeout[12]),
    .X(net106));
 sg13g2_buf_1 input108 (.A(io_config_timeout[13]),
    .X(net107));
 sg13g2_buf_1 input109 (.A(io_config_timeout[14]),
    .X(net108));
 sg13g2_buf_1 input110 (.A(io_config_timeout[15]),
    .X(net109));
 sg13g2_buf_1 input111 (.A(io_config_timeout[1]),
    .X(net110));
 sg13g2_buf_1 input112 (.A(io_config_timeout[2]),
    .X(net111));
 sg13g2_buf_1 input113 (.A(io_config_timeout[3]),
    .X(net112));
 sg13g2_buf_1 input114 (.A(io_config_timeout[4]),
    .X(net113));
 sg13g2_buf_1 input115 (.A(io_config_timeout[5]),
    .X(net114));
 sg13g2_buf_1 input116 (.A(io_config_timeout[6]),
    .X(net115));
 sg13g2_buf_1 input117 (.A(io_config_timeout[7]),
    .X(net116));
 sg13g2_buf_1 input118 (.A(io_config_timeout[8]),
    .X(net117));
 sg13g2_buf_1 input119 (.A(io_config_timeout[9]),
    .X(net118));
 sg13g2_buf_1 input120 (.A(io_i2c_scl_read),
    .X(net119));
 sg13g2_buf_1 input121 (.A(io_i2c_sda_read),
    .X(net120));
 sg13g2_buf_1 input122 (.A(io_rsp_payload_data[0]),
    .X(net121));
 sg13g2_buf_1 input123 (.A(io_rsp_payload_data[1]),
    .X(net122));
 sg13g2_buf_1 input124 (.A(io_rsp_payload_data[2]),
    .X(net123));
 sg13g2_buf_1 input125 (.A(io_rsp_payload_data[3]),
    .X(net124));
 sg13g2_buf_1 input126 (.A(io_rsp_payload_data[4]),
    .X(net125));
 sg13g2_buf_1 input127 (.A(io_rsp_payload_data[5]),
    .X(net126));
 sg13g2_buf_1 input128 (.A(io_rsp_payload_data[6]),
    .X(net127));
 sg13g2_buf_1 input129 (.A(io_rsp_payload_data[7]),
    .X(net128));
 sg13g2_buf_1 input130 (.A(io_rsp_payload_error),
    .X(net129));
 sg13g2_buf_1 input131 (.A(io_rsp_valid),
    .X(net130));
 sg13g2_buf_1 input132 (.A(reset),
    .X(net131));
 sg13g2_buf_1 input80 (.A(io_cmd_ready),
    .X(net79));
 sg13g2_buf_1 input81 (.A(io_config_clockDivider[0]),
    .X(net80));
 sg13g2_buf_1 input82 (.A(io_config_clockDivider[10]),
    .X(net81));
 sg13g2_buf_1 input83 (.A(io_config_clockDivider[11]),
    .X(net82));
 sg13g2_buf_1 input84 (.A(io_config_clockDivider[12]),
    .X(net83));
 sg13g2_buf_1 input85 (.A(io_config_clockDivider[13]),
    .X(net84));
 sg13g2_buf_1 input86 (.A(io_config_clockDivider[14]),
    .X(net85));
 sg13g2_buf_1 input87 (.A(io_config_clockDivider[15]),
    .X(net86));
 sg13g2_buf_1 input88 (.A(io_config_clockDivider[1]),
    .X(net87));
 sg13g2_buf_1 input89 (.A(io_config_clockDivider[2]),
    .X(net88));
 sg13g2_buf_1 input90 (.A(io_config_clockDivider[3]),
    .X(net89));
 sg13g2_buf_1 input91 (.A(io_config_clockDivider[4]),
    .X(net90));
 sg13g2_buf_1 input92 (.A(io_config_clockDivider[5]),
    .X(net91));
 sg13g2_buf_1 input93 (.A(io_config_clockDivider[6]),
    .X(net92));
 sg13g2_buf_1 input94 (.A(io_config_clockDivider[7]),
    .X(net93));
 sg13g2_buf_1 input95 (.A(io_config_clockDivider[8]),
    .X(net94));
 sg13g2_buf_1 input96 (.A(io_config_clockDivider[9]),
    .X(net95));
 sg13g2_buf_1 input97 (.A(io_config_deviceAddr[0]),
    .X(net96));
 sg13g2_buf_1 input98 (.A(io_config_deviceAddr[1]),
    .X(net97));
 sg13g2_buf_1 input99 (.A(io_config_deviceAddr[2]),
    .X(net98));
 sg13g2_nand2b_1 \io_i2c_scl_read_buffercc/_3_  (.Y(\io_i2c_scl_read_buffercc/_0_ ),
    .B(net131),
    .A_N(net119));
 sg13g2_nand2b_1 \io_i2c_scl_read_buffercc/_4_  (.Y(\io_i2c_scl_read_buffercc/_1_ ),
    .B(net200),
    .A_N(\io_i2c_scl_read_buffercc/buffers_0 ));
 sg13g2_dfrbpq_1 \io_i2c_scl_read_buffercc/buffers_0$_SDFF_PN1_  (.RESET_B(net75),
    .D(\io_i2c_scl_read_buffercc/_0_ ),
    .Q(\io_i2c_scl_read_buffercc/buffers_0 ),
    .CLK(clknet_4_2_0_clock));
 sg13g2_tiehi \io_i2c_scl_read_buffercc/buffers_0$_SDFF_PN1__76  (.L_HI(net75));
 sg13g2_dfrbpq_1 \io_i2c_scl_read_buffercc/buffers_1$_SDFF_PN1_  (.RESET_B(net76),
    .D(\io_i2c_scl_read_buffercc/_1_ ),
    .Q(_zz_filter_sampler_sclSamples_0),
    .CLK(clknet_4_3_0_clock));
 sg13g2_tiehi \io_i2c_scl_read_buffercc/buffers_1$_SDFF_PN1__77  (.L_HI(net76));
 sg13g2_nand2b_1 \io_i2c_sda_read_buffercc/_3_  (.Y(\io_i2c_sda_read_buffercc/_0_ ),
    .B(net131),
    .A_N(net120));
 sg13g2_nand2b_1 \io_i2c_sda_read_buffercc/_4_  (.Y(\io_i2c_sda_read_buffercc/_1_ ),
    .B(net199),
    .A_N(\io_i2c_sda_read_buffercc/buffers_0 ));
 sg13g2_dfrbpq_1 \io_i2c_sda_read_buffercc/buffers_0$_SDFF_PN1_  (.RESET_B(net77),
    .D(\io_i2c_sda_read_buffercc/_0_ ),
    .Q(\io_i2c_sda_read_buffercc/buffers_0 ),
    .CLK(clknet_4_2_0_clock));
 sg13g2_tiehi \io_i2c_sda_read_buffercc/buffers_0$_SDFF_PN1__78  (.L_HI(net77));
 sg13g2_dfrbpq_1 \io_i2c_sda_read_buffercc/buffers_1$_SDFF_PN1_  (.RESET_B(net78),
    .D(\io_i2c_sda_read_buffercc/_1_ ),
    .Q(_zz_filter_sampler_sdaSamples_0),
    .CLK(clknet_4_3_0_clock));
 sg13g2_tiehi \io_i2c_sda_read_buffercc/buffers_1$_SDFF_PN1__79  (.L_HI(net78));
 sg13g2_buf_1 output133 (.A(net132),
    .X(io_cmd_payload_data[0]));
 sg13g2_buf_1 output134 (.A(net133),
    .X(io_cmd_payload_data[1]));
 sg13g2_buf_1 output135 (.A(net134),
    .X(io_cmd_payload_data[2]));
 sg13g2_buf_1 output136 (.A(net135),
    .X(io_cmd_payload_data[3]));
 sg13g2_buf_1 output137 (.A(net136),
    .X(io_cmd_payload_data[4]));
 sg13g2_buf_1 output138 (.A(net137),
    .X(io_cmd_payload_data[5]));
 sg13g2_buf_1 output139 (.A(net138),
    .X(io_cmd_payload_data[6]));
 sg13g2_buf_1 output140 (.A(net139),
    .X(io_cmd_payload_data[7]));
 sg13g2_buf_1 output141 (.A(net140),
    .X(io_cmd_payload_read));
 sg13g2_buf_1 output142 (.A(net141),
    .X(io_cmd_payload_reg));
 sg13g2_buf_1 output143 (.A(net142),
    .X(io_cmd_valid));
 sg13g2_buf_1 output144 (.A(net143),
    .X(io_i2c_sda_write));
 sg13g2_buf_1 output145 (.A(net144),
    .X(io_rsp_ready));
 sg13g2_buf_1 place186 (.A(net186),
    .X(net185));
 sg13g2_buf_1 place187 (.A(_294_),
    .X(net186));
 sg13g2_buf_1 place188 (.A(_288_),
    .X(net187));
 sg13g2_buf_1 place189 (.A(_209_),
    .X(net188));
 sg13g2_buf_1 place190 (.A(_203_),
    .X(net189));
 sg13g2_buf_1 place191 (.A(_301_),
    .X(net190));
 sg13g2_buf_1 place192 (.A(_148_),
    .X(net191));
 sg13g2_buf_1 place193 (.A(net144),
    .X(net192));
 sg13g2_buf_1 place194 (.A(\filter_timer_counter[12] ),
    .X(net193));
 sg13g2_buf_1 place195 (.A(filter_scl),
    .X(net194));
 sg13g2_buf_1 place196 (.A(\ctrl_frameCounter[0] ),
    .X(net195));
 sg13g2_buf_1 place197 (.A(\_zz_ctrl_sdaWrite_1[0] ),
    .X(net196));
 sg13g2_buf_1 place198 (.A(net198),
    .X(net197));
 sg13g2_buf_1 place199 (.A(_116_),
    .X(net198));
 sg13g2_buf_1 place200 (.A(net200),
    .X(net199));
 sg13g2_buf_1 place201 (.A(net131),
    .X(net200));
 sg13g2_dfrbpq_1 \timeout_transmission$_SDFFE_PP0P_  (.RESET_B(net58),
    .D(_057_),
    .Q(timeout_transmission),
    .CLK(clknet_4_12_0_clock));
 sg13g2_tiehi \timeout_transmission$_SDFFE_PP0P__59  (.L_HI(net58));
 sg13g2_dfrbpq_1 \timeout_value[0]$_SDFFE_PN0P_  (.RESET_B(net59),
    .D(_058_),
    .Q(\timeout_value[0] ),
    .CLK(clknet_4_7_0_clock));
 sg13g2_tiehi \timeout_value[0]$_SDFFE_PN0P__60  (.L_HI(net59));
 sg13g2_dfrbpq_1 \timeout_value[10]$_SDFFE_PN0P_  (.RESET_B(net60),
    .D(_059_),
    .Q(\timeout_value[10] ),
    .CLK(clknet_4_13_0_clock));
 sg13g2_tiehi \timeout_value[10]$_SDFFE_PN0P__61  (.L_HI(net60));
 sg13g2_dfrbpq_1 \timeout_value[11]$_SDFFE_PN0P_  (.RESET_B(net61),
    .D(_060_),
    .Q(\timeout_value[11] ),
    .CLK(clknet_4_13_0_clock));
 sg13g2_tiehi \timeout_value[11]$_SDFFE_PN0P__62  (.L_HI(net61));
 sg13g2_dfrbpq_1 \timeout_value[12]$_SDFFE_PN0P_  (.RESET_B(net62),
    .D(_061_),
    .Q(\timeout_value[12] ),
    .CLK(clknet_4_14_0_clock));
 sg13g2_tiehi \timeout_value[12]$_SDFFE_PN0P__63  (.L_HI(net62));
 sg13g2_dfrbpq_1 \timeout_value[13]$_SDFFE_PN0P_  (.RESET_B(net63),
    .D(_062_),
    .Q(\timeout_value[13] ),
    .CLK(clknet_4_14_0_clock));
 sg13g2_tiehi \timeout_value[13]$_SDFFE_PN0P__64  (.L_HI(net63));
 sg13g2_dfrbpq_1 \timeout_value[14]$_SDFFE_PN0P_  (.RESET_B(net64),
    .D(_063_),
    .Q(\timeout_value[14] ),
    .CLK(clknet_4_14_0_clock));
 sg13g2_tiehi \timeout_value[14]$_SDFFE_PN0P__65  (.L_HI(net64));
 sg13g2_dfrbpq_1 \timeout_value[15]$_SDFFE_PN0P_  (.RESET_B(net65),
    .D(_064_),
    .Q(\timeout_value[15] ),
    .CLK(clknet_4_15_0_clock));
 sg13g2_tiehi \timeout_value[15]$_SDFFE_PN0P__66  (.L_HI(net65));
 sg13g2_dfrbpq_1 \timeout_value[1]$_SDFFE_PN0P_  (.RESET_B(net66),
    .D(_065_),
    .Q(\timeout_value[1] ),
    .CLK(clknet_4_6_0_clock));
 sg13g2_tiehi \timeout_value[1]$_SDFFE_PN0P__67  (.L_HI(net66));
 sg13g2_dfrbpq_1 \timeout_value[2]$_SDFFE_PN0P_  (.RESET_B(net67),
    .D(_066_),
    .Q(\timeout_value[2] ),
    .CLK(clknet_4_6_0_clock));
 sg13g2_tiehi \timeout_value[2]$_SDFFE_PN0P__68  (.L_HI(net67));
 sg13g2_dfrbpq_1 \timeout_value[3]$_SDFFE_PN0P_  (.RESET_B(net68),
    .D(_067_),
    .Q(\timeout_value[3] ),
    .CLK(clknet_4_13_0_clock));
 sg13g2_tiehi \timeout_value[3]$_SDFFE_PN0P__69  (.L_HI(net68));
 sg13g2_dfrbpq_1 \timeout_value[4]$_SDFFE_PN0P_  (.RESET_B(net69),
    .D(_068_),
    .Q(\timeout_value[4] ),
    .CLK(clknet_4_15_0_clock));
 sg13g2_tiehi \timeout_value[4]$_SDFFE_PN0P__70  (.L_HI(net69));
 sg13g2_dfrbpq_1 \timeout_value[5]$_SDFFE_PN0P_  (.RESET_B(net70),
    .D(_069_),
    .Q(\timeout_value[5] ),
    .CLK(clknet_4_15_0_clock));
 sg13g2_tiehi \timeout_value[5]$_SDFFE_PN0P__71  (.L_HI(net70));
 sg13g2_dfrbpq_1 \timeout_value[6]$_SDFFE_PN0P_  (.RESET_B(net71),
    .D(_070_),
    .Q(\timeout_value[6] ),
    .CLK(clknet_4_15_0_clock));
 sg13g2_tiehi \timeout_value[6]$_SDFFE_PN0P__72  (.L_HI(net71));
 sg13g2_dfrbpq_1 \timeout_value[7]$_SDFFE_PN0P_  (.RESET_B(net72),
    .D(_071_),
    .Q(\timeout_value[7] ),
    .CLK(clknet_4_14_0_clock));
 sg13g2_tiehi \timeout_value[7]$_SDFFE_PN0P__73  (.L_HI(net72));
 sg13g2_dfrbpq_1 \timeout_value[8]$_SDFFE_PN0P_  (.RESET_B(net73),
    .D(_072_),
    .Q(\timeout_value[8] ),
    .CLK(clknet_4_13_0_clock));
 sg13g2_tiehi \timeout_value[8]$_SDFFE_PN0P__74  (.L_HI(net73));
 sg13g2_dfrbpq_1 \timeout_value[9]$_SDFFE_PN0P_  (.RESET_B(net74),
    .D(_073_),
    .Q(\timeout_value[9] ),
    .CLK(clknet_4_13_0_clock));
 sg13g2_tiehi \timeout_value[9]$_SDFFE_PN0P__75  (.L_HI(net74));
 assign io_i2c_interrupts[0] = io_interrupts[0];
endmodule
