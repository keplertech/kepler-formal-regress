module aes_cipher_top (clk,
    done,
    ld,
    rst,
    key,
    text_in,
    text_out);
 input clk;
 output done;
 input ld;
 input rst;
 input [127:0] key;
 input [127:0] text_in;
 output [127:0] text_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire net4738;
 wire net4736;
 wire net4733;
 wire net4734;
 wire net4774;
 wire net4820;
 wire net4818;
 wire net4815;
 wire net4814;
 wire net4730;
 wire net4775;
 wire net4729;
 wire net4751;
 wire net4753;
 wire net4747;
 wire net4745;
 wire net4742;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire net4822;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire net4811;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire net4741;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire net4744;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire net4740;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire net4702;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire net4752;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire net4750;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire net4684;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire net4755;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire net4683;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire net4754;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire net4646;
 wire net4625;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01067_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire net4644;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire net4647;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire net4616;
 wire net4591;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01088_;
 wire net4617;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire net4611;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire net4571;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire net4580;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire net4569;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire net4573;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire net4517;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire net4522;
 wire _01130_;
 wire net4520;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire net4521;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire net4518;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire net4480;
 wire net4474;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire net4482;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire net4481;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire net4426;
 wire net6322;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire net4432;
 wire _01172_;
 wire net4429;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire net4438;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire net4427;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire net5942;
 wire net5793;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire net5982;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire net5945;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire net5960;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire net5746;
 wire net5663;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire net5742;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire net5744;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire net5436;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01266_;
 wire _01267_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01289_;
 wire _01290_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01312_;
 wire _01313_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01327_;
 wire _01328_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01334_;
 wire _01335_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01348_;
 wire _01349_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01355_;
 wire _01356_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01369_;
 wire _01370_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01376_;
 wire _01377_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01397_;
 wire _01398_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire net5743;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire net5775;
 wire net5774;
 wire net5740;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire net5739;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire net5735;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire net5725;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire net5711;
 wire _01739_;
 wire net5689;
 wire _01741_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire net5683;
 wire _01750_;
 wire _01752_;
 wire _01753_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire net5674;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire net5664;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01789_;
 wire _01790_;
 wire net5659;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire net5658;
 wire net5657;
 wire _01797_;
 wire _01798_;
 wire net5644;
 wire net5653;
 wire _01801_;
 wire _01802_;
 wire net5639;
 wire _01804_;
 wire net5638;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire net5623;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire net5609;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01861_;
 wire _01862_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01874_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire net5480;
 wire _01911_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02023_;
 wire _02024_;
 wire _02026_;
 wire _02027_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire net5156;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02398_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02416_;
 wire _02417_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02462_;
 wire _02463_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02494_;
 wire _02495_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02538_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03080_;
 wire _03082_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03121_;
 wire _03123_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03165_;
 wire _03166_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03181_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03210_;
 wire _03211_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03755_;
 wire _03756_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03791_;
 wire _03793_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03807_;
 wire _03809_;
 wire _03810_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03825_;
 wire _03826_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03861_;
 wire _03862_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03894_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03928_;
 wire _03929_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03942_;
 wire _03943_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04471_;
 wire _04472_;
 wire _04474_;
 wire _04475_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04485_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04509_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04526_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04580_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04675_;
 wire _04676_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05130_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05142_;
 wire _05143_;
 wire _05146_;
 wire _05147_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05159_;
 wire _05161_;
 wire _05162_;
 wire _05165_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05189_;
 wire _05190_;
 wire _05193_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05199_;
 wire _05200_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05209_;
 wire _05210_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05278_;
 wire _05279_;
 wire _05281_;
 wire _05283_;
 wire _05284_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05819_;
 wire _05820_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05828_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05855_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05882_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05899_;
 wire _05902_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06504_;
 wire _06505_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06520_;
 wire _06522_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06558_;
 wire _06560_;
 wire _06563_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06575_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06592_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06601_;
 wire _06602_;
 wire _06605_;
 wire _06606_;
 wire _06609_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06618_;
 wire _06619_;
 wire _06621_;
 wire _06622_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06654_;
 wire _06656_;
 wire _06657_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07196_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07219_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07258_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07270_;
 wire _07271_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07278_;
 wire _07279_;
 wire _07282_;
 wire _07283_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07774_;
 wire _07775_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07786_;
 wire _07787_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07799_;
 wire _07800_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07811_;
 wire _07812_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07823_;
 wire _07824_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07835_;
 wire _07836_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07847_;
 wire _07848_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07859_;
 wire _07860_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07871_;
 wire _07872_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07883_;
 wire _07884_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07895_;
 wire _07896_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire net4864;
 wire net4863;
 wire net4862;
 wire net4861;
 wire net4860;
 wire net4859;
 wire net4858;
 wire net4857;
 wire net4856;
 wire net4855;
 wire net4854;
 wire net4853;
 wire net4850;
 wire net4851;
 wire net4852;
 wire net4849;
 wire net4848;
 wire net4847;
 wire net4845;
 wire net4846;
 wire net4844;
 wire net4841;
 wire net4842;
 wire net4840;
 wire net4843;
 wire net4839;
 wire net4838;
 wire net4835;
 wire net4834;
 wire net4836;
 wire net4837;
 wire net4833;
 wire net4832;
 wire net4831;
 wire net4828;
 wire net4829;
 wire net4830;
 wire net4827;
 wire net4825;
 wire net4826;
 wire net4824;
 wire _08030_;
 wire net4823;
 wire _08035_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08060_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire net4821;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire net4819;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire net4816;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire net4813;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire net4810;
 wire _08107_;
 wire _08108_;
 wire net4812;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire net4809;
 wire _08124_;
 wire net4807;
 wire net4806;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire net4804;
 wire _08134_;
 wire net4805;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire net4803;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire net4808;
 wire _08147_;
 wire _08148_;
 wire net4802;
 wire _08150_;
 wire _08151_;
 wire net4817;
 wire _08153_;
 wire net4801;
 wire net4800;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08161_;
 wire net4799;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire net4798;
 wire net4797;
 wire _08168_;
 wire _08169_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire net4796;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire net4794;
 wire _08195_;
 wire _08196_;
 wire net4793;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire net4792;
 wire _08204_;
 wire net4790;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire net4789;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire net4795;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire net4791;
 wire _08239_;
 wire _08240_;
 wire net4788;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire net4787;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire net4784;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire net4782;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire net4783;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire net4785;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire net4786;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire net4779;
 wire net4778;
 wire net4777;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire net4776;
 wire _08653_;
 wire _08654_;
 wire net4780;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire net4781;
 wire _08676_;
 wire _08677_;
 wire net4773;
 wire _08679_;
 wire _08680_;
 wire net4771;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire net4770;
 wire net4769;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire net4768;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire net4772;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire net4767;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire net4765;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire net4764;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire net4761;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire net4763;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire net4762;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire net4759;
 wire _08828_;
 wire _08829_;
 wire net4757;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire net4756;
 wire _08856_;
 wire _08857_;
 wire net4766;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire net4758;
 wire _08904_;
 wire _08905_;
 wire net4760;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire net4749;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire net4748;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire net4746;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire net4743;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire net4739;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire net4737;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire net4735;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire net4732;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire net4731;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire net4728;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire net4727;
 wire net4726;
 wire _09039_;
 wire _09040_;
 wire net4725;
 wire _09042_;
 wire _09043_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire net4724;
 wire net4722;
 wire _09057_;
 wire net4721;
 wire net4717;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire net4715;
 wire _09068_;
 wire net4716;
 wire net4714;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire net4718;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire net4713;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire net4712;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire net4711;
 wire _09100_;
 wire net4719;
 wire _09102_;
 wire _09103_;
 wire net4720;
 wire _09105_;
 wire net4710;
 wire _09107_;
 wire net4709;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire net4723;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire net4708;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire net4707;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire net4706;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09191_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire net4705;
 wire _09212_;
 wire net4704;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09235_;
 wire _09236_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire net4703;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire net4701;
 wire net4700;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire net4699;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire net4698;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09593_;
 wire _09594_;
 wire net4697;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire net4696;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09611_;
 wire _09612_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire net4695;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire net4694;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire net4693;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09648_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire net4692;
 wire net4691;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire net4690;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire net4689;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire net4688;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire net4687;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire net4686;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire net4685;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire net4681;
 wire net4682;
 wire _10118_;
 wire _10119_;
 wire net4680;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire net4677;
 wire _10133_;
 wire _10134_;
 wire net4676;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire net4675;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire net4674;
 wire _10149_;
 wire net4673;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire net4678;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire net4672;
 wire _10168_;
 wire net4679;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire net4671;
 wire _10176_;
 wire net4670;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire net4669;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire net4667;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire net4668;
 wire _10212_;
 wire _10213_;
 wire net4666;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10226_;
 wire net4665;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10258_;
 wire _10259_;
 wire net4664;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire net4661;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire net4662;
 wire _10295_;
 wire net4658;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire net4660;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire net4659;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire net4656;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire net4657;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire _10563_;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire _10582_;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire _10602_;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire _10609_;
 wire _10610_;
 wire _10611_;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire _10618_;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire _10632_;
 wire _10633_;
 wire _10634_;
 wire _10635_;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire _10652_;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire net4663;
 wire net4655;
 wire net4654;
 wire _10675_;
 wire _10676_;
 wire net4653;
 wire net4652;
 wire _10679_;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire net4651;
 wire _10689_;
 wire net4650;
 wire _10691_;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire net4649;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10727_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire net4648;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire _10741_;
 wire net4645;
 wire _10743_;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire net4643;
 wire net4642;
 wire _10750_;
 wire _10751_;
 wire _10752_;
 wire _10753_;
 wire _10756_;
 wire _10757_;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10765_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10773_;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10780_;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire _10787_;
 wire net4641;
 wire _10790_;
 wire _10791_;
 wire net4639;
 wire _10793_;
 wire _10794_;
 wire net4638;
 wire _10796_;
 wire _10797_;
 wire _10798_;
 wire _10799_;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire _10807_;
 wire _10808_;
 wire _10809_;
 wire _10810_;
 wire _10811_;
 wire _10812_;
 wire _10813_;
 wire _10814_;
 wire net4636;
 wire net4635;
 wire _10817_;
 wire _10818_;
 wire net4634;
 wire net4633;
 wire _10821_;
 wire _10822_;
 wire net4637;
 wire _10824_;
 wire _10825_;
 wire _10826_;
 wire _10827_;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire _10831_;
 wire _10832_;
 wire _10833_;
 wire _10834_;
 wire _10835_;
 wire _10836_;
 wire net4632;
 wire net4640;
 wire _10839_;
 wire _10840_;
 wire _10841_;
 wire _10842_;
 wire _10843_;
 wire _10844_;
 wire net4631;
 wire _10847_;
 wire _10848_;
 wire _10849_;
 wire _10850_;
 wire _10852_;
 wire net4630;
 wire _10854_;
 wire _10855_;
 wire _10856_;
 wire _10857_;
 wire _10858_;
 wire _10859_;
 wire _10860_;
 wire _10861_;
 wire net4629;
 wire net4628;
 wire net4626;
 wire _10865_;
 wire _10866_;
 wire _10867_;
 wire _10868_;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire _10872_;
 wire _10873_;
 wire _10874_;
 wire _10875_;
 wire _10876_;
 wire _10877_;
 wire _10878_;
 wire _10879_;
 wire net4624;
 wire _10881_;
 wire _10882_;
 wire net4622;
 wire _10884_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire _10889_;
 wire net4621;
 wire _10891_;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire net4619;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire net4620;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire net4623;
 wire _10908_;
 wire net4627;
 wire _10910_;
 wire _10911_;
 wire _10912_;
 wire _10913_;
 wire _10914_;
 wire _10915_;
 wire _10916_;
 wire _10917_;
 wire _10918_;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10923_;
 wire _10924_;
 wire _10926_;
 wire _10927_;
 wire net4618;
 wire _10929_;
 wire _10931_;
 wire _10932_;
 wire _10933_;
 wire _10934_;
 wire _10935_;
 wire _10937_;
 wire _10938_;
 wire _10939_;
 wire _10940_;
 wire _10941_;
 wire _10942_;
 wire _10943_;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire _10947_;
 wire _10948_;
 wire _10949_;
 wire _10950_;
 wire _10951_;
 wire _10952_;
 wire _10953_;
 wire _10954_;
 wire _10955_;
 wire _10956_;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire _10960_;
 wire _10961_;
 wire _10962_;
 wire _10963_;
 wire _10964_;
 wire _10965_;
 wire _10966_;
 wire _10967_;
 wire _10968_;
 wire _10969_;
 wire _10970_;
 wire _10971_;
 wire _10972_;
 wire _10973_;
 wire _10975_;
 wire _10976_;
 wire _10977_;
 wire _10978_;
 wire _10979_;
 wire _10980_;
 wire _10981_;
 wire _10982_;
 wire _10983_;
 wire _10984_;
 wire _10985_;
 wire _10986_;
 wire _10987_;
 wire _10988_;
 wire _10989_;
 wire _10990_;
 wire _10991_;
 wire _10992_;
 wire _10993_;
 wire _10994_;
 wire _10995_;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire _10999_;
 wire _11000_;
 wire _11001_;
 wire _11002_;
 wire _11003_;
 wire _11004_;
 wire _11005_;
 wire _11006_;
 wire _11007_;
 wire _11008_;
 wire _11009_;
 wire _11010_;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire _11015_;
 wire _11016_;
 wire _11017_;
 wire _11018_;
 wire _11019_;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire _11025_;
 wire _11026_;
 wire _11027_;
 wire _11028_;
 wire _11029_;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire _11034_;
 wire _11035_;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire _11043_;
 wire _11044_;
 wire _11045_;
 wire _11046_;
 wire _11047_;
 wire _11048_;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11052_;
 wire _11053_;
 wire _11054_;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire _11058_;
 wire _11059_;
 wire _11060_;
 wire _11061_;
 wire _11062_;
 wire _11063_;
 wire _11064_;
 wire _11065_;
 wire _11066_;
 wire _11067_;
 wire _11068_;
 wire _11069_;
 wire _11070_;
 wire _11071_;
 wire _11072_;
 wire _11073_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire _11077_;
 wire _11078_;
 wire _11079_;
 wire _11080_;
 wire _11081_;
 wire _11082_;
 wire _11083_;
 wire _11084_;
 wire _11085_;
 wire _11086_;
 wire _11087_;
 wire _11088_;
 wire _11089_;
 wire _11090_;
 wire _11091_;
 wire _11092_;
 wire _11093_;
 wire _11094_;
 wire _11095_;
 wire _11096_;
 wire _11097_;
 wire _11098_;
 wire _11099_;
 wire _11100_;
 wire _11101_;
 wire _11102_;
 wire _11103_;
 wire _11104_;
 wire _11105_;
 wire _11106_;
 wire _11107_;
 wire _11108_;
 wire _11109_;
 wire _11110_;
 wire _11111_;
 wire _11112_;
 wire _11113_;
 wire _11114_;
 wire _11115_;
 wire _11116_;
 wire _11117_;
 wire _11118_;
 wire _11119_;
 wire _11120_;
 wire _11121_;
 wire _11122_;
 wire _11123_;
 wire _11124_;
 wire _11125_;
 wire _11126_;
 wire _11127_;
 wire _11128_;
 wire _11129_;
 wire _11130_;
 wire _11131_;
 wire _11132_;
 wire _11133_;
 wire _11134_;
 wire _11135_;
 wire _11136_;
 wire _11137_;
 wire _11138_;
 wire _11139_;
 wire _11140_;
 wire _11141_;
 wire _11142_;
 wire _11143_;
 wire _11144_;
 wire _11145_;
 wire _11146_;
 wire _11147_;
 wire _11148_;
 wire _11149_;
 wire _11150_;
 wire _11151_;
 wire _11152_;
 wire _11153_;
 wire _11154_;
 wire _11155_;
 wire _11156_;
 wire _11157_;
 wire _11158_;
 wire _11159_;
 wire _11160_;
 wire _11161_;
 wire _11162_;
 wire _11163_;
 wire _11164_;
 wire _11165_;
 wire _11166_;
 wire _11167_;
 wire _11168_;
 wire _11169_;
 wire _11170_;
 wire _11171_;
 wire _11172_;
 wire _11173_;
 wire _11174_;
 wire _11175_;
 wire _11176_;
 wire _11177_;
 wire _11178_;
 wire _11179_;
 wire _11180_;
 wire _11181_;
 wire _11182_;
 wire _11183_;
 wire _11184_;
 wire _11185_;
 wire _11186_;
 wire _11187_;
 wire _11188_;
 wire _11189_;
 wire _11190_;
 wire _11191_;
 wire _11192_;
 wire _11193_;
 wire _11194_;
 wire _11195_;
 wire _11196_;
 wire _11197_;
 wire _11198_;
 wire _11199_;
 wire _11200_;
 wire _11201_;
 wire _11202_;
 wire _11203_;
 wire _11204_;
 wire _11205_;
 wire _11206_;
 wire _11207_;
 wire _11208_;
 wire _11209_;
 wire _11210_;
 wire _11211_;
 wire _11212_;
 wire _11213_;
 wire _11214_;
 wire _11215_;
 wire _11216_;
 wire _11217_;
 wire _11218_;
 wire _11219_;
 wire _11220_;
 wire _11221_;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire _11225_;
 wire _11226_;
 wire _11227_;
 wire _11228_;
 wire _11229_;
 wire _11230_;
 wire _11231_;
 wire _11232_;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11237_;
 wire _11238_;
 wire _11239_;
 wire _11240_;
 wire _11241_;
 wire _11242_;
 wire _11243_;
 wire _11244_;
 wire _11245_;
 wire _11246_;
 wire _11247_;
 wire _11248_;
 wire _11249_;
 wire _11250_;
 wire _11251_;
 wire _11252_;
 wire _11253_;
 wire _11254_;
 wire _11255_;
 wire _11256_;
 wire _11257_;
 wire _11258_;
 wire _11259_;
 wire _11260_;
 wire _11261_;
 wire _11262_;
 wire _11263_;
 wire _11264_;
 wire _11265_;
 wire _11266_;
 wire _11267_;
 wire _11268_;
 wire _11269_;
 wire _11270_;
 wire _11271_;
 wire _11272_;
 wire _11273_;
 wire _11274_;
 wire _11275_;
 wire _11276_;
 wire _11277_;
 wire _11278_;
 wire _11279_;
 wire _11280_;
 wire _11281_;
 wire _11282_;
 wire _11283_;
 wire _11284_;
 wire _11285_;
 wire _11286_;
 wire _11287_;
 wire _11288_;
 wire _11289_;
 wire _11290_;
 wire _11291_;
 wire _11292_;
 wire _11293_;
 wire _11294_;
 wire _11295_;
 wire _11296_;
 wire _11297_;
 wire _11298_;
 wire _11299_;
 wire _11300_;
 wire _11301_;
 wire _11302_;
 wire _11303_;
 wire _11304_;
 wire _11305_;
 wire _11306_;
 wire _11307_;
 wire _11308_;
 wire _11309_;
 wire _11310_;
 wire _11311_;
 wire _11312_;
 wire _11313_;
 wire _11314_;
 wire _11315_;
 wire _11316_;
 wire _11317_;
 wire _11318_;
 wire _11319_;
 wire _11320_;
 wire _11321_;
 wire _11322_;
 wire _11323_;
 wire _11324_;
 wire _11325_;
 wire _11326_;
 wire _11327_;
 wire _11328_;
 wire _11329_;
 wire _11330_;
 wire _11331_;
 wire _11332_;
 wire _11333_;
 wire _11334_;
 wire _11335_;
 wire _11336_;
 wire _11337_;
 wire _11338_;
 wire _11339_;
 wire _11340_;
 wire _11341_;
 wire _11342_;
 wire _11343_;
 wire _11344_;
 wire _11345_;
 wire _11346_;
 wire _11347_;
 wire _11348_;
 wire _11349_;
 wire _11350_;
 wire _11351_;
 wire _11352_;
 wire _11353_;
 wire _11354_;
 wire _11355_;
 wire _11356_;
 wire _11357_;
 wire _11358_;
 wire _11359_;
 wire _11360_;
 wire _11361_;
 wire _11362_;
 wire _11363_;
 wire _11364_;
 wire _11365_;
 wire _11366_;
 wire _11367_;
 wire _11368_;
 wire _11369_;
 wire _11370_;
 wire _11371_;
 wire _11372_;
 wire _11373_;
 wire _11374_;
 wire _11375_;
 wire _11376_;
 wire _11377_;
 wire _11378_;
 wire _11379_;
 wire _11380_;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire _11384_;
 wire _11385_;
 wire _11386_;
 wire _11387_;
 wire _11388_;
 wire _11389_;
 wire _11390_;
 wire _11391_;
 wire _11392_;
 wire _11393_;
 wire _11394_;
 wire _11395_;
 wire _11396_;
 wire _11397_;
 wire _11398_;
 wire _11399_;
 wire _11400_;
 wire _11401_;
 wire _11402_;
 wire _11403_;
 wire _11404_;
 wire _11405_;
 wire _11406_;
 wire _11407_;
 wire _11408_;
 wire _11409_;
 wire _11410_;
 wire _11411_;
 wire _11412_;
 wire _11413_;
 wire _11414_;
 wire _11415_;
 wire _11416_;
 wire _11417_;
 wire _11418_;
 wire _11419_;
 wire _11420_;
 wire _11421_;
 wire _11422_;
 wire _11423_;
 wire _11424_;
 wire _11425_;
 wire _11426_;
 wire _11427_;
 wire _11428_;
 wire _11429_;
 wire _11430_;
 wire _11431_;
 wire _11432_;
 wire _11433_;
 wire _11434_;
 wire _11435_;
 wire _11436_;
 wire _11437_;
 wire _11438_;
 wire _11439_;
 wire _11440_;
 wire _11441_;
 wire _11442_;
 wire _11443_;
 wire _11444_;
 wire _11445_;
 wire _11446_;
 wire _11447_;
 wire _11448_;
 wire net4614;
 wire _11450_;
 wire net4613;
 wire _11452_;
 wire net4615;
 wire _11454_;
 wire _11455_;
 wire _11456_;
 wire _11457_;
 wire net4612;
 wire net4610;
 wire net4609;
 wire net4608;
 wire _11462_;
 wire _11463_;
 wire _11464_;
 wire _11465_;
 wire net4607;
 wire _11467_;
 wire _11468_;
 wire _11469_;
 wire _11470_;
 wire _11471_;
 wire _11472_;
 wire _11473_;
 wire _11474_;
 wire _11475_;
 wire _11476_;
 wire _11477_;
 wire net4606;
 wire _11480_;
 wire _11481_;
 wire _11482_;
 wire _11483_;
 wire _11484_;
 wire _11485_;
 wire _11486_;
 wire _11487_;
 wire _11488_;
 wire _11489_;
 wire _11490_;
 wire net4605;
 wire _11493_;
 wire net4604;
 wire _11496_;
 wire _11497_;
 wire _11498_;
 wire _11499_;
 wire _11501_;
 wire _11502_;
 wire _11503_;
 wire _11504_;
 wire _11505_;
 wire _11506_;
 wire _11507_;
 wire _11508_;
 wire _11509_;
 wire _11510_;
 wire net4602;
 wire net4603;
 wire _11513_;
 wire _11514_;
 wire _11515_;
 wire _11516_;
 wire _11517_;
 wire _11518_;
 wire _11519_;
 wire net4601;
 wire net4600;
 wire _11522_;
 wire _11523_;
 wire net4599;
 wire net4597;
 wire net4598;
 wire _11527_;
 wire _11528_;
 wire net4596;
 wire _11530_;
 wire _11531_;
 wire net4594;
 wire _11533_;
 wire _11534_;
 wire _11535_;
 wire _11536_;
 wire _11537_;
 wire net4593;
 wire net4592;
 wire _11540_;
 wire _11541_;
 wire _11542_;
 wire _11543_;
 wire net4595;
 wire _11546_;
 wire _11547_;
 wire net4590;
 wire _11549_;
 wire _11550_;
 wire _11551_;
 wire _11552_;
 wire _11553_;
 wire _11554_;
 wire net4589;
 wire _11556_;
 wire _11557_;
 wire _11558_;
 wire _11559_;
 wire _11561_;
 wire _11562_;
 wire _11563_;
 wire _11564_;
 wire _11565_;
 wire _11566_;
 wire _11567_;
 wire _11568_;
 wire _11569_;
 wire _11570_;
 wire _11571_;
 wire _11572_;
 wire _11573_;
 wire _11574_;
 wire _11575_;
 wire _11576_;
 wire net4588;
 wire _11578_;
 wire _11579_;
 wire _11580_;
 wire _11581_;
 wire _11582_;
 wire _11583_;
 wire _11584_;
 wire _11585_;
 wire _11586_;
 wire _11587_;
 wire _11588_;
 wire _11589_;
 wire _11590_;
 wire _11591_;
 wire _11592_;
 wire _11593_;
 wire _11594_;
 wire _11595_;
 wire _11596_;
 wire _11597_;
 wire _11598_;
 wire _11599_;
 wire _11600_;
 wire net4586;
 wire _11602_;
 wire _11603_;
 wire _11604_;
 wire _11605_;
 wire _11606_;
 wire net4587;
 wire _11608_;
 wire _11609_;
 wire _11610_;
 wire _11611_;
 wire net4585;
 wire net4584;
 wire _11614_;
 wire net4583;
 wire _11617_;
 wire _11618_;
 wire _11619_;
 wire _11620_;
 wire _11621_;
 wire _11622_;
 wire _11623_;
 wire _11624_;
 wire _11625_;
 wire _11627_;
 wire _11628_;
 wire _11629_;
 wire _11630_;
 wire _11631_;
 wire net4582;
 wire _11633_;
 wire _11634_;
 wire _11635_;
 wire _11636_;
 wire _11637_;
 wire _11638_;
 wire _11639_;
 wire _11640_;
 wire _11641_;
 wire _11642_;
 wire net4581;
 wire _11644_;
 wire _11645_;
 wire net4579;
 wire _11647_;
 wire _11648_;
 wire _11649_;
 wire _11650_;
 wire _11651_;
 wire _11652_;
 wire _11653_;
 wire _11654_;
 wire net4578;
 wire _11656_;
 wire _11657_;
 wire _11658_;
 wire _11659_;
 wire _11660_;
 wire _11661_;
 wire net4577;
 wire _11663_;
 wire _11664_;
 wire _11665_;
 wire _11666_;
 wire _11667_;
 wire _11668_;
 wire _11669_;
 wire _11670_;
 wire _11671_;
 wire _11672_;
 wire _11673_;
 wire _11674_;
 wire _11675_;
 wire _11676_;
 wire _11677_;
 wire _11678_;
 wire _11679_;
 wire _11680_;
 wire _11681_;
 wire _11682_;
 wire _11683_;
 wire _11684_;
 wire _11685_;
 wire _11686_;
 wire _11687_;
 wire _11688_;
 wire _11689_;
 wire _11690_;
 wire _11691_;
 wire _11692_;
 wire _11693_;
 wire _11694_;
 wire _11695_;
 wire _11696_;
 wire _11697_;
 wire _11698_;
 wire _11699_;
 wire _11700_;
 wire _11701_;
 wire _11702_;
 wire _11703_;
 wire _11704_;
 wire _11705_;
 wire _11706_;
 wire _11707_;
 wire _11708_;
 wire _11709_;
 wire _11710_;
 wire _11711_;
 wire _11712_;
 wire _11713_;
 wire _11714_;
 wire _11715_;
 wire _11716_;
 wire _11717_;
 wire _11718_;
 wire _11719_;
 wire _11720_;
 wire _11721_;
 wire _11722_;
 wire _11723_;
 wire _11724_;
 wire _11725_;
 wire _11726_;
 wire _11727_;
 wire _11728_;
 wire _11729_;
 wire _11730_;
 wire _11731_;
 wire _11732_;
 wire _11733_;
 wire _11734_;
 wire _11735_;
 wire _11736_;
 wire _11737_;
 wire _11738_;
 wire _11739_;
 wire _11740_;
 wire _11741_;
 wire _11742_;
 wire _11743_;
 wire _11744_;
 wire _11745_;
 wire _11746_;
 wire _11747_;
 wire _11748_;
 wire _11749_;
 wire _11750_;
 wire _11751_;
 wire _11752_;
 wire _11753_;
 wire _11754_;
 wire _11755_;
 wire _11756_;
 wire _11757_;
 wire _11758_;
 wire _11759_;
 wire _11760_;
 wire _11761_;
 wire _11762_;
 wire _11763_;
 wire _11764_;
 wire _11765_;
 wire _11766_;
 wire _11767_;
 wire _11768_;
 wire _11769_;
 wire _11770_;
 wire _11771_;
 wire _11772_;
 wire _11773_;
 wire _11774_;
 wire _11775_;
 wire _11776_;
 wire _11777_;
 wire _11778_;
 wire _11779_;
 wire _11780_;
 wire _11781_;
 wire _11782_;
 wire _11783_;
 wire _11784_;
 wire _11785_;
 wire _11786_;
 wire _11787_;
 wire _11788_;
 wire _11789_;
 wire _11790_;
 wire _11791_;
 wire _11792_;
 wire _11793_;
 wire _11794_;
 wire _11795_;
 wire _11796_;
 wire _11797_;
 wire _11798_;
 wire _11799_;
 wire _11800_;
 wire _11801_;
 wire _11802_;
 wire _11803_;
 wire _11804_;
 wire _11805_;
 wire _11806_;
 wire _11807_;
 wire _11808_;
 wire _11809_;
 wire _11810_;
 wire _11811_;
 wire _11812_;
 wire _11813_;
 wire _11814_;
 wire _11815_;
 wire _11816_;
 wire _11817_;
 wire _11818_;
 wire _11819_;
 wire _11820_;
 wire _11821_;
 wire _11822_;
 wire _11823_;
 wire _11824_;
 wire _11825_;
 wire _11826_;
 wire _11827_;
 wire _11828_;
 wire _11829_;
 wire _11830_;
 wire _11831_;
 wire _11832_;
 wire _11833_;
 wire _11834_;
 wire _11835_;
 wire _11836_;
 wire _11837_;
 wire _11838_;
 wire _11839_;
 wire _11840_;
 wire _11841_;
 wire _11842_;
 wire _11843_;
 wire _11844_;
 wire _11845_;
 wire _11846_;
 wire _11847_;
 wire _11848_;
 wire _11849_;
 wire _11850_;
 wire _11851_;
 wire _11852_;
 wire _11853_;
 wire _11854_;
 wire _11855_;
 wire _11856_;
 wire _11857_;
 wire _11858_;
 wire _11859_;
 wire _11860_;
 wire _11861_;
 wire _11862_;
 wire _11863_;
 wire _11864_;
 wire _11865_;
 wire _11866_;
 wire _11867_;
 wire _11868_;
 wire _11869_;
 wire _11870_;
 wire _11871_;
 wire _11872_;
 wire _11873_;
 wire _11874_;
 wire _11875_;
 wire _11876_;
 wire _11877_;
 wire _11878_;
 wire _11879_;
 wire _11880_;
 wire _11881_;
 wire _11882_;
 wire _11883_;
 wire _11884_;
 wire _11885_;
 wire _11886_;
 wire _11887_;
 wire _11888_;
 wire _11889_;
 wire _11890_;
 wire _11891_;
 wire _11892_;
 wire _11893_;
 wire _11894_;
 wire _11895_;
 wire _11896_;
 wire _11897_;
 wire _11898_;
 wire _11899_;
 wire _11900_;
 wire _11901_;
 wire _11902_;
 wire _11903_;
 wire _11904_;
 wire _11905_;
 wire _11906_;
 wire _11907_;
 wire _11908_;
 wire _11909_;
 wire _11910_;
 wire _11911_;
 wire _11912_;
 wire _11913_;
 wire _11914_;
 wire _11915_;
 wire _11916_;
 wire _11917_;
 wire _11918_;
 wire _11919_;
 wire _11920_;
 wire _11921_;
 wire _11922_;
 wire _11923_;
 wire _11924_;
 wire _11925_;
 wire _11926_;
 wire _11927_;
 wire _11928_;
 wire _11929_;
 wire _11930_;
 wire _11931_;
 wire _11932_;
 wire _11933_;
 wire _11934_;
 wire _11935_;
 wire _11936_;
 wire _11937_;
 wire _11938_;
 wire _11939_;
 wire _11940_;
 wire _11941_;
 wire _11942_;
 wire _11943_;
 wire _11944_;
 wire _11945_;
 wire _11946_;
 wire _11947_;
 wire _11948_;
 wire _11949_;
 wire _11950_;
 wire _11951_;
 wire _11952_;
 wire _11953_;
 wire _11954_;
 wire _11955_;
 wire _11956_;
 wire _11957_;
 wire _11958_;
 wire _11959_;
 wire _11960_;
 wire _11961_;
 wire _11962_;
 wire _11963_;
 wire _11964_;
 wire _11965_;
 wire _11966_;
 wire _11967_;
 wire _11968_;
 wire _11969_;
 wire _11970_;
 wire _11971_;
 wire _11972_;
 wire _11973_;
 wire _11974_;
 wire _11975_;
 wire _11976_;
 wire _11977_;
 wire _11978_;
 wire _11979_;
 wire _11980_;
 wire _11981_;
 wire _11982_;
 wire _11983_;
 wire _11984_;
 wire _11985_;
 wire _11986_;
 wire _11987_;
 wire _11988_;
 wire _11989_;
 wire _11990_;
 wire _11991_;
 wire _11992_;
 wire _11993_;
 wire _11994_;
 wire _11995_;
 wire _11996_;
 wire _11997_;
 wire _11998_;
 wire _11999_;
 wire _12000_;
 wire _12001_;
 wire _12002_;
 wire _12003_;
 wire _12004_;
 wire _12005_;
 wire _12006_;
 wire _12007_;
 wire _12008_;
 wire _12009_;
 wire _12010_;
 wire _12011_;
 wire _12012_;
 wire _12013_;
 wire _12014_;
 wire _12015_;
 wire _12016_;
 wire _12017_;
 wire _12018_;
 wire _12019_;
 wire _12020_;
 wire _12021_;
 wire _12022_;
 wire _12023_;
 wire _12024_;
 wire _12025_;
 wire _12026_;
 wire _12027_;
 wire _12028_;
 wire _12029_;
 wire _12030_;
 wire _12031_;
 wire _12032_;
 wire _12033_;
 wire _12034_;
 wire _12035_;
 wire _12036_;
 wire _12037_;
 wire _12038_;
 wire _12039_;
 wire _12040_;
 wire _12041_;
 wire _12042_;
 wire _12043_;
 wire _12044_;
 wire _12045_;
 wire _12046_;
 wire _12047_;
 wire _12048_;
 wire _12049_;
 wire _12050_;
 wire _12051_;
 wire _12052_;
 wire _12053_;
 wire _12054_;
 wire _12055_;
 wire _12056_;
 wire _12057_;
 wire _12058_;
 wire _12059_;
 wire _12060_;
 wire _12061_;
 wire _12062_;
 wire _12063_;
 wire _12064_;
 wire _12065_;
 wire _12066_;
 wire _12067_;
 wire _12068_;
 wire _12069_;
 wire _12070_;
 wire _12071_;
 wire _12072_;
 wire _12073_;
 wire _12074_;
 wire _12075_;
 wire _12076_;
 wire _12077_;
 wire _12078_;
 wire _12079_;
 wire _12080_;
 wire _12081_;
 wire _12082_;
 wire _12083_;
 wire _12084_;
 wire _12085_;
 wire _12086_;
 wire _12087_;
 wire _12088_;
 wire _12089_;
 wire _12090_;
 wire _12091_;
 wire _12092_;
 wire _12093_;
 wire _12094_;
 wire _12095_;
 wire _12096_;
 wire _12097_;
 wire _12098_;
 wire _12099_;
 wire _12100_;
 wire _12101_;
 wire _12102_;
 wire _12103_;
 wire _12104_;
 wire _12105_;
 wire _12106_;
 wire _12107_;
 wire _12108_;
 wire _12109_;
 wire _12110_;
 wire _12111_;
 wire _12112_;
 wire _12113_;
 wire _12114_;
 wire _12115_;
 wire _12116_;
 wire _12117_;
 wire _12118_;
 wire _12119_;
 wire _12120_;
 wire _12121_;
 wire _12122_;
 wire _12123_;
 wire _12124_;
 wire _12125_;
 wire _12126_;
 wire _12127_;
 wire _12128_;
 wire _12129_;
 wire _12130_;
 wire _12131_;
 wire _12132_;
 wire _12133_;
 wire _12134_;
 wire _12135_;
 wire _12136_;
 wire _12137_;
 wire _12138_;
 wire _12139_;
 wire _12140_;
 wire _12141_;
 wire _12142_;
 wire _12143_;
 wire _12144_;
 wire _12145_;
 wire _12146_;
 wire _12147_;
 wire _12148_;
 wire _12149_;
 wire _12150_;
 wire net4576;
 wire _12152_;
 wire net4575;
 wire _12154_;
 wire _12155_;
 wire _12156_;
 wire _12157_;
 wire _12158_;
 wire _12159_;
 wire _12160_;
 wire _12161_;
 wire _12162_;
 wire _12163_;
 wire _12164_;
 wire _12165_;
 wire _12166_;
 wire _12167_;
 wire _12168_;
 wire _12169_;
 wire _12170_;
 wire _12171_;
 wire _12172_;
 wire _12173_;
 wire _12174_;
 wire net4574;
 wire _12176_;
 wire _12177_;
 wire _12178_;
 wire _12179_;
 wire _12180_;
 wire _12181_;
 wire _12182_;
 wire net4567;
 wire net4566;
 wire _12185_;
 wire net4568;
 wire _12187_;
 wire _12188_;
 wire _12189_;
 wire _12190_;
 wire _12191_;
 wire _12192_;
 wire _12193_;
 wire _12194_;
 wire _12195_;
 wire _12196_;
 wire _12197_;
 wire _12198_;
 wire _12199_;
 wire _12200_;
 wire _12201_;
 wire net4572;
 wire net4570;
 wire _12204_;
 wire _12205_;
 wire _12206_;
 wire _12207_;
 wire _12208_;
 wire net4563;
 wire net4562;
 wire _12211_;
 wire _12212_;
 wire _12213_;
 wire _12214_;
 wire _12215_;
 wire _12216_;
 wire _12217_;
 wire _12218_;
 wire _12219_;
 wire _12220_;
 wire net4559;
 wire net4558;
 wire _12223_;
 wire _12224_;
 wire _12225_;
 wire _12226_;
 wire net4557;
 wire _12228_;
 wire _12229_;
 wire _12230_;
 wire net4556;
 wire _12232_;
 wire net4554;
 wire _12234_;
 wire _12235_;
 wire _12236_;
 wire _12237_;
 wire _12238_;
 wire _12239_;
 wire net4555;
 wire net4552;
 wire _12242_;
 wire _12243_;
 wire _12244_;
 wire _12245_;
 wire net4551;
 wire _12247_;
 wire _12248_;
 wire net4550;
 wire _12250_;
 wire _12251_;
 wire _12252_;
 wire _12253_;
 wire net4549;
 wire _12255_;
 wire _12256_;
 wire net4548;
 wire _12258_;
 wire _12259_;
 wire net4547;
 wire net4560;
 wire _12262_;
 wire _12263_;
 wire _12264_;
 wire _12265_;
 wire _12266_;
 wire net4553;
 wire net4546;
 wire _12269_;
 wire _12270_;
 wire _12271_;
 wire _12272_;
 wire _12273_;
 wire _12274_;
 wire _12275_;
 wire _12276_;
 wire _12277_;
 wire net4544;
 wire _12279_;
 wire net4545;
 wire _12281_;
 wire _12282_;
 wire net4543;
 wire net4564;
 wire _12285_;
 wire _12286_;
 wire _12287_;
 wire net4561;
 wire _12289_;
 wire _12290_;
 wire _12291_;
 wire _12292_;
 wire _12293_;
 wire _12294_;
 wire _12295_;
 wire _12296_;
 wire _12297_;
 wire _12298_;
 wire _12299_;
 wire _12300_;
 wire net4539;
 wire net4538;
 wire _12303_;
 wire _12304_;
 wire _12305_;
 wire _12306_;
 wire _12307_;
 wire _12308_;
 wire _12309_;
 wire _12310_;
 wire _12311_;
 wire _12312_;
 wire _12313_;
 wire _12314_;
 wire _12315_;
 wire _12316_;
 wire _12317_;
 wire _12318_;
 wire _12319_;
 wire _12320_;
 wire _12321_;
 wire _12322_;
 wire net4541;
 wire _12324_;
 wire _12325_;
 wire _12326_;
 wire net4537;
 wire _12328_;
 wire _12329_;
 wire _12330_;
 wire _12331_;
 wire _12332_;
 wire net4540;
 wire _12334_;
 wire _12335_;
 wire _12336_;
 wire _12337_;
 wire _12338_;
 wire net4536;
 wire _12340_;
 wire _12341_;
 wire _12342_;
 wire _12343_;
 wire _12344_;
 wire _12345_;
 wire _12346_;
 wire _12347_;
 wire _12348_;
 wire _12349_;
 wire _12350_;
 wire _12351_;
 wire _12352_;
 wire _12353_;
 wire net4535;
 wire _12355_;
 wire _12356_;
 wire _12357_;
 wire _12358_;
 wire _12359_;
 wire _12360_;
 wire _12361_;
 wire _12362_;
 wire _12363_;
 wire _12364_;
 wire _12365_;
 wire _12366_;
 wire net4532;
 wire _12368_;
 wire _12369_;
 wire _12370_;
 wire _12371_;
 wire _12372_;
 wire net4531;
 wire _12374_;
 wire _12375_;
 wire _12376_;
 wire _12377_;
 wire _12378_;
 wire _12379_;
 wire _12380_;
 wire _12381_;
 wire _12382_;
 wire net4530;
 wire _12384_;
 wire _12385_;
 wire _12386_;
 wire _12387_;
 wire _12388_;
 wire _12389_;
 wire _12390_;
 wire _12391_;
 wire _12392_;
 wire net4529;
 wire _12394_;
 wire _12395_;
 wire net4528;
 wire _12397_;
 wire net4527;
 wire _12399_;
 wire _12400_;
 wire _12401_;
 wire _12402_;
 wire _12403_;
 wire _12404_;
 wire _12405_;
 wire _12406_;
 wire _12407_;
 wire _12408_;
 wire _12409_;
 wire _12410_;
 wire _12411_;
 wire _12412_;
 wire _12413_;
 wire _12414_;
 wire _12415_;
 wire _12416_;
 wire _12417_;
 wire _12418_;
 wire _12419_;
 wire _12420_;
 wire _12421_;
 wire _12422_;
 wire _12423_;
 wire _12424_;
 wire _12425_;
 wire _12426_;
 wire _12427_;
 wire _12428_;
 wire _12429_;
 wire _12430_;
 wire _12431_;
 wire _12432_;
 wire _12433_;
 wire _12434_;
 wire _12435_;
 wire _12436_;
 wire _12437_;
 wire net4526;
 wire _12439_;
 wire _12440_;
 wire _12441_;
 wire _12442_;
 wire net4525;
 wire _12444_;
 wire _12445_;
 wire _12446_;
 wire _12447_;
 wire _12448_;
 wire _12449_;
 wire _12450_;
 wire _12451_;
 wire _12452_;
 wire net4533;
 wire _12454_;
 wire _12455_;
 wire _12456_;
 wire _12457_;
 wire _12458_;
 wire _12459_;
 wire _12460_;
 wire _12461_;
 wire _12462_;
 wire _12463_;
 wire _12464_;
 wire _12465_;
 wire _12466_;
 wire _12467_;
 wire _12468_;
 wire _12469_;
 wire _12470_;
 wire _12471_;
 wire _12472_;
 wire _12473_;
 wire _12474_;
 wire _12475_;
 wire _12476_;
 wire _12477_;
 wire _12478_;
 wire _12479_;
 wire _12480_;
 wire _12481_;
 wire _12482_;
 wire _12483_;
 wire _12484_;
 wire _12485_;
 wire _12486_;
 wire _12487_;
 wire _12488_;
 wire _12489_;
 wire _12490_;
 wire _12491_;
 wire _12492_;
 wire _12493_;
 wire _12494_;
 wire _12495_;
 wire _12496_;
 wire _12497_;
 wire _12498_;
 wire _12499_;
 wire _12500_;
 wire _12501_;
 wire _12502_;
 wire _12503_;
 wire net4524;
 wire _12505_;
 wire _12506_;
 wire _12507_;
 wire _12508_;
 wire _12509_;
 wire _12510_;
 wire _12511_;
 wire _12512_;
 wire _12513_;
 wire _12514_;
 wire _12515_;
 wire _12516_;
 wire _12517_;
 wire _12518_;
 wire _12519_;
 wire _12520_;
 wire _12521_;
 wire _12522_;
 wire _12523_;
 wire _12524_;
 wire _12525_;
 wire _12526_;
 wire _12527_;
 wire _12528_;
 wire _12529_;
 wire _12530_;
 wire _12531_;
 wire _12532_;
 wire _12533_;
 wire _12534_;
 wire _12535_;
 wire _12536_;
 wire _12537_;
 wire _12538_;
 wire net4523;
 wire _12540_;
 wire _12541_;
 wire _12542_;
 wire _12543_;
 wire _12544_;
 wire _12545_;
 wire _12546_;
 wire _12547_;
 wire _12548_;
 wire _12549_;
 wire _12550_;
 wire _12551_;
 wire _12552_;
 wire _12553_;
 wire _12554_;
 wire _12555_;
 wire _12556_;
 wire _12557_;
 wire _12558_;
 wire _12559_;
 wire _12560_;
 wire _12561_;
 wire _12562_;
 wire _12563_;
 wire _12564_;
 wire _12565_;
 wire _12566_;
 wire _12567_;
 wire _12568_;
 wire _12569_;
 wire _12570_;
 wire _12571_;
 wire _12572_;
 wire _12573_;
 wire _12574_;
 wire _12575_;
 wire _12576_;
 wire _12577_;
 wire _12578_;
 wire _12579_;
 wire _12580_;
 wire _12581_;
 wire _12582_;
 wire _12583_;
 wire _12584_;
 wire _12585_;
 wire _12586_;
 wire _12587_;
 wire _12588_;
 wire _12589_;
 wire _12590_;
 wire _12591_;
 wire _12592_;
 wire _12593_;
 wire _12594_;
 wire _12595_;
 wire _12596_;
 wire _12597_;
 wire _12598_;
 wire _12599_;
 wire _12600_;
 wire _12601_;
 wire _12602_;
 wire _12603_;
 wire _12604_;
 wire _12605_;
 wire _12606_;
 wire _12607_;
 wire _12608_;
 wire _12609_;
 wire _12610_;
 wire _12611_;
 wire _12612_;
 wire _12613_;
 wire _12614_;
 wire _12615_;
 wire _12616_;
 wire _12617_;
 wire _12618_;
 wire _12619_;
 wire _12620_;
 wire _12621_;
 wire _12622_;
 wire _12623_;
 wire _12624_;
 wire _12625_;
 wire _12626_;
 wire _12627_;
 wire _12628_;
 wire _12629_;
 wire _12630_;
 wire _12631_;
 wire _12632_;
 wire _12633_;
 wire _12634_;
 wire _12635_;
 wire _12636_;
 wire _12637_;
 wire _12638_;
 wire _12639_;
 wire _12640_;
 wire _12641_;
 wire _12642_;
 wire _12643_;
 wire _12644_;
 wire _12645_;
 wire _12646_;
 wire _12647_;
 wire _12648_;
 wire _12649_;
 wire _12650_;
 wire _12651_;
 wire _12652_;
 wire _12653_;
 wire _12654_;
 wire _12655_;
 wire _12656_;
 wire _12657_;
 wire _12658_;
 wire _12659_;
 wire _12660_;
 wire _12661_;
 wire _12662_;
 wire _12663_;
 wire _12664_;
 wire _12665_;
 wire _12666_;
 wire _12667_;
 wire _12668_;
 wire _12669_;
 wire _12670_;
 wire _12671_;
 wire _12672_;
 wire _12673_;
 wire _12674_;
 wire _12675_;
 wire _12676_;
 wire _12677_;
 wire _12678_;
 wire _12679_;
 wire _12680_;
 wire _12681_;
 wire _12682_;
 wire _12683_;
 wire _12684_;
 wire _12685_;
 wire _12686_;
 wire _12687_;
 wire _12688_;
 wire _12689_;
 wire _12690_;
 wire _12691_;
 wire _12692_;
 wire _12693_;
 wire _12694_;
 wire _12695_;
 wire _12696_;
 wire _12697_;
 wire _12698_;
 wire _12699_;
 wire _12700_;
 wire _12701_;
 wire _12702_;
 wire _12703_;
 wire _12704_;
 wire _12705_;
 wire _12706_;
 wire _12707_;
 wire _12708_;
 wire _12709_;
 wire _12710_;
 wire _12711_;
 wire _12712_;
 wire _12713_;
 wire _12714_;
 wire _12715_;
 wire _12716_;
 wire _12717_;
 wire _12718_;
 wire _12719_;
 wire _12720_;
 wire _12721_;
 wire _12722_;
 wire _12723_;
 wire _12724_;
 wire _12725_;
 wire _12726_;
 wire _12727_;
 wire _12728_;
 wire _12729_;
 wire _12730_;
 wire _12731_;
 wire _12732_;
 wire _12733_;
 wire _12734_;
 wire _12735_;
 wire _12736_;
 wire _12737_;
 wire _12738_;
 wire _12739_;
 wire _12740_;
 wire _12741_;
 wire _12742_;
 wire _12743_;
 wire _12744_;
 wire _12745_;
 wire _12746_;
 wire _12747_;
 wire _12748_;
 wire _12749_;
 wire _12750_;
 wire _12751_;
 wire _12752_;
 wire _12753_;
 wire _12754_;
 wire _12755_;
 wire _12756_;
 wire _12757_;
 wire _12758_;
 wire _12759_;
 wire _12760_;
 wire _12761_;
 wire _12762_;
 wire _12763_;
 wire _12764_;
 wire _12765_;
 wire _12766_;
 wire _12767_;
 wire _12768_;
 wire _12769_;
 wire _12770_;
 wire _12771_;
 wire _12772_;
 wire _12773_;
 wire _12774_;
 wire _12775_;
 wire _12776_;
 wire _12777_;
 wire _12778_;
 wire _12779_;
 wire _12780_;
 wire _12781_;
 wire _12782_;
 wire _12783_;
 wire _12784_;
 wire _12785_;
 wire _12786_;
 wire _12787_;
 wire _12788_;
 wire _12789_;
 wire _12790_;
 wire _12791_;
 wire _12792_;
 wire _12793_;
 wire _12794_;
 wire _12795_;
 wire _12796_;
 wire _12797_;
 wire _12798_;
 wire _12799_;
 wire _12800_;
 wire _12801_;
 wire _12802_;
 wire _12803_;
 wire _12804_;
 wire _12805_;
 wire _12806_;
 wire _12807_;
 wire _12808_;
 wire _12809_;
 wire _12810_;
 wire _12811_;
 wire _12812_;
 wire _12813_;
 wire _12814_;
 wire _12815_;
 wire _12816_;
 wire _12817_;
 wire _12818_;
 wire _12819_;
 wire _12820_;
 wire _12821_;
 wire _12822_;
 wire _12823_;
 wire _12824_;
 wire net4534;
 wire _12826_;
 wire _12827_;
 wire _12828_;
 wire _12829_;
 wire _12830_;
 wire _12831_;
 wire _12832_;
 wire _12833_;
 wire _12834_;
 wire _12835_;
 wire _12836_;
 wire _12837_;
 wire _12838_;
 wire _12839_;
 wire _12840_;
 wire _12841_;
 wire _12842_;
 wire _12843_;
 wire _12844_;
 wire _12845_;
 wire _12846_;
 wire _12847_;
 wire _12848_;
 wire _12849_;
 wire _12850_;
 wire _12851_;
 wire _12852_;
 wire _12853_;
 wire _12854_;
 wire _12855_;
 wire _12856_;
 wire _12857_;
 wire _12858_;
 wire _12859_;
 wire _12860_;
 wire _12861_;
 wire _12862_;
 wire _12863_;
 wire _12864_;
 wire _12865_;
 wire _12866_;
 wire net4519;
 wire _12868_;
 wire _12869_;
 wire _12870_;
 wire _12871_;
 wire _12872_;
 wire _12873_;
 wire _12874_;
 wire net4516;
 wire net4515;
 wire net4513;
 wire _12878_;
 wire _12879_;
 wire net4542;
 wire _12881_;
 wire _12882_;
 wire _12883_;
 wire _12884_;
 wire _12885_;
 wire _12886_;
 wire _12887_;
 wire _12888_;
 wire _12889_;
 wire _12890_;
 wire _12891_;
 wire _12892_;
 wire _12893_;
 wire _12894_;
 wire net4512;
 wire net4514;
 wire _12897_;
 wire net4509;
 wire net4508;
 wire net4507;
 wire net4506;
 wire net4510;
 wire _12903_;
 wire _12904_;
 wire _12905_;
 wire _12906_;
 wire _12907_;
 wire _12908_;
 wire _12909_;
 wire _12910_;
 wire _12911_;
 wire _12912_;
 wire _12913_;
 wire _12914_;
 wire _12915_;
 wire _12916_;
 wire net4511;
 wire net4505;
 wire _12919_;
 wire _12920_;
 wire _12921_;
 wire net4565;
 wire _12923_;
 wire _12924_;
 wire _12925_;
 wire _12927_;
 wire _12928_;
 wire _12929_;
 wire _12930_;
 wire _12931_;
 wire _12932_;
 wire _12933_;
 wire _12934_;
 wire _12935_;
 wire _12936_;
 wire _12937_;
 wire _12938_;
 wire _12939_;
 wire net4504;
 wire _12942_;
 wire _12943_;
 wire _12944_;
 wire _12945_;
 wire net4502;
 wire _12947_;
 wire _12948_;
 wire net4501;
 wire _12950_;
 wire _12951_;
 wire net4500;
 wire _12953_;
 wire _12954_;
 wire _12955_;
 wire _12956_;
 wire _12957_;
 wire _12958_;
 wire _12959_;
 wire _12960_;
 wire _12961_;
 wire net4503;
 wire _12963_;
 wire _12964_;
 wire _12965_;
 wire _12966_;
 wire net4499;
 wire _12969_;
 wire _12970_;
 wire _12971_;
 wire net4498;
 wire _12973_;
 wire _12974_;
 wire net4497;
 wire _12976_;
 wire _12977_;
 wire _12978_;
 wire _12979_;
 wire _12980_;
 wire _12981_;
 wire _12983_;
 wire _12985_;
 wire _12986_;
 wire _12987_;
 wire _12988_;
 wire _12989_;
 wire _12990_;
 wire _12991_;
 wire _12992_;
 wire _12993_;
 wire _12994_;
 wire net4496;
 wire _12996_;
 wire _12997_;
 wire _12999_;
 wire _13000_;
 wire _13001_;
 wire net4495;
 wire _13003_;
 wire _13004_;
 wire _13005_;
 wire _13006_;
 wire _13007_;
 wire _13008_;
 wire _13009_;
 wire _13010_;
 wire _13011_;
 wire _13012_;
 wire _13013_;
 wire _13014_;
 wire _13015_;
 wire _13016_;
 wire net4494;
 wire _13018_;
 wire _13019_;
 wire _13020_;
 wire _13021_;
 wire _13022_;
 wire _13023_;
 wire _13024_;
 wire _13025_;
 wire _13026_;
 wire _13027_;
 wire _13028_;
 wire _13029_;
 wire _13030_;
 wire _13031_;
 wire _13032_;
 wire _13033_;
 wire _13034_;
 wire _13035_;
 wire _13036_;
 wire _13037_;
 wire net4493;
 wire _13039_;
 wire _13040_;
 wire _13041_;
 wire _13042_;
 wire _13043_;
 wire _13044_;
 wire _13045_;
 wire _13046_;
 wire net4492;
 wire _13048_;
 wire _13050_;
 wire _13051_;
 wire _13052_;
 wire _13053_;
 wire _13054_;
 wire _13055_;
 wire _13056_;
 wire _13057_;
 wire _13058_;
 wire _13060_;
 wire _13061_;
 wire _13062_;
 wire _13063_;
 wire _13064_;
 wire _13065_;
 wire _13066_;
 wire _13068_;
 wire _13069_;
 wire _13070_;
 wire _13071_;
 wire _13072_;
 wire _13073_;
 wire _13074_;
 wire _13075_;
 wire _13076_;
 wire _13077_;
 wire _13078_;
 wire _13079_;
 wire _13080_;
 wire net4491;
 wire _13082_;
 wire net4487;
 wire _13084_;
 wire _13085_;
 wire _13086_;
 wire _13087_;
 wire _13088_;
 wire _13089_;
 wire _13090_;
 wire _13091_;
 wire _13092_;
 wire _13093_;
 wire _13094_;
 wire _13095_;
 wire net4488;
 wire _13097_;
 wire net4486;
 wire _13099_;
 wire _13100_;
 wire _13101_;
 wire _13102_;
 wire _13103_;
 wire net4484;
 wire _13105_;
 wire _13106_;
 wire net4485;
 wire _13108_;
 wire _13109_;
 wire _13110_;
 wire _13111_;
 wire _13112_;
 wire _13113_;
 wire _13114_;
 wire _13115_;
 wire _13116_;
 wire net4489;
 wire _13118_;
 wire _13119_;
 wire _13120_;
 wire net4490;
 wire _13122_;
 wire _13123_;
 wire _13124_;
 wire _13125_;
 wire _13126_;
 wire _13127_;
 wire _13128_;
 wire _13129_;
 wire _13130_;
 wire _13131_;
 wire _13132_;
 wire _13133_;
 wire _13134_;
 wire _13135_;
 wire _13136_;
 wire _13137_;
 wire _13138_;
 wire _13139_;
 wire _13140_;
 wire _13141_;
 wire _13142_;
 wire _13143_;
 wire _13144_;
 wire _13145_;
 wire _13146_;
 wire _13147_;
 wire _13148_;
 wire _13149_;
 wire _13150_;
 wire _13151_;
 wire _13152_;
 wire _13153_;
 wire _13154_;
 wire _13155_;
 wire _13156_;
 wire _13157_;
 wire _13158_;
 wire _13159_;
 wire _13160_;
 wire _13161_;
 wire _13162_;
 wire _13163_;
 wire _13164_;
 wire _13165_;
 wire _13166_;
 wire _13167_;
 wire _13168_;
 wire _13169_;
 wire _13170_;
 wire _13171_;
 wire _13172_;
 wire _13173_;
 wire _13174_;
 wire _13175_;
 wire _13176_;
 wire _13177_;
 wire _13178_;
 wire _13179_;
 wire _13180_;
 wire _13181_;
 wire net4483;
 wire _13183_;
 wire _13184_;
 wire _13185_;
 wire _13186_;
 wire _13187_;
 wire _13188_;
 wire _13189_;
 wire _13190_;
 wire _13191_;
 wire _13192_;
 wire _13193_;
 wire _13194_;
 wire _13195_;
 wire _13196_;
 wire _13197_;
 wire _13198_;
 wire _13199_;
 wire _13200_;
 wire _13201_;
 wire _13202_;
 wire _13203_;
 wire _13204_;
 wire _13205_;
 wire _13206_;
 wire _13207_;
 wire _13208_;
 wire _13210_;
 wire _13211_;
 wire _13212_;
 wire _13213_;
 wire _13214_;
 wire _13215_;
 wire _13216_;
 wire _13217_;
 wire _13218_;
 wire _13219_;
 wire _13220_;
 wire _13221_;
 wire _13222_;
 wire _13223_;
 wire _13224_;
 wire _13225_;
 wire _13226_;
 wire _13227_;
 wire _13228_;
 wire _13229_;
 wire _13230_;
 wire _13231_;
 wire _13232_;
 wire _13233_;
 wire _13234_;
 wire _13235_;
 wire _13236_;
 wire _13237_;
 wire _13238_;
 wire _13239_;
 wire _13240_;
 wire _13241_;
 wire _13242_;
 wire _13243_;
 wire _13244_;
 wire _13245_;
 wire _13246_;
 wire _13247_;
 wire _13248_;
 wire _13249_;
 wire _13250_;
 wire _13251_;
 wire _13252_;
 wire _13253_;
 wire _13254_;
 wire _13255_;
 wire _13256_;
 wire _13257_;
 wire _13258_;
 wire _13259_;
 wire _13260_;
 wire _13261_;
 wire _13262_;
 wire _13263_;
 wire _13264_;
 wire _13265_;
 wire _13266_;
 wire _13267_;
 wire _13268_;
 wire _13269_;
 wire _13270_;
 wire _13271_;
 wire _13272_;
 wire _13273_;
 wire _13274_;
 wire _13275_;
 wire _13276_;
 wire _13277_;
 wire _13278_;
 wire _13279_;
 wire _13280_;
 wire _13281_;
 wire _13282_;
 wire _13283_;
 wire _13284_;
 wire _13285_;
 wire _13286_;
 wire _13287_;
 wire _13288_;
 wire _13289_;
 wire _13290_;
 wire _13291_;
 wire _13292_;
 wire _13293_;
 wire _13294_;
 wire _13295_;
 wire _13296_;
 wire _13297_;
 wire _13298_;
 wire _13299_;
 wire _13300_;
 wire _13301_;
 wire _13302_;
 wire _13303_;
 wire _13304_;
 wire _13305_;
 wire _13306_;
 wire _13307_;
 wire _13308_;
 wire _13309_;
 wire _13310_;
 wire _13311_;
 wire _13312_;
 wire _13313_;
 wire _13314_;
 wire _13315_;
 wire _13316_;
 wire _13317_;
 wire _13318_;
 wire _13319_;
 wire _13320_;
 wire _13321_;
 wire _13322_;
 wire _13323_;
 wire _13324_;
 wire _13325_;
 wire _13326_;
 wire _13327_;
 wire _13328_;
 wire _13329_;
 wire _13330_;
 wire _13331_;
 wire _13332_;
 wire _13333_;
 wire _13334_;
 wire _13335_;
 wire _13336_;
 wire _13337_;
 wire _13338_;
 wire _13339_;
 wire _13340_;
 wire _13341_;
 wire _13342_;
 wire _13343_;
 wire _13344_;
 wire _13345_;
 wire _13346_;
 wire _13347_;
 wire _13348_;
 wire _13349_;
 wire _13350_;
 wire _13351_;
 wire _13352_;
 wire _13353_;
 wire _13354_;
 wire _13355_;
 wire _13356_;
 wire _13357_;
 wire _13358_;
 wire _13359_;
 wire _13360_;
 wire _13361_;
 wire _13362_;
 wire _13363_;
 wire _13364_;
 wire _13365_;
 wire _13366_;
 wire _13367_;
 wire _13368_;
 wire _13369_;
 wire _13370_;
 wire _13371_;
 wire _13372_;
 wire _13373_;
 wire _13374_;
 wire _13375_;
 wire _13376_;
 wire _13377_;
 wire _13378_;
 wire _13379_;
 wire _13380_;
 wire _13381_;
 wire _13382_;
 wire _13383_;
 wire _13384_;
 wire _13385_;
 wire _13386_;
 wire _13387_;
 wire _13388_;
 wire _13389_;
 wire _13390_;
 wire _13391_;
 wire _13392_;
 wire _13393_;
 wire _13394_;
 wire _13395_;
 wire _13396_;
 wire _13397_;
 wire _13398_;
 wire _13399_;
 wire _13400_;
 wire _13401_;
 wire _13402_;
 wire _13403_;
 wire _13404_;
 wire _13405_;
 wire _13406_;
 wire _13407_;
 wire _13408_;
 wire _13409_;
 wire _13410_;
 wire _13411_;
 wire _13412_;
 wire _13413_;
 wire _13414_;
 wire _13415_;
 wire _13416_;
 wire _13417_;
 wire _13418_;
 wire _13419_;
 wire _13420_;
 wire _13421_;
 wire _13422_;
 wire _13423_;
 wire _13424_;
 wire _13425_;
 wire _13426_;
 wire _13427_;
 wire _13428_;
 wire _13429_;
 wire _13430_;
 wire _13431_;
 wire _13432_;
 wire _13433_;
 wire _13434_;
 wire _13435_;
 wire _13436_;
 wire _13437_;
 wire _13438_;
 wire _13439_;
 wire _13440_;
 wire _13441_;
 wire _13442_;
 wire _13443_;
 wire _13444_;
 wire _13445_;
 wire _13446_;
 wire _13447_;
 wire _13448_;
 wire _13449_;
 wire _13450_;
 wire _13451_;
 wire _13452_;
 wire _13453_;
 wire _13454_;
 wire _13455_;
 wire _13456_;
 wire _13457_;
 wire _13458_;
 wire _13459_;
 wire _13460_;
 wire _13461_;
 wire _13462_;
 wire _13463_;
 wire _13464_;
 wire _13465_;
 wire _13466_;
 wire _13467_;
 wire _13468_;
 wire _13469_;
 wire _13470_;
 wire _13471_;
 wire _13472_;
 wire _13473_;
 wire _13474_;
 wire _13475_;
 wire _13476_;
 wire _13477_;
 wire _13478_;
 wire _13479_;
 wire _13480_;
 wire _13481_;
 wire _13482_;
 wire _13483_;
 wire _13484_;
 wire _13485_;
 wire _13486_;
 wire _13487_;
 wire _13488_;
 wire _13489_;
 wire _13490_;
 wire _13491_;
 wire _13492_;
 wire _13493_;
 wire _13494_;
 wire _13495_;
 wire _13496_;
 wire _13497_;
 wire _13498_;
 wire _13499_;
 wire _13500_;
 wire _13501_;
 wire _13502_;
 wire _13503_;
 wire _13504_;
 wire _13505_;
 wire _13506_;
 wire _13507_;
 wire _13508_;
 wire _13509_;
 wire _13510_;
 wire _13511_;
 wire _13512_;
 wire _13513_;
 wire _13514_;
 wire _13515_;
 wire _13516_;
 wire _13517_;
 wire _13518_;
 wire _13519_;
 wire _13520_;
 wire _13521_;
 wire _13522_;
 wire _13523_;
 wire _13524_;
 wire _13525_;
 wire _13526_;
 wire _13527_;
 wire _13528_;
 wire _13529_;
 wire _13530_;
 wire _13531_;
 wire _13532_;
 wire _13533_;
 wire _13534_;
 wire _13535_;
 wire _13536_;
 wire _13537_;
 wire _13538_;
 wire _13539_;
 wire _13540_;
 wire _13541_;
 wire _13542_;
 wire _13543_;
 wire _13544_;
 wire _13546_;
 wire _13547_;
 wire _13548_;
 wire _13549_;
 wire _13550_;
 wire _13551_;
 wire _13552_;
 wire _13553_;
 wire _13554_;
 wire _13555_;
 wire _13556_;
 wire _13557_;
 wire _13558_;
 wire _13559_;
 wire _13560_;
 wire _13561_;
 wire _13562_;
 wire _13563_;
 wire _13564_;
 wire _13565_;
 wire _13566_;
 wire _13567_;
 wire _13568_;
 wire _13569_;
 wire _13570_;
 wire _13571_;
 wire _13573_;
 wire _13574_;
 wire _13575_;
 wire _13576_;
 wire _13578_;
 wire _13579_;
 wire _13580_;
 wire net4479;
 wire _13582_;
 wire _13583_;
 wire _13584_;
 wire _13585_;
 wire _13586_;
 wire _13587_;
 wire _13588_;
 wire _13589_;
 wire _13590_;
 wire _13591_;
 wire _13592_;
 wire _13593_;
 wire _13594_;
 wire _13595_;
 wire net4478;
 wire _13597_;
 wire _13598_;
 wire _13599_;
 wire _13600_;
 wire _13601_;
 wire _13602_;
 wire _13603_;
 wire _13604_;
 wire _13605_;
 wire _13606_;
 wire _13607_;
 wire _13608_;
 wire _13609_;
 wire _13610_;
 wire _13611_;
 wire _13612_;
 wire _13613_;
 wire _13614_;
 wire _13615_;
 wire _13616_;
 wire net4476;
 wire _13618_;
 wire _13619_;
 wire _13620_;
 wire _13621_;
 wire _13622_;
 wire _13623_;
 wire _13624_;
 wire _13625_;
 wire _13626_;
 wire _13627_;
 wire _13628_;
 wire net4477;
 wire _13630_;
 wire net4475;
 wire _13632_;
 wire _13633_;
 wire _13634_;
 wire _13635_;
 wire _13636_;
 wire _13637_;
 wire _13638_;
 wire _13639_;
 wire net4473;
 wire _13641_;
 wire _13642_;
 wire _13643_;
 wire _13644_;
 wire _13645_;
 wire net4472;
 wire net4470;
 wire _13648_;
 wire _13649_;
 wire net4469;
 wire _13651_;
 wire _13652_;
 wire net4468;
 wire _13654_;
 wire _13655_;
 wire net4466;
 wire _13657_;
 wire _13658_;
 wire _13659_;
 wire net4467;
 wire _13661_;
 wire net4471;
 wire _13663_;
 wire _13664_;
 wire _13665_;
 wire _13666_;
 wire _13667_;
 wire _13668_;
 wire _13669_;
 wire _13670_;
 wire _13671_;
 wire _13672_;
 wire _13673_;
 wire _13674_;
 wire _13675_;
 wire _13676_;
 wire _13677_;
 wire _13678_;
 wire net4463;
 wire net4462;
 wire _13681_;
 wire _13682_;
 wire net4459;
 wire net4460;
 wire _13685_;
 wire _13686_;
 wire _13687_;
 wire net4464;
 wire _13689_;
 wire _13690_;
 wire _13691_;
 wire _13692_;
 wire net4461;
 wire _13694_;
 wire net4458;
 wire _13696_;
 wire _13697_;
 wire _13698_;
 wire net4465;
 wire _13700_;
 wire _13701_;
 wire _13702_;
 wire net4456;
 wire _13704_;
 wire net4455;
 wire _13706_;
 wire _13707_;
 wire net4453;
 wire net4451;
 wire _13710_;
 wire _13711_;
 wire _13712_;
 wire _13713_;
 wire _13714_;
 wire net4450;
 wire _13716_;
 wire _13717_;
 wire _13718_;
 wire _13719_;
 wire _13720_;
 wire _13721_;
 wire _13722_;
 wire _13723_;
 wire _13724_;
 wire _13725_;
 wire _13726_;
 wire _13727_;
 wire _13728_;
 wire net4449;
 wire _13730_;
 wire _13731_;
 wire net4447;
 wire _13733_;
 wire _13734_;
 wire _13735_;
 wire _13736_;
 wire _13737_;
 wire _13738_;
 wire net4446;
 wire _13740_;
 wire _13741_;
 wire _13742_;
 wire net4448;
 wire net4445;
 wire _13745_;
 wire _13746_;
 wire _13747_;
 wire net4443;
 wire _13749_;
 wire _13750_;
 wire _13751_;
 wire net4444;
 wire _13753_;
 wire _13754_;
 wire _13755_;
 wire _13756_;
 wire net4442;
 wire _13758_;
 wire _13759_;
 wire net4441;
 wire _13761_;
 wire _13762_;
 wire _13763_;
 wire _13764_;
 wire _13765_;
 wire _13766_;
 wire _13767_;
 wire _13768_;
 wire _13769_;
 wire _13770_;
 wire _13771_;
 wire _13772_;
 wire _13773_;
 wire net4452;
 wire net4440;
 wire _13776_;
 wire net4439;
 wire _13778_;
 wire _13779_;
 wire _13780_;
 wire net4437;
 wire _13782_;
 wire _13783_;
 wire _13784_;
 wire _13785_;
 wire _13786_;
 wire _13787_;
 wire _13788_;
 wire net4436;
 wire _13790_;
 wire _13791_;
 wire _13792_;
 wire _13793_;
 wire _13794_;
 wire _13795_;
 wire _13796_;
 wire _13797_;
 wire _13798_;
 wire _13799_;
 wire _13800_;
 wire _13801_;
 wire _13802_;
 wire _13803_;
 wire _13804_;
 wire _13805_;
 wire _13806_;
 wire _13807_;
 wire _13808_;
 wire _13809_;
 wire _13810_;
 wire _13811_;
 wire _13812_;
 wire _13813_;
 wire _13814_;
 wire _13815_;
 wire _13816_;
 wire _13817_;
 wire _13818_;
 wire _13819_;
 wire _13820_;
 wire _13821_;
 wire _13822_;
 wire _13823_;
 wire _13824_;
 wire _13825_;
 wire _13826_;
 wire _13827_;
 wire _13828_;
 wire net4434;
 wire _13830_;
 wire _13831_;
 wire _13832_;
 wire _13833_;
 wire _13834_;
 wire _13835_;
 wire _13836_;
 wire _13837_;
 wire _13838_;
 wire _13839_;
 wire _13840_;
 wire _13841_;
 wire _13842_;
 wire _13843_;
 wire _13844_;
 wire _13845_;
 wire _13846_;
 wire _13847_;
 wire _13848_;
 wire _13849_;
 wire _13850_;
 wire _13851_;
 wire _13852_;
 wire _13853_;
 wire _13854_;
 wire _13855_;
 wire _13856_;
 wire _13857_;
 wire _13858_;
 wire _13859_;
 wire _13860_;
 wire _13861_;
 wire _13862_;
 wire _13863_;
 wire _13864_;
 wire _13865_;
 wire _13866_;
 wire _13867_;
 wire _13868_;
 wire _13869_;
 wire _13870_;
 wire _13871_;
 wire _13872_;
 wire _13873_;
 wire _13874_;
 wire _13875_;
 wire _13876_;
 wire _13877_;
 wire _13878_;
 wire _13879_;
 wire _13880_;
 wire _13881_;
 wire _13882_;
 wire net4435;
 wire _13884_;
 wire net4433;
 wire _13886_;
 wire _13887_;
 wire _13888_;
 wire _13889_;
 wire _13890_;
 wire _13891_;
 wire _13892_;
 wire _13893_;
 wire _13894_;
 wire _13895_;
 wire _13896_;
 wire _13897_;
 wire _13898_;
 wire _13899_;
 wire _13900_;
 wire _13901_;
 wire _13902_;
 wire _13903_;
 wire _13904_;
 wire _13905_;
 wire _13906_;
 wire _13907_;
 wire _13908_;
 wire _13909_;
 wire _13910_;
 wire _13911_;
 wire _13912_;
 wire _13913_;
 wire _13914_;
 wire _13915_;
 wire _13916_;
 wire _13917_;
 wire _13918_;
 wire _13919_;
 wire _13920_;
 wire _13921_;
 wire _13922_;
 wire _13923_;
 wire _13924_;
 wire _13925_;
 wire _13926_;
 wire _13927_;
 wire _13928_;
 wire _13929_;
 wire _13930_;
 wire _13931_;
 wire _13932_;
 wire _13933_;
 wire _13934_;
 wire _13935_;
 wire _13936_;
 wire _13937_;
 wire _13938_;
 wire _13939_;
 wire _13940_;
 wire _13941_;
 wire _13942_;
 wire _13943_;
 wire _13944_;
 wire _13945_;
 wire _13946_;
 wire _13947_;
 wire _13948_;
 wire _13949_;
 wire _13950_;
 wire _13951_;
 wire _13952_;
 wire _13953_;
 wire _13954_;
 wire _13955_;
 wire _13956_;
 wire _13957_;
 wire _13958_;
 wire _13959_;
 wire _13960_;
 wire _13961_;
 wire _13962_;
 wire _13963_;
 wire _13964_;
 wire _13965_;
 wire _13966_;
 wire _13967_;
 wire _13968_;
 wire _13969_;
 wire _13970_;
 wire _13971_;
 wire _13972_;
 wire _13973_;
 wire _13974_;
 wire _13975_;
 wire _13976_;
 wire _13977_;
 wire _13978_;
 wire _13979_;
 wire _13980_;
 wire _13981_;
 wire _13982_;
 wire _13983_;
 wire _13984_;
 wire _13985_;
 wire _13986_;
 wire _13987_;
 wire _13988_;
 wire _13989_;
 wire _13990_;
 wire _13991_;
 wire _13992_;
 wire _13993_;
 wire _13994_;
 wire _13995_;
 wire _13996_;
 wire _13997_;
 wire _13998_;
 wire _13999_;
 wire _14000_;
 wire _14001_;
 wire _14002_;
 wire _14003_;
 wire _14004_;
 wire _14005_;
 wire _14006_;
 wire _14007_;
 wire _14008_;
 wire _14009_;
 wire _14010_;
 wire _14011_;
 wire _14012_;
 wire _14013_;
 wire _14014_;
 wire _14015_;
 wire _14016_;
 wire _14017_;
 wire _14018_;
 wire _14019_;
 wire _14020_;
 wire _14021_;
 wire _14022_;
 wire _14023_;
 wire _14024_;
 wire _14025_;
 wire _14026_;
 wire _14027_;
 wire _14028_;
 wire _14029_;
 wire _14030_;
 wire _14031_;
 wire _14032_;
 wire _14033_;
 wire _14034_;
 wire _14035_;
 wire _14036_;
 wire _14037_;
 wire _14038_;
 wire _14039_;
 wire _14040_;
 wire _14041_;
 wire _14042_;
 wire _14043_;
 wire _14044_;
 wire _14045_;
 wire _14046_;
 wire _14047_;
 wire _14048_;
 wire _14049_;
 wire _14050_;
 wire _14051_;
 wire _14052_;
 wire _14053_;
 wire _14054_;
 wire _14055_;
 wire _14056_;
 wire _14057_;
 wire _14058_;
 wire _14059_;
 wire _14060_;
 wire _14061_;
 wire _14062_;
 wire _14063_;
 wire _14064_;
 wire _14065_;
 wire _14066_;
 wire _14067_;
 wire _14068_;
 wire _14069_;
 wire _14070_;
 wire _14071_;
 wire _14072_;
 wire _14073_;
 wire _14074_;
 wire _14075_;
 wire _14076_;
 wire _14077_;
 wire _14078_;
 wire _14079_;
 wire _14080_;
 wire _14081_;
 wire _14082_;
 wire _14083_;
 wire _14084_;
 wire _14085_;
 wire _14086_;
 wire _14087_;
 wire _14088_;
 wire _14089_;
 wire _14090_;
 wire _14091_;
 wire _14092_;
 wire _14093_;
 wire _14094_;
 wire _14095_;
 wire _14096_;
 wire _14097_;
 wire _14098_;
 wire _14099_;
 wire _14100_;
 wire _14101_;
 wire _14102_;
 wire _14103_;
 wire _14104_;
 wire _14105_;
 wire _14106_;
 wire _14107_;
 wire _14108_;
 wire _14109_;
 wire _14110_;
 wire _14111_;
 wire _14112_;
 wire _14113_;
 wire _14114_;
 wire _14115_;
 wire _14116_;
 wire _14117_;
 wire _14118_;
 wire _14119_;
 wire _14120_;
 wire _14121_;
 wire _14122_;
 wire _14123_;
 wire _14124_;
 wire _14125_;
 wire _14126_;
 wire _14127_;
 wire _14128_;
 wire _14129_;
 wire _14130_;
 wire _14131_;
 wire _14132_;
 wire _14133_;
 wire _14134_;
 wire _14135_;
 wire _14136_;
 wire _14137_;
 wire _14138_;
 wire _14139_;
 wire _14140_;
 wire _14141_;
 wire _14142_;
 wire _14143_;
 wire _14144_;
 wire _14145_;
 wire _14146_;
 wire _14147_;
 wire _14148_;
 wire _14149_;
 wire _14150_;
 wire _14151_;
 wire _14152_;
 wire _14153_;
 wire _14154_;
 wire _14155_;
 wire _14156_;
 wire _14157_;
 wire _14158_;
 wire _14159_;
 wire _14160_;
 wire _14161_;
 wire _14162_;
 wire _14163_;
 wire _14164_;
 wire _14165_;
 wire _14166_;
 wire _14167_;
 wire _14168_;
 wire _14169_;
 wire _14170_;
 wire _14171_;
 wire _14172_;
 wire _14173_;
 wire _14174_;
 wire _14175_;
 wire _14176_;
 wire _14177_;
 wire _14178_;
 wire _14179_;
 wire _14180_;
 wire _14181_;
 wire _14182_;
 wire _14183_;
 wire _14184_;
 wire _14185_;
 wire _14186_;
 wire _14187_;
 wire _14188_;
 wire _14189_;
 wire _14190_;
 wire _14191_;
 wire _14192_;
 wire _14193_;
 wire _14194_;
 wire _14195_;
 wire _14196_;
 wire _14197_;
 wire _14198_;
 wire _14199_;
 wire _14200_;
 wire _14201_;
 wire _14202_;
 wire _14203_;
 wire _14204_;
 wire _14205_;
 wire _14206_;
 wire _14207_;
 wire _14208_;
 wire _14209_;
 wire _14210_;
 wire _14211_;
 wire _14212_;
 wire _14213_;
 wire _14214_;
 wire _14215_;
 wire _14216_;
 wire _14217_;
 wire _14218_;
 wire _14219_;
 wire _14220_;
 wire _14221_;
 wire _14222_;
 wire _14223_;
 wire _14224_;
 wire _14225_;
 wire _14226_;
 wire _14227_;
 wire _14228_;
 wire _14229_;
 wire _14230_;
 wire _14231_;
 wire _14232_;
 wire _14233_;
 wire _14234_;
 wire _14235_;
 wire _14236_;
 wire _14237_;
 wire _14238_;
 wire _14239_;
 wire _14240_;
 wire _14241_;
 wire _14242_;
 wire _14243_;
 wire _14244_;
 wire _14245_;
 wire _14246_;
 wire _14247_;
 wire _14248_;
 wire _14249_;
 wire _14250_;
 wire _14251_;
 wire _14252_;
 wire _14253_;
 wire _14254_;
 wire _14255_;
 wire _14256_;
 wire _14257_;
 wire _14258_;
 wire _14259_;
 wire _14260_;
 wire _14261_;
 wire _14262_;
 wire _14263_;
 wire _14264_;
 wire _14265_;
 wire _14266_;
 wire net4425;
 wire _14268_;
 wire _14269_;
 wire _14270_;
 wire net4431;
 wire _14272_;
 wire _14273_;
 wire _14274_;
 wire _14275_;
 wire _14276_;
 wire _14277_;
 wire _14278_;
 wire _14279_;
 wire _14280_;
 wire _14281_;
 wire _14282_;
 wire _14283_;
 wire _14284_;
 wire _14285_;
 wire _14286_;
 wire _14287_;
 wire net4430;
 wire net4428;
 wire _14290_;
 wire net4424;
 wire _14292_;
 wire clknet_leaf_5_clk;
 wire _14294_;
 wire net6685;
 wire _14296_;
 wire _14297_;
 wire _14298_;
 wire _14299_;
 wire _14300_;
 wire _14301_;
 wire _14302_;
 wire _14303_;
 wire _14304_;
 wire _14305_;
 wire _14306_;
 wire _14307_;
 wire net6684;
 wire _14309_;
 wire _14310_;
 wire _14311_;
 wire _14312_;
 wire _14313_;
 wire _14314_;
 wire net6680;
 wire _14316_;
 wire _14317_;
 wire _14318_;
 wire _14319_;
 wire net6683;
 wire _14321_;
 wire _14322_;
 wire _14323_;
 wire clknet_leaf_11_clk;
 wire _14325_;
 wire _14326_;
 wire _14327_;
 wire _14328_;
 wire _14329_;
 wire _14330_;
 wire _14331_;
 wire _14332_;
 wire _14333_;
 wire _14334_;
 wire _14335_;
 wire _14336_;
 wire _14337_;
 wire _14338_;
 wire _14339_;
 wire net6674;
 wire _14341_;
 wire _14342_;
 wire _14343_;
 wire _14344_;
 wire _14345_;
 wire _14346_;
 wire _14347_;
 wire _14348_;
 wire _14349_;
 wire _14350_;
 wire _14351_;
 wire net6465;
 wire _14353_;
 wire _14355_;
 wire _14357_;
 wire net6382;
 wire _14360_;
 wire _14361_;
 wire _14362_;
 wire _14363_;
 wire _14364_;
 wire _14365_;
 wire _14366_;
 wire _14367_;
 wire _14368_;
 wire _14370_;
 wire _14371_;
 wire _14372_;
 wire _14373_;
 wire _14374_;
 wire _14375_;
 wire net6327;
 wire _14378_;
 wire net6325;
 wire _14380_;
 wire _14381_;
 wire net6324;
 wire _14383_;
 wire _14384_;
 wire _14385_;
 wire _14386_;
 wire net6323;
 wire _14388_;
 wire _14389_;
 wire _14390_;
 wire _14391_;
 wire _14392_;
 wire _14393_;
 wire net6321;
 wire _14396_;
 wire _14397_;
 wire _14398_;
 wire _14399_;
 wire _14400_;
 wire _14401_;
 wire _14403_;
 wire _14404_;
 wire _14405_;
 wire _14406_;
 wire _14407_;
 wire _14408_;
 wire _14409_;
 wire _14410_;
 wire _14411_;
 wire _14412_;
 wire _14413_;
 wire _14414_;
 wire _14415_;
 wire _14416_;
 wire _14417_;
 wire _14418_;
 wire _14419_;
 wire _14420_;
 wire _14421_;
 wire net6311;
 wire _14423_;
 wire net6310;
 wire _14425_;
 wire _14426_;
 wire net6309;
 wire _14428_;
 wire net6318;
 wire _14431_;
 wire _14434_;
 wire _14435_;
 wire _14436_;
 wire _14437_;
 wire _14438_;
 wire _14439_;
 wire _14440_;
 wire _14441_;
 wire _14442_;
 wire _14443_;
 wire _14444_;
 wire _14445_;
 wire _14446_;
 wire _14447_;
 wire _14448_;
 wire _14449_;
 wire _14450_;
 wire net6302;
 wire _14452_;
 wire _14453_;
 wire _14454_;
 wire _14455_;
 wire net6301;
 wire net6299;
 wire _14458_;
 wire _14459_;
 wire _14460_;
 wire _14461_;
 wire _14462_;
 wire _14463_;
 wire _14465_;
 wire net6297;
 wire _14467_;
 wire _14468_;
 wire _14469_;
 wire _14470_;
 wire _14471_;
 wire _14472_;
 wire _14474_;
 wire _14475_;
 wire _14476_;
 wire _14477_;
 wire _14478_;
 wire _14479_;
 wire _14480_;
 wire _14481_;
 wire _14482_;
 wire _14483_;
 wire _14484_;
 wire _14485_;
 wire net6296;
 wire _14487_;
 wire _14489_;
 wire _14490_;
 wire _14491_;
 wire _14492_;
 wire _14493_;
 wire _14494_;
 wire _14495_;
 wire _14496_;
 wire _14497_;
 wire _14498_;
 wire _14499_;
 wire _14500_;
 wire _14501_;
 wire _14502_;
 wire _14503_;
 wire _14504_;
 wire _14505_;
 wire net6156;
 wire _14507_;
 wire _14508_;
 wire _14509_;
 wire _14510_;
 wire _14511_;
 wire _14512_;
 wire _14513_;
 wire _14514_;
 wire _14515_;
 wire _14516_;
 wire _14517_;
 wire _14518_;
 wire _14519_;
 wire _14520_;
 wire _14521_;
 wire _14522_;
 wire _14523_;
 wire _14524_;
 wire _14525_;
 wire _14526_;
 wire _14527_;
 wire _14528_;
 wire _14529_;
 wire _14530_;
 wire _14531_;
 wire _14532_;
 wire net6115;
 wire _14534_;
 wire _14535_;
 wire _14536_;
 wire _14537_;
 wire _14538_;
 wire _14539_;
 wire _14540_;
 wire _14541_;
 wire net6102;
 wire _14543_;
 wire _14544_;
 wire _14545_;
 wire _14546_;
 wire _14547_;
 wire _14548_;
 wire _14549_;
 wire _14550_;
 wire _14551_;
 wire _14552_;
 wire _14553_;
 wire _14554_;
 wire _14555_;
 wire _14556_;
 wire _14557_;
 wire _14558_;
 wire _14559_;
 wire _14560_;
 wire _14561_;
 wire _14562_;
 wire _14563_;
 wire _14564_;
 wire _14565_;
 wire _14566_;
 wire _14567_;
 wire _14568_;
 wire _14569_;
 wire _14570_;
 wire _14571_;
 wire _14572_;
 wire _14573_;
 wire _14574_;
 wire _14575_;
 wire _14576_;
 wire _14577_;
 wire _14578_;
 wire _14579_;
 wire _14580_;
 wire _14581_;
 wire _14582_;
 wire _14583_;
 wire _14584_;
 wire _14585_;
 wire _14586_;
 wire _14587_;
 wire _14588_;
 wire _14589_;
 wire _14590_;
 wire _14591_;
 wire _14592_;
 wire _14593_;
 wire _14594_;
 wire _14595_;
 wire _14596_;
 wire _14597_;
 wire _14598_;
 wire _14599_;
 wire _14600_;
 wire _14601_;
 wire _14602_;
 wire _14603_;
 wire _14604_;
 wire _14605_;
 wire _14606_;
 wire _14607_;
 wire _14608_;
 wire _14609_;
 wire _14610_;
 wire _14611_;
 wire _14612_;
 wire _14613_;
 wire _14614_;
 wire _14615_;
 wire _14616_;
 wire _14617_;
 wire _14618_;
 wire _14619_;
 wire _14620_;
 wire _14621_;
 wire _14622_;
 wire _14623_;
 wire _14624_;
 wire _14625_;
 wire _14626_;
 wire _14627_;
 wire _14628_;
 wire _14629_;
 wire _14630_;
 wire _14631_;
 wire _14632_;
 wire _14633_;
 wire _14634_;
 wire _14635_;
 wire _14636_;
 wire _14637_;
 wire _14638_;
 wire _14639_;
 wire _14640_;
 wire _14641_;
 wire _14642_;
 wire _14643_;
 wire _14644_;
 wire _14645_;
 wire _14646_;
 wire _14647_;
 wire _14648_;
 wire _14649_;
 wire _14650_;
 wire _14651_;
 wire _14652_;
 wire _14653_;
 wire _14654_;
 wire _14655_;
 wire _14656_;
 wire _14657_;
 wire _14658_;
 wire _14659_;
 wire _14660_;
 wire _14661_;
 wire _14662_;
 wire _14663_;
 wire _14664_;
 wire _14665_;
 wire _14666_;
 wire _14667_;
 wire _14668_;
 wire _14669_;
 wire _14670_;
 wire _14671_;
 wire _14672_;
 wire _14673_;
 wire _14674_;
 wire _14675_;
 wire _14676_;
 wire _14677_;
 wire _14678_;
 wire _14679_;
 wire _14680_;
 wire _14681_;
 wire _14682_;
 wire _14683_;
 wire _14684_;
 wire _14685_;
 wire _14686_;
 wire _14687_;
 wire _14688_;
 wire _14689_;
 wire _14690_;
 wire _14691_;
 wire _14692_;
 wire _14693_;
 wire _14694_;
 wire _14695_;
 wire _14696_;
 wire _14697_;
 wire _14698_;
 wire _14699_;
 wire _14700_;
 wire _14701_;
 wire _14702_;
 wire _14703_;
 wire _14704_;
 wire _14705_;
 wire _14706_;
 wire _14707_;
 wire _14708_;
 wire _14709_;
 wire _14710_;
 wire _14711_;
 wire _14712_;
 wire _14713_;
 wire _14714_;
 wire _14715_;
 wire _14716_;
 wire _14717_;
 wire _14718_;
 wire _14719_;
 wire _14720_;
 wire _14721_;
 wire _14722_;
 wire _14723_;
 wire _14724_;
 wire _14725_;
 wire _14726_;
 wire _14727_;
 wire _14728_;
 wire _14729_;
 wire _14730_;
 wire _14731_;
 wire _14732_;
 wire _14733_;
 wire _14734_;
 wire _14735_;
 wire _14736_;
 wire _14737_;
 wire _14738_;
 wire _14739_;
 wire _14740_;
 wire _14741_;
 wire _14742_;
 wire _14743_;
 wire _14744_;
 wire _14745_;
 wire _14746_;
 wire _14747_;
 wire _14748_;
 wire _14749_;
 wire _14750_;
 wire _14751_;
 wire _14752_;
 wire _14753_;
 wire _14754_;
 wire _14755_;
 wire _14756_;
 wire _14757_;
 wire _14758_;
 wire _14759_;
 wire _14760_;
 wire _14761_;
 wire _14762_;
 wire _14763_;
 wire _14764_;
 wire _14765_;
 wire _14766_;
 wire _14767_;
 wire _14768_;
 wire _14769_;
 wire _14770_;
 wire _14771_;
 wire _14772_;
 wire _14773_;
 wire _14774_;
 wire _14775_;
 wire _14776_;
 wire _14777_;
 wire _14778_;
 wire _14779_;
 wire _14780_;
 wire _14781_;
 wire _14782_;
 wire _14783_;
 wire _14784_;
 wire _14785_;
 wire _14786_;
 wire _14787_;
 wire _14788_;
 wire _14789_;
 wire _14790_;
 wire _14791_;
 wire _14792_;
 wire _14793_;
 wire _14794_;
 wire _14795_;
 wire _14796_;
 wire _14797_;
 wire _14798_;
 wire _14799_;
 wire _14800_;
 wire _14801_;
 wire _14802_;
 wire _14803_;
 wire _14804_;
 wire _14805_;
 wire _14806_;
 wire _14807_;
 wire _14808_;
 wire _14809_;
 wire _14810_;
 wire _14811_;
 wire _14812_;
 wire _14813_;
 wire _14814_;
 wire _14815_;
 wire _14816_;
 wire _14817_;
 wire _14818_;
 wire _14819_;
 wire _14820_;
 wire _14821_;
 wire _14822_;
 wire _14823_;
 wire _14824_;
 wire _14825_;
 wire _14826_;
 wire _14827_;
 wire _14828_;
 wire _14829_;
 wire _14830_;
 wire _14831_;
 wire _14832_;
 wire _14833_;
 wire _14834_;
 wire _14835_;
 wire _14836_;
 wire _14837_;
 wire _14838_;
 wire _14839_;
 wire _14840_;
 wire _14841_;
 wire _14842_;
 wire _14843_;
 wire _14844_;
 wire _14845_;
 wire _14846_;
 wire _14847_;
 wire _14848_;
 wire _14849_;
 wire _14850_;
 wire _14851_;
 wire _14852_;
 wire _14853_;
 wire _14854_;
 wire _14855_;
 wire _14856_;
 wire _14857_;
 wire _14858_;
 wire _14859_;
 wire _14860_;
 wire _14861_;
 wire _14862_;
 wire _14863_;
 wire _14864_;
 wire _14865_;
 wire _14866_;
 wire _14867_;
 wire _14868_;
 wire _14869_;
 wire _14870_;
 wire _14871_;
 wire _14872_;
 wire _14873_;
 wire _14874_;
 wire _14875_;
 wire _14876_;
 wire _14877_;
 wire _14878_;
 wire _14879_;
 wire _14880_;
 wire _14881_;
 wire _14882_;
 wire _14883_;
 wire _14884_;
 wire _14885_;
 wire _14886_;
 wire _14887_;
 wire _14888_;
 wire _14889_;
 wire _14890_;
 wire _14891_;
 wire _14892_;
 wire _14893_;
 wire _14894_;
 wire _14895_;
 wire _14896_;
 wire _14897_;
 wire _14898_;
 wire _14899_;
 wire _14900_;
 wire _14901_;
 wire _14902_;
 wire _14903_;
 wire _14904_;
 wire _14905_;
 wire _14906_;
 wire _14907_;
 wire _14908_;
 wire _14909_;
 wire _14910_;
 wire _14911_;
 wire _14912_;
 wire _14913_;
 wire _14914_;
 wire _14915_;
 wire _14916_;
 wire _14917_;
 wire _14918_;
 wire _14919_;
 wire _14920_;
 wire _14921_;
 wire _14922_;
 wire _14923_;
 wire _14924_;
 wire _14925_;
 wire _14926_;
 wire _14927_;
 wire _14928_;
 wire _14929_;
 wire _14930_;
 wire _14931_;
 wire _14932_;
 wire _14933_;
 wire _14934_;
 wire _14935_;
 wire _14936_;
 wire _14937_;
 wire _14938_;
 wire _14939_;
 wire _14940_;
 wire _14941_;
 wire _14942_;
 wire _14943_;
 wire _14944_;
 wire _14945_;
 wire _14946_;
 wire _14947_;
 wire _14948_;
 wire _14949_;
 wire _14950_;
 wire _14951_;
 wire _14952_;
 wire _14953_;
 wire _14954_;
 wire _14955_;
 wire _14956_;
 wire _14957_;
 wire _14958_;
 wire _14959_;
 wire _14960_;
 wire _14961_;
 wire _14962_;
 wire _14963_;
 wire _14964_;
 wire _14965_;
 wire _14966_;
 wire _14967_;
 wire _14969_;
 wire _14970_;
 wire _14971_;
 wire _14972_;
 wire _14973_;
 wire _14974_;
 wire _14975_;
 wire _14976_;
 wire _14977_;
 wire _14978_;
 wire _14979_;
 wire _14980_;
 wire _14981_;
 wire _14982_;
 wire _14983_;
 wire _14984_;
 wire _14985_;
 wire _14986_;
 wire _14987_;
 wire _14988_;
 wire _14989_;
 wire net5941;
 wire _14991_;
 wire _14992_;
 wire _14993_;
 wire net5940;
 wire _14995_;
 wire _14996_;
 wire _14997_;
 wire _14998_;
 wire _14999_;
 wire net5947;
 wire _15002_;
 wire _15003_;
 wire _15004_;
 wire _15005_;
 wire _15006_;
 wire _15007_;
 wire _15008_;
 wire _15009_;
 wire _15010_;
 wire _15011_;
 wire _15012_;
 wire _15013_;
 wire _15014_;
 wire _15015_;
 wire _15016_;
 wire _15017_;
 wire _15018_;
 wire _15019_;
 wire _15020_;
 wire _15021_;
 wire _15022_;
 wire _15023_;
 wire _15024_;
 wire _15025_;
 wire _15026_;
 wire _15027_;
 wire _15028_;
 wire _15029_;
 wire _15030_;
 wire net5936;
 wire _15032_;
 wire net5932;
 wire _15034_;
 wire _15035_;
 wire _15037_;
 wire _15039_;
 wire _15040_;
 wire _15041_;
 wire _15042_;
 wire _15043_;
 wire _15044_;
 wire _15045_;
 wire _15046_;
 wire _15047_;
 wire _15048_;
 wire _15049_;
 wire _15050_;
 wire _15051_;
 wire net5862;
 wire _15053_;
 wire _15054_;
 wire _15055_;
 wire net5851;
 wire net5853;
 wire net5850;
 wire _15059_;
 wire _15060_;
 wire _15061_;
 wire net5846;
 wire _15063_;
 wire _15064_;
 wire net5845;
 wire _15066_;
 wire _15067_;
 wire _15068_;
 wire _15069_;
 wire _15070_;
 wire _15071_;
 wire net5855;
 wire _15073_;
 wire _15074_;
 wire _15075_;
 wire _15076_;
 wire _15077_;
 wire _15078_;
 wire _15079_;
 wire _15080_;
 wire net5854;
 wire _15082_;
 wire _15083_;
 wire _15084_;
 wire _15085_;
 wire _15086_;
 wire _15087_;
 wire net5844;
 wire _15090_;
 wire _15091_;
 wire _15092_;
 wire _15093_;
 wire _15094_;
 wire _15095_;
 wire _15097_;
 wire _15098_;
 wire _15099_;
 wire _15101_;
 wire _15102_;
 wire net5819;
 wire _15104_;
 wire net5817;
 wire _15106_;
 wire _15107_;
 wire _15109_;
 wire _15110_;
 wire _15111_;
 wire _15112_;
 wire _15114_;
 wire net5812;
 wire _15116_;
 wire _15117_;
 wire _15118_;
 wire net5811;
 wire _15120_;
 wire _15121_;
 wire net5809;
 wire _15123_;
 wire _15124_;
 wire net5808;
 wire net5802;
 wire _15127_;
 wire net5801;
 wire net5810;
 wire _15130_;
 wire _15131_;
 wire _15132_;
 wire _15133_;
 wire _15134_;
 wire _15135_;
 wire _15136_;
 wire _15137_;
 wire _15138_;
 wire _15139_;
 wire net5800;
 wire _15141_;
 wire _15142_;
 wire _15143_;
 wire _15144_;
 wire _15145_;
 wire _15146_;
 wire _15147_;
 wire net5799;
 wire _15149_;
 wire _15150_;
 wire _15151_;
 wire net5798;
 wire _15153_;
 wire _15154_;
 wire _15155_;
 wire _15156_;
 wire _15157_;
 wire _15158_;
 wire net5795;
 wire net5794;
 wire _15161_;
 wire _15162_;
 wire _15163_;
 wire _15164_;
 wire _15165_;
 wire net5796;
 wire _15167_;
 wire _15168_;
 wire _15169_;
 wire _15170_;
 wire _15171_;
 wire _15172_;
 wire _15173_;
 wire _15174_;
 wire _15175_;
 wire _15176_;
 wire _15177_;
 wire net5782;
 wire _15179_;
 wire _15180_;
 wire net5781;
 wire _15182_;
 wire _15183_;
 wire _15184_;
 wire _15185_;
 wire _15186_;
 wire _15187_;
 wire _15188_;
 wire _15189_;
 wire _15190_;
 wire _15191_;
 wire _15192_;
 wire net5789;
 wire _15194_;
 wire _15195_;
 wire _15196_;
 wire _15197_;
 wire _15198_;
 wire _15199_;
 wire _15200_;
 wire _15201_;
 wire net5779;
 wire _15203_;
 wire _15204_;
 wire _15205_;
 wire _15206_;
 wire _15207_;
 wire _15208_;
 wire _15209_;
 wire _15210_;
 wire _15211_;
 wire _15212_;
 wire _15213_;
 wire _15214_;
 wire _15215_;
 wire _15216_;
 wire _15217_;
 wire _15218_;
 wire _15219_;
 wire _15220_;
 wire _15221_;
 wire _15222_;
 wire _15223_;
 wire _15224_;
 wire _15225_;
 wire _15226_;
 wire _15227_;
 wire _15228_;
 wire _15229_;
 wire _15230_;
 wire _15231_;
 wire net5778;
 wire _15233_;
 wire _15234_;
 wire _15235_;
 wire _15236_;
 wire _15237_;
 wire _15238_;
 wire _15239_;
 wire _15240_;
 wire _15241_;
 wire _15242_;
 wire _15243_;
 wire _15245_;
 wire _15246_;
 wire _15247_;
 wire _15248_;
 wire _15249_;
 wire _15250_;
 wire _15251_;
 wire _15252_;
 wire _15253_;
 wire _15254_;
 wire _15255_;
 wire _15256_;
 wire _15257_;
 wire _15258_;
 wire _15259_;
 wire _15260_;
 wire _15261_;
 wire _15262_;
 wire _15263_;
 wire _15264_;
 wire _15265_;
 wire _15266_;
 wire _15267_;
 wire _15268_;
 wire _15269_;
 wire _15270_;
 wire _15271_;
 wire _15272_;
 wire _15273_;
 wire _15274_;
 wire _15275_;
 wire _15276_;
 wire _15277_;
 wire _15278_;
 wire _15279_;
 wire _15280_;
 wire _15281_;
 wire _15282_;
 wire _15283_;
 wire _15284_;
 wire _15286_;
 wire _15287_;
 wire _15288_;
 wire _15289_;
 wire _15290_;
 wire _15291_;
 wire _15292_;
 wire _15293_;
 wire _15294_;
 wire _15295_;
 wire _15296_;
 wire _15297_;
 wire _15298_;
 wire _15299_;
 wire _15300_;
 wire _15301_;
 wire _15302_;
 wire _15303_;
 wire _15304_;
 wire _15305_;
 wire _15306_;
 wire _15307_;
 wire _15308_;
 wire _15309_;
 wire _15310_;
 wire _15311_;
 wire _15312_;
 wire _15313_;
 wire _15314_;
 wire _15315_;
 wire _15316_;
 wire _15317_;
 wire _15318_;
 wire _15319_;
 wire _15320_;
 wire _15321_;
 wire _15322_;
 wire _15323_;
 wire _15324_;
 wire _15325_;
 wire _15326_;
 wire _15327_;
 wire _15328_;
 wire _15329_;
 wire _15330_;
 wire _15331_;
 wire _15332_;
 wire _15333_;
 wire _15334_;
 wire _15335_;
 wire _15336_;
 wire _15337_;
 wire _15338_;
 wire _15339_;
 wire _15340_;
 wire _15341_;
 wire _15342_;
 wire _15343_;
 wire _15344_;
 wire _15345_;
 wire _15346_;
 wire _15347_;
 wire _15348_;
 wire _15349_;
 wire _15350_;
 wire _15351_;
 wire _15352_;
 wire _15353_;
 wire _15354_;
 wire _15355_;
 wire _15356_;
 wire _15357_;
 wire _15358_;
 wire _15359_;
 wire _15360_;
 wire _15361_;
 wire _15362_;
 wire _15363_;
 wire _15364_;
 wire _15365_;
 wire _15366_;
 wire _15367_;
 wire _15368_;
 wire _15369_;
 wire _15370_;
 wire _15371_;
 wire _15372_;
 wire _15373_;
 wire _15374_;
 wire _15375_;
 wire _15376_;
 wire _15377_;
 wire _15378_;
 wire _15379_;
 wire _15380_;
 wire _15381_;
 wire _15382_;
 wire _15383_;
 wire _15384_;
 wire _15385_;
 wire _15386_;
 wire _15387_;
 wire _15388_;
 wire _15389_;
 wire _15390_;
 wire _15391_;
 wire _15392_;
 wire _15393_;
 wire _15394_;
 wire _15395_;
 wire _15396_;
 wire _15397_;
 wire _15398_;
 wire _15399_;
 wire _15400_;
 wire _15401_;
 wire _15402_;
 wire _15403_;
 wire _15404_;
 wire _15405_;
 wire _15406_;
 wire _15407_;
 wire _15408_;
 wire _15409_;
 wire _15410_;
 wire _15411_;
 wire _15412_;
 wire _15413_;
 wire _15414_;
 wire _15415_;
 wire _15416_;
 wire _15417_;
 wire _15418_;
 wire _15419_;
 wire _15420_;
 wire _15421_;
 wire _15422_;
 wire _15423_;
 wire _15424_;
 wire _15425_;
 wire _15426_;
 wire _15427_;
 wire _15428_;
 wire _15429_;
 wire _15430_;
 wire _15431_;
 wire _15432_;
 wire _15433_;
 wire _15434_;
 wire _15435_;
 wire _15436_;
 wire _15437_;
 wire _15438_;
 wire _15439_;
 wire _15440_;
 wire _15441_;
 wire _15442_;
 wire _15443_;
 wire _15444_;
 wire _15445_;
 wire _15446_;
 wire _15447_;
 wire _15448_;
 wire _15449_;
 wire _15450_;
 wire _15451_;
 wire _15452_;
 wire _15453_;
 wire _15454_;
 wire _15455_;
 wire _15456_;
 wire _15457_;
 wire _15458_;
 wire _15459_;
 wire _15460_;
 wire _15461_;
 wire _15462_;
 wire _15463_;
 wire _15464_;
 wire _15465_;
 wire _15466_;
 wire _15467_;
 wire _15468_;
 wire _15469_;
 wire _15470_;
 wire _15471_;
 wire _15472_;
 wire _15473_;
 wire _15474_;
 wire _15475_;
 wire _15476_;
 wire _15477_;
 wire _15478_;
 wire _15479_;
 wire _15480_;
 wire _15481_;
 wire _15482_;
 wire _15483_;
 wire _15484_;
 wire _15485_;
 wire _15486_;
 wire _15487_;
 wire _15488_;
 wire _15489_;
 wire _15490_;
 wire _15491_;
 wire _15492_;
 wire _15493_;
 wire _15494_;
 wire _15495_;
 wire _15496_;
 wire _15497_;
 wire _15498_;
 wire _15499_;
 wire _15500_;
 wire _15501_;
 wire _15502_;
 wire _15503_;
 wire _15504_;
 wire _15505_;
 wire _15506_;
 wire _15507_;
 wire _15508_;
 wire _15509_;
 wire _15510_;
 wire _15511_;
 wire _15512_;
 wire _15513_;
 wire _15514_;
 wire _15515_;
 wire _15516_;
 wire _15517_;
 wire _15518_;
 wire _15519_;
 wire _15520_;
 wire _15521_;
 wire _15522_;
 wire _15523_;
 wire _15524_;
 wire _15525_;
 wire _15526_;
 wire _15527_;
 wire _15528_;
 wire _15529_;
 wire _15530_;
 wire _15531_;
 wire _15532_;
 wire _15533_;
 wire _15534_;
 wire _15535_;
 wire _15536_;
 wire _15537_;
 wire _15538_;
 wire _15539_;
 wire _15540_;
 wire _15541_;
 wire _15542_;
 wire _15543_;
 wire _15544_;
 wire _15545_;
 wire _15546_;
 wire _15547_;
 wire _15548_;
 wire _15549_;
 wire _15550_;
 wire _15551_;
 wire _15552_;
 wire _15553_;
 wire _15554_;
 wire _15555_;
 wire _15556_;
 wire _15557_;
 wire _15558_;
 wire _15559_;
 wire _15560_;
 wire _15561_;
 wire _15562_;
 wire _15563_;
 wire _15564_;
 wire _15565_;
 wire _15566_;
 wire _15567_;
 wire _15568_;
 wire _15569_;
 wire _15570_;
 wire _15571_;
 wire _15572_;
 wire _15573_;
 wire _15574_;
 wire _15575_;
 wire _15576_;
 wire _15577_;
 wire _15578_;
 wire _15579_;
 wire _15580_;
 wire _15581_;
 wire _15582_;
 wire _15583_;
 wire _15584_;
 wire _15585_;
 wire _15586_;
 wire _15587_;
 wire _15588_;
 wire _15589_;
 wire _15590_;
 wire _15591_;
 wire _15592_;
 wire _15593_;
 wire _15594_;
 wire _15595_;
 wire _15596_;
 wire _15597_;
 wire _15598_;
 wire _15599_;
 wire _15600_;
 wire _15601_;
 wire _15602_;
 wire _15603_;
 wire _15604_;
 wire _15605_;
 wire _15606_;
 wire _15607_;
 wire _15608_;
 wire _15609_;
 wire _15610_;
 wire _15611_;
 wire _15612_;
 wire _15613_;
 wire _15614_;
 wire _15615_;
 wire _15616_;
 wire _15617_;
 wire _15618_;
 wire _15619_;
 wire _15620_;
 wire _15621_;
 wire _15622_;
 wire _15623_;
 wire _15624_;
 wire _15625_;
 wire _15626_;
 wire _15627_;
 wire _15628_;
 wire _15629_;
 wire _15630_;
 wire _15631_;
 wire _15632_;
 wire _15633_;
 wire _15634_;
 wire _15635_;
 wire _15636_;
 wire _15637_;
 wire _15638_;
 wire _15639_;
 wire _15640_;
 wire _15641_;
 wire _15642_;
 wire _15643_;
 wire _15644_;
 wire _15645_;
 wire _15646_;
 wire _15647_;
 wire _15648_;
 wire _15649_;
 wire _15650_;
 wire _15651_;
 wire _15652_;
 wire _15653_;
 wire _15654_;
 wire _15655_;
 wire _15656_;
 wire _15657_;
 wire _15658_;
 wire _15659_;
 wire _15660_;
 wire _15661_;
 wire _15662_;
 wire _15663_;
 wire _15664_;
 wire _15665_;
 wire _15666_;
 wire _15667_;
 wire _15668_;
 wire _15669_;
 wire _15670_;
 wire _15671_;
 wire _15672_;
 wire _15673_;
 wire _15674_;
 wire _15675_;
 wire _15676_;
 wire _15677_;
 wire _15678_;
 wire _15679_;
 wire _15680_;
 wire _15681_;
 wire _15682_;
 wire _15683_;
 wire _15684_;
 wire _15685_;
 wire _15686_;
 wire _15687_;
 wire _15688_;
 wire _15689_;
 wire _15690_;
 wire _15691_;
 wire _15692_;
 wire _15693_;
 wire _15694_;
 wire _15695_;
 wire _15696_;
 wire _15697_;
 wire _15698_;
 wire _15699_;
 wire _15700_;
 wire _15701_;
 wire _15702_;
 wire _15703_;
 wire _15704_;
 wire _15705_;
 wire _15706_;
 wire _15707_;
 wire _15708_;
 wire _15709_;
 wire _15710_;
 wire _15711_;
 wire _15712_;
 wire _15713_;
 wire _15714_;
 wire _15715_;
 wire _15716_;
 wire _15717_;
 wire _15718_;
 wire _15719_;
 wire _15720_;
 wire _15721_;
 wire _15722_;
 wire _15723_;
 wire _15724_;
 wire _15725_;
 wire _15726_;
 wire _15727_;
 wire _15728_;
 wire _15729_;
 wire _15730_;
 wire _15731_;
 wire _15732_;
 wire _15733_;
 wire _15734_;
 wire _15735_;
 wire _15736_;
 wire _15737_;
 wire _15738_;
 wire _15739_;
 wire _15740_;
 wire _15741_;
 wire _15742_;
 wire _15743_;
 wire _15744_;
 wire _15745_;
 wire _15746_;
 wire _15747_;
 wire _15748_;
 wire _15749_;
 wire _15750_;
 wire _15751_;
 wire _15752_;
 wire _15753_;
 wire _15754_;
 wire _15755_;
 wire _15756_;
 wire _15757_;
 wire _15758_;
 wire _15759_;
 wire _15760_;
 wire _15761_;
 wire _15762_;
 wire _15763_;
 wire _15764_;
 wire _15765_;
 wire _15766_;
 wire _15767_;
 wire _15768_;
 wire _15769_;
 wire _15770_;
 wire _15771_;
 wire _15772_;
 wire _15773_;
 wire _15774_;
 wire _15775_;
 wire _15776_;
 wire _15777_;
 wire _15778_;
 wire _15779_;
 wire _15780_;
 wire _15781_;
 wire _15782_;
 wire _15783_;
 wire _15784_;
 wire _15785_;
 wire _15786_;
 wire _15787_;
 wire _15788_;
 wire _15789_;
 wire _15790_;
 wire _15791_;
 wire _15792_;
 wire _15793_;
 wire _15794_;
 wire _15795_;
 wire _15796_;
 wire _15797_;
 wire _15798_;
 wire _15799_;
 wire _15800_;
 wire _15801_;
 wire _15802_;
 wire _15803_;
 wire _15804_;
 wire _15805_;
 wire _15806_;
 wire _15807_;
 wire _15808_;
 wire _15809_;
 wire _15810_;
 wire _15811_;
 wire _15812_;
 wire _15813_;
 wire _15814_;
 wire _15815_;
 wire _15816_;
 wire _15817_;
 wire _15818_;
 wire _15819_;
 wire _15820_;
 wire _15821_;
 wire _15822_;
 wire _15823_;
 wire _15824_;
 wire _15825_;
 wire _15826_;
 wire _15827_;
 wire _15828_;
 wire _15829_;
 wire _15830_;
 wire _15831_;
 wire _15832_;
 wire _15833_;
 wire _15834_;
 wire _15835_;
 wire _15836_;
 wire _15837_;
 wire _15838_;
 wire net259;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire \u0.r0.rcnt[0] ;
 wire \u0.r0.rcnt[1] ;
 wire \u0.r0.rcnt_next[0] ;
 wire net4865;
 wire net4866;
 wire net4867;
 wire net4868;
 wire net4869;
 wire net4870;
 wire net4871;
 wire net4872;
 wire net4873;
 wire net4874;
 wire net4875;
 wire net4876;
 wire net4877;
 wire net4878;
 wire net4883;
 wire net4879;
 wire net4880;
 wire net4881;
 wire net4882;
 wire net4884;
 wire net4885;
 wire net4887;
 wire net4886;
 wire net4888;
 wire net4889;
 wire net4890;
 wire net4893;
 wire net4892;
 wire net4891;
 wire net4894;
 wire net4895;
 wire net4896;
 wire net4897;
 wire net4898;
 wire net4899;
 wire net4901;
 wire net4900;
 wire net4902;
 wire net4903;
 wire net4904;
 wire net4906;
 wire net4905;
 wire net4907;
 wire net4911;
 wire net4908;
 wire net4909;
 wire net4910;
 wire net4912;
 wire net4913;
 wire net4914;
 wire net4915;
 wire net4916;
 wire net4918;
 wire net4917;
 wire net4919;
 wire net4935;
 wire net4920;
 wire net4933;
 wire net4921;
 wire net4924;
 wire net4923;
 wire net4922;
 wire net4928;
 wire net4925;
 wire net4927;
 wire net4926;
 wire net4929;
 wire net4930;
 wire net4931;
 wire net4932;
 wire net4934;
 wire net4936;
 wire net4937;
 wire net4938;
 wire net4939;
 wire net4943;
 wire net4940;
 wire net4941;
 wire net4942;
 wire net4944;
 wire net4945;
 wire net4946;
 wire net4947;
 wire net4950;
 wire net4948;
 wire net4949;
 wire net4951;
 wire net4952;
 wire net4953;
 wire net4954;
 wire net4955;
 wire net4956;
 wire net4957;
 wire net4958;
 wire net4959;
 wire net4960;
 wire net4961;
 wire net4962;
 wire net4963;
 wire net4964;
 wire net4965;
 wire net4966;
 wire net4967;
 wire net4971;
 wire net4968;
 wire net4969;
 wire net4970;
 wire net4972;
 wire net4973;
 wire net4974;
 wire net4975;
 wire net4976;
 wire net4977;
 wire net4978;
 wire net4979;
 wire net4980;
 wire net4981;
 wire net4982;
 wire net4983;
 wire net4984;
 wire net4985;
 wire net4987;
 wire net4986;
 wire net4988;
 wire net4990;
 wire net4989;
 wire net4991;
 wire net4992;
 wire net4998;
 wire net5002;
 wire net4993;
 wire net4997;
 wire net4994;
 wire net4995;
 wire net4996;
 wire net5000;
 wire net4999;
 wire net5001;
 wire net5007;
 wire net5003;
 wire net5004;
 wire net5005;
 wire net5006;
 wire net5008;
 wire net5019;
 wire net5009;
 wire net5011;
 wire net5010;
 wire net5012;
 wire net5013;
 wire net5015;
 wire net5014;
 wire net5016;
 wire net5017;
 wire net5018;
 wire net5026;
 wire net5025;
 wire net5023;
 wire net5020;
 wire net5021;
 wire net5022;
 wire net5024;
 wire net5027;
 wire net5028;
 wire net5029;
 wire net5030;
 wire net5031;
 wire net5032;
 wire net5033;
 wire net5034;
 wire net5036;
 wire net5035;
 wire net5037;
 wire net5038;
 wire net5045;
 wire net5039;
 wire net5044;
 wire net5041;
 wire net5040;
 wire net5042;
 wire net5043;
 wire net5052;
 wire net5046;
 wire net5047;
 wire net5048;
 wire net5049;
 wire net5050;
 wire net5051;
 wire net5053;
 wire net5054;
 wire net5055;
 wire net5056;
 wire net5057;
 wire net5058;
 wire net5059;
 wire net5060;
 wire net5061;
 wire net5062;
 wire net5063;
 wire net5064;
 wire net5065;
 wire net5066;
 wire net5067;
 wire net5068;
 wire net5069;
 wire net5070;
 wire net5071;
 wire net5072;
 wire net5073;
 wire net5074;
 wire net5076;
 wire net5075;
 wire net5083;
 wire net5077;
 wire net5081;
 wire net5078;
 wire net5080;
 wire net5079;
 wire net5082;
 wire net5084;
 wire net5085;
 wire net5089;
 wire net5086;
 wire net5088;
 wire net5087;
 wire net5090;
 wire net5091;
 wire net5092;
 wire net5093;
 wire net5099;
 wire net5094;
 wire net5095;
 wire net5096;
 wire net5097;
 wire net5098;
 wire net5102;
 wire net5100;
 wire net5101;
 wire net5103;
 wire net5104;
 wire net5106;
 wire net5105;
 wire net5107;
 wire net5108;
 wire net5109;
 wire net5110;
 wire net5111;
 wire net5114;
 wire net5112;
 wire net5113;
 wire net5115;
 wire net5118;
 wire net5116;
 wire net5117;
 wire net5119;
 wire net5120;
 wire net5121;
 wire net5122;
 wire net5123;
 wire net5124;
 wire net5125;
 wire net5126;
 wire net5130;
 wire net5127;
 wire net5128;
 wire net5129;
 wire net5131;
 wire net5132;
 wire net5133;
 wire net5134;
 wire net5135;
 wire net5136;
 wire net5139;
 wire net5137;
 wire net5138;
 wire net5141;
 wire net5140;
 wire net5142;
 wire net5143;
 wire net5145;
 wire net5144;
 wire net5155;
 wire net5154;
 wire net5153;
 wire net5152;
 wire net5151;
 wire net5147;
 wire net5146;
 wire net5150;
 wire net5149;
 wire net5148;
 wire net5158;
 wire net5157;
 wire net5159;
 wire net5160;
 wire net5161;
 wire net5162;
 wire net5164;
 wire net5163;
 wire net5165;
 wire net5166;
 wire net5167;
 wire net5168;
 wire net5169;
 wire net5170;
 wire net5171;
 wire net5173;
 wire net5172;
 wire net5174;
 wire net5175;
 wire net5176;
 wire net5177;
 wire net5178;
 wire net5179;
 wire net5180;
 wire net5181;
 wire net5182;
 wire net5183;
 wire net5184;
 wire net5191;
 wire net5185;
 wire net5186;
 wire net5187;
 wire net5189;
 wire net5188;
 wire net5190;
 wire net5192;
 wire net5193;
 wire net5194;
 wire net5195;
 wire net5196;
 wire net5197;
 wire net5198;
 wire net5199;
 wire net5200;
 wire net5201;
 wire net5202;
 wire net5203;
 wire net5204;
 wire net5206;
 wire net5205;
 wire net5207;
 wire net5208;
 wire net5209;
 wire net5210;
 wire net5211;
 wire net5221;
 wire net5212;
 wire net5220;
 wire net5217;
 wire net5213;
 wire net5214;
 wire net5215;
 wire net5216;
 wire net5218;
 wire net5219;
 wire net5222;
 wire net5223;
 wire net5224;
 wire net5228;
 wire net5226;
 wire net5225;
 wire net5227;
 wire net5229;
 wire net5230;
 wire net5231;
 wire net5232;
 wire net5233;
 wire net5234;
 wire net5235;
 wire net5236;
 wire net5237;
 wire net5238;
 wire net5239;
 wire net5240;
 wire net5241;
 wire net5242;
 wire net5245;
 wire net5243;
 wire net5244;
 wire net5246;
 wire net5247;
 wire net5248;
 wire net5249;
 wire net5250;
 wire net5251;
 wire net5252;
 wire net5257;
 wire net5253;
 wire net5254;
 wire net5255;
 wire net5256;
 wire net5258;
 wire net5259;
 wire net5260;
 wire net5261;
 wire net5263;
 wire net5262;
 wire net5264;
 wire net5265;
 wire net5266;
 wire net5268;
 wire net5267;
 wire net5270;
 wire net5269;
 wire net5271;
 wire net5272;
 wire net5274;
 wire net5273;
 wire net5275;
 wire net5276;
 wire net5277;
 wire net5279;
 wire net5278;
 wire net5280;
 wire net5281;
 wire net5282;
 wire net5283;
 wire net5284;
 wire net5285;
 wire net5286;
 wire net5287;
 wire net5288;
 wire net5289;
 wire net5290;
 wire net5291;
 wire net5292;
 wire net5293;
 wire net5294;
 wire net5295;
 wire net5296;
 wire net5297;
 wire net5298;
 wire net5299;
 wire net5300;
 wire net5301;
 wire net5302;
 wire net5303;
 wire net5308;
 wire net5306;
 wire net5304;
 wire net5305;
 wire net5307;
 wire net5309;
 wire net5310;
 wire net5311;
 wire net5318;
 wire net5314;
 wire net5312;
 wire net5313;
 wire net5315;
 wire net5316;
 wire net5317;
 wire net5319;
 wire net5320;
 wire net5321;
 wire net5322;
 wire net5323;
 wire net5324;
 wire net5325;
 wire net5326;
 wire net5327;
 wire net5328;
 wire net5329;
 wire net5330;
 wire net5331;
 wire net5332;
 wire net5333;
 wire net5334;
 wire net5337;
 wire net5335;
 wire net5336;
 wire net5341;
 wire net5338;
 wire net5339;
 wire net5340;
 wire net5345;
 wire net5342;
 wire net5343;
 wire net5344;
 wire net5346;
 wire net5349;
 wire net5347;
 wire net5350;
 wire net5348;
 wire net5351;
 wire net5353;
 wire net5352;
 wire net5354;
 wire net5355;
 wire net5356;
 wire net5360;
 wire net5357;
 wire net5358;
 wire net5359;
 wire net5361;
 wire net5362;
 wire net5363;
 wire net5364;
 wire net5365;
 wire net5366;
 wire net5367;
 wire net5368;
 wire net5370;
 wire net5377;
 wire net5371;
 wire net5376;
 wire net5369;
 wire net5372;
 wire net5374;
 wire net5373;
 wire net5375;
 wire net5379;
 wire net5378;
 wire net5380;
 wire net5381;
 wire net5382;
 wire net5383;
 wire net5385;
 wire net5384;
 wire net5387;
 wire net5386;
 wire net5388;
 wire net5389;
 wire net5393;
 wire net5392;
 wire net5390;
 wire net5394;
 wire net5391;
 wire net5398;
 wire net5397;
 wire net5395;
 wire net5396;
 wire net5400;
 wire net5399;
 wire net5403;
 wire net5402;
 wire net5401;
 wire net5404;
 wire net5405;
 wire net5411;
 wire net5410;
 wire net5409;
 wire net5408;
 wire net5406;
 wire net5407;
 wire net5412;
 wire net5414;
 wire net5413;
 wire net5415;
 wire net5419;
 wire net5416;
 wire net5418;
 wire net5417;
 wire net5420;
 wire net5422;
 wire net5421;
 wire net5424;
 wire net5423;
 wire net5426;
 wire net5425;
 wire net5429;
 wire net5427;
 wire net5428;
 wire net5433;
 wire net5432;
 wire net5431;
 wire net5430;
 wire net5435;
 wire net5434;
 wire net5437;
 wire net5438;
 wire net5443;
 wire net5441;
 wire net5439;
 wire net5440;
 wire net5442;
 wire net5446;
 wire net5445;
 wire net5444;
 wire net5447;
 wire net5448;
 wire net5451;
 wire net5449;
 wire net5450;
 wire net5452;
 wire net5454;
 wire net5453;
 wire net5456;
 wire net5455;
 wire net5458;
 wire net5457;
 wire net5459;
 wire net5460;
 wire net5461;
 wire net5462;
 wire net5475;
 wire net5465;
 wire net5463;
 wire net5464;
 wire net5466;
 wire net5473;
 wire net5471;
 wire net5470;
 wire net5469;
 wire net5468;
 wire net5467;
 wire net5472;
 wire net5474;
 wire net5479;
 wire net5478;
 wire net5477;
 wire net5476;
 wire net5481;
 wire net5482;
 wire net5487;
 wire net5486;
 wire net5484;
 wire net5483;
 wire net5485;
 wire net5488;
 wire net5489;
 wire net5492;
 wire net5491;
 wire net5490;
 wire net5495;
 wire net5493;
 wire net5494;
 wire net5499;
 wire net5500;
 wire net5498;
 wire net5496;
 wire net5497;
 wire net5501;
 wire net5502;
 wire net5503;
 wire net5504;
 wire net5505;
 wire net5506;
 wire net5508;
 wire net5507;
 wire net5509;
 wire net5514;
 wire net5510;
 wire net5511;
 wire net5512;
 wire net5513;
 wire net5516;
 wire net5515;
 wire net5517;
 wire net5518;
 wire net5519;
 wire net5520;
 wire net5521;
 wire net5522;
 wire net5524;
 wire net5523;
 wire net5525;
 wire net5526;
 wire net5527;
 wire net5528;
 wire net5529;
 wire net5530;
 wire net5532;
 wire net5531;
 wire net5533;
 wire net5534;
 wire net5535;
 wire net5536;
 wire net5537;
 wire net5538;
 wire net5541;
 wire net5540;
 wire net5539;
 wire net5542;
 wire net5543;
 wire net5546;
 wire net5545;
 wire net5544;
 wire net5547;
 wire net5548;
 wire net5550;
 wire net5549;
 wire net5553;
 wire net5552;
 wire net5551;
 wire net5554;
 wire net5555;
 wire net5556;
 wire net5557;
 wire net5558;
 wire net5559;
 wire net5560;
 wire net5561;
 wire net5562;
 wire net5563;
 wire net5564;
 wire net5565;
 wire net5566;
 wire net5567;
 wire net5568;
 wire net5569;
 wire net5570;
 wire net5571;
 wire net5572;
 wire net5573;
 wire net5580;
 wire net5574;
 wire net5577;
 wire net5575;
 wire net5579;
 wire net5578;
 wire net5576;
 wire net5581;
 wire net5582;
 wire net5583;
 wire net5585;
 wire net5584;
 wire net5587;
 wire net5586;
 wire net5588;
 wire net5589;
 wire net5590;
 wire net5593;
 wire net5591;
 wire net5594;
 wire net5592;
 wire net5599;
 wire net5598;
 wire net5597;
 wire net5596;
 wire net5595;
 wire net5600;
 wire net5601;
 wire net5603;
 wire net5602;
 wire net5604;
 wire net5614;
 wire net5613;
 wire net5606;
 wire net5605;
 wire net5612;
 wire net5610;
 wire net5611;
 wire net5607;
 wire net5608;
 wire net5615;
 wire net5616;
 wire net5619;
 wire net5618;
 wire net5617;
 wire net5622;
 wire net5620;
 wire net5621;
 wire net5630;
 wire net5624;
 wire net5629;
 wire net5626;
 wire net5625;
 wire net5628;
 wire net5627;
 wire net5631;
 wire net5634;
 wire net5633;
 wire net5632;
 wire net5635;
 wire net5636;
 wire net5637;
 wire net5654;
 wire net5655;
 wire net5652;
 wire net5642;
 wire net5641;
 wire net5651;
 wire net5640;
 wire net5643;
 wire net5650;
 wire net5649;
 wire net5648;
 wire net5645;
 wire net5647;
 wire net5646;
 wire net5656;
 wire net5661;
 wire net5660;
 wire net5662;
 wire net5666;
 wire net5665;
 wire net5668;
 wire net5667;
 wire net5669;
 wire net5672;
 wire net5671;
 wire net5670;
 wire net5673;
 wire net5675;
 wire net5676;
 wire net5678;
 wire net5677;
 wire net5679;
 wire net5680;
 wire net5686;
 wire net5687;
 wire net5685;
 wire net5681;
 wire net5682;
 wire net5684;
 wire net5691;
 wire net5688;
 wire net5706;
 wire net5695;
 wire net5690;
 wire net5692;
 wire net5694;
 wire net5693;
 wire net5699;
 wire net5698;
 wire net5697;
 wire net5696;
 wire net5701;
 wire net5700;
 wire net5705;
 wire net5704;
 wire net5703;
 wire net5702;
 wire net5709;
 wire net5708;
 wire net5707;
 wire net5710;
 wire net5734;
 wire net5712;
 wire net5713;
 wire net5714;
 wire net5723;
 wire net5722;
 wire net5721;
 wire net5715;
 wire net5718;
 wire net5717;
 wire net5716;
 wire net5720;
 wire net5719;
 wire net5732;
 wire net5731;
 wire net5730;
 wire net5729;
 wire net5724;
 wire net5728;
 wire net5727;
 wire net5726;
 wire net5733;
 wire net5738;
 wire net5737;
 wire net5736;
 wire net5747;
 wire net5741;
 wire net5776;
 wire net5745;
 wire net5763;
 wire net5749;
 wire net5748;
 wire net5762;
 wire net5750;
 wire net5761;
 wire net5752;
 wire net5751;
 wire net5760;
 wire net5758;
 wire net5759;
 wire net5757;
 wire net5756;
 wire net5755;
 wire net5753;
 wire net5754;
 wire net5766;
 wire net5765;
 wire net5764;
 wire net5773;
 wire net5771;
 wire net5770;
 wire net5769;
 wire net5768;
 wire net5767;
 wire net5772;
 wire net5791;
 wire net5777;
 wire net5790;
 wire net5780;
 wire net5787;
 wire net5786;
 wire net5785;
 wire net5784;
 wire net5783;
 wire net5788;
 wire net5792;
 wire net5797;
 wire net5803;
 wire net5807;
 wire net5805;
 wire net5804;
 wire net5806;
 wire net5813;
 wire net5816;
 wire net5815;
 wire net5814;
 wire net5820;
 wire net5821;
 wire net5818;
 wire net5822;
 wire net5827;
 wire net5823;
 wire net5826;
 wire net5825;
 wire net5824;
 wire net5842;
 wire net5834;
 wire net5833;
 wire net5832;
 wire net5831;
 wire net5843;
 wire net5830;
 wire net5828;
 wire net5829;
 wire net5840;
 wire net5839;
 wire net5838;
 wire net5837;
 wire net5836;
 wire net5835;
 wire net5841;
 wire net5847;
 wire net5856;
 wire net5848;
 wire net5849;
 wire net5852;
 wire net5857;
 wire net5858;
 wire net5861;
 wire net5859;
 wire net5860;
 wire net5863;
 wire net5864;
 wire net5865;
 wire net5867;
 wire net5866;
 wire net5868;
 wire net5869;
 wire net5870;
 wire net5871;
 wire net5873;
 wire net5872;
 wire net5874;
 wire net5876;
 wire net5875;
 wire net5878;
 wire net5877;
 wire net5879;
 wire net5880;
 wire net5886;
 wire net5885;
 wire net5881;
 wire net5882;
 wire net5883;
 wire net5884;
 wire net5891;
 wire net5890;
 wire net5887;
 wire net5888;
 wire net5889;
 wire net5893;
 wire net5892;
 wire net5894;
 wire net5899;
 wire net5895;
 wire net5897;
 wire net5896;
 wire net5898;
 wire net5905;
 wire net5904;
 wire net5901;
 wire net5900;
 wire net5902;
 wire net5903;
 wire net5906;
 wire net5907;
 wire net5910;
 wire net5909;
 wire net5908;
 wire net5917;
 wire net5916;
 wire net5914;
 wire net5915;
 wire net5913;
 wire net5912;
 wire net5911;
 wire net5920;
 wire net5918;
 wire net5919;
 wire net5921;
 wire net5930;
 wire net5922;
 wire net5923;
 wire net5929;
 wire net5924;
 wire net5928;
 wire net5927;
 wire net5926;
 wire net5925;
 wire net5931;
 wire net5933;
 wire net5935;
 wire net5934;
 wire net5937;
 wire net5946;
 wire net5939;
 wire net5938;
 wire net5948;
 wire net5943;
 wire net5944;
 wire net5950;
 wire net5949;
 wire net5961;
 wire net5951;
 wire net5962;
 wire net5952;
 wire net5959;
 wire net5953;
 wire net5958;
 wire net5957;
 wire net5954;
 wire net5956;
 wire net5955;
 wire net5964;
 wire net5963;
 wire net5965;
 wire net5966;
 wire net5967;
 wire net5968;
 wire net5970;
 wire net5969;
 wire net5971;
 wire net5972;
 wire net5973;
 wire net5979;
 wire net5974;
 wire net5980;
 wire net5975;
 wire net5978;
 wire net5976;
 wire net5977;
 wire net5990;
 wire net5987;
 wire net5983;
 wire net5981;
 wire net5991;
 wire net5984;
 wire net5985;
 wire net5986;
 wire net5989;
 wire net5988;
 wire net6003;
 wire net5997;
 wire net5993;
 wire net5992;
 wire net5996;
 wire net5995;
 wire net5994;
 wire net5999;
 wire net5998;
 wire net6002;
 wire net6000;
 wire net6001;
 wire net6004;
 wire net6007;
 wire net6006;
 wire net6005;
 wire net6008;
 wire net6009;
 wire net6016;
 wire net6010;
 wire net6017;
 wire net6024;
 wire net6023;
 wire net6022;
 wire net6011;
 wire net6012;
 wire net6013;
 wire net6014;
 wire net6015;
 wire net6020;
 wire net6019;
 wire net6018;
 wire net6021;
 wire net6026;
 wire net6025;
 wire net6028;
 wire net6027;
 wire net6031;
 wire net6030;
 wire net6029;
 wire net6043;
 wire net6042;
 wire net6038;
 wire net6032;
 wire net6044;
 wire net6033;
 wire net6034;
 wire net6035;
 wire net6036;
 wire net6037;
 wire net6039;
 wire net6040;
 wire net6041;
 wire net6045;
 wire net6050;
 wire net6051;
 wire net6052;
 wire net6048;
 wire net6047;
 wire net6046;
 wire net6049;
 wire net6063;
 wire net6053;
 wire net6065;
 wire net6064;
 wire net6066;
 wire net6067;
 wire net6054;
 wire net6055;
 wire net6056;
 wire net6057;
 wire net6058;
 wire net6062;
 wire net6059;
 wire net6060;
 wire net6061;
 wire net6069;
 wire net6068;
 wire net6071;
 wire net6070;
 wire net6074;
 wire net6073;
 wire net6072;
 wire net6075;
 wire net6076;
 wire net6078;
 wire net6077;
 wire net6081;
 wire net6080;
 wire net6079;
 wire net6082;
 wire net6093;
 wire net6092;
 wire net6083;
 wire net6099;
 wire net6098;
 wire net6097;
 wire net6096;
 wire net6094;
 wire net6095;
 wire net6084;
 wire net6085;
 wire net6086;
 wire net6087;
 wire net6088;
 wire net6089;
 wire net6090;
 wire net6091;
 wire net6100;
 wire net6101;
 wire net6107;
 wire net6106;
 wire net6105;
 wire net6104;
 wire net6103;
 wire net6111;
 wire net6114;
 wire net6113;
 wire net6112;
 wire net6110;
 wire net6108;
 wire net6109;
 wire net6121;
 wire net6120;
 wire net6119;
 wire net6116;
 wire net6122;
 wire net6117;
 wire net6118;
 wire net6124;
 wire net6123;
 wire net6126;
 wire net6125;
 wire net6127;
 wire net6128;
 wire net6133;
 wire net6132;
 wire net6131;
 wire net6130;
 wire net6129;
 wire net6136;
 wire net6134;
 wire net6135;
 wire net6137;
 wire net6138;
 wire net6139;
 wire net6140;
 wire net6141;
 wire net6142;
 wire net6145;
 wire net6144;
 wire net6143;
 wire net6151;
 wire net6150;
 wire net6149;
 wire net6148;
 wire net6147;
 wire net6146;
 wire net6152;
 wire net6155;
 wire net6154;
 wire net6153;
 wire net6157;
 wire net6158;
 wire net6159;
 wire net6160;
 wire net6161;
 wire net6162;
 wire net6163;
 wire net6164;
 wire net6165;
 wire net6166;
 wire net6167;
 wire net6168;
 wire net6169;
 wire net6170;
 wire net6171;
 wire net6172;
 wire net6173;
 wire net6174;
 wire net6191;
 wire net6179;
 wire net6206;
 wire net6175;
 wire net6176;
 wire net6177;
 wire net6178;
 wire net6185;
 wire net6180;
 wire net6181;
 wire net6182;
 wire net6183;
 wire net6184;
 wire net6186;
 wire net6187;
 wire net6188;
 wire net6189;
 wire net6190;
 wire net6192;
 wire net6205;
 wire net6204;
 wire net6198;
 wire net6193;
 wire net6194;
 wire net6195;
 wire net6196;
 wire net6197;
 wire net6203;
 wire net6199;
 wire net6202;
 wire net6200;
 wire net6201;
 wire net6207;
 wire net6214;
 wire net6213;
 wire net6212;
 wire net6210;
 wire net6209;
 wire net6208;
 wire net6211;
 wire net6225;
 wire net6215;
 wire net6226;
 wire net6216;
 wire net6217;
 wire net6218;
 wire net6219;
 wire net6223;
 wire net6220;
 wire net6221;
 wire net6222;
 wire net6224;
 wire net6227;
 wire net6229;
 wire net6228;
 wire net6231;
 wire net6230;
 wire net6233;
 wire net6232;
 wire net6234;
 wire net6237;
 wire net6236;
 wire net6235;
 wire net6238;
 wire net6239;
 wire net6240;
 wire net6241;
 wire net6246;
 wire net6245;
 wire net6242;
 wire net6243;
 wire net6244;
 wire net6248;
 wire net6247;
 wire net6256;
 wire net6250;
 wire net6249;
 wire net6253;
 wire net6252;
 wire net6251;
 wire net6255;
 wire net6254;
 wire net6266;
 wire net6257;
 wire net6258;
 wire net6265;
 wire net6259;
 wire net6260;
 wire net6261;
 wire net6262;
 wire net6263;
 wire net6264;
 wire net6267;
 wire net6268;
 wire net6270;
 wire net6271;
 wire net6272;
 wire net6277;
 wire net6269;
 wire net6274;
 wire net6273;
 wire net6276;
 wire net6275;
 wire net6292;
 wire net6291;
 wire net6290;
 wire net6278;
 wire net6289;
 wire net6279;
 wire net6280;
 wire net6281;
 wire net6282;
 wire net6283;
 wire net6284;
 wire net6285;
 wire net6286;
 wire net6287;
 wire net6288;
 wire net6293;
 wire net6295;
 wire net6294;
 wire net6300;
 wire net6298;
 wire net6303;
 wire net6304;
 wire net6307;
 wire net6306;
 wire net6305;
 wire net6308;
 wire net6317;
 wire net6313;
 wire net6312;
 wire net6314;
 wire net6315;
 wire net6316;
 wire net6330;
 wire net6320;
 wire net6319;
 wire net6329;
 wire net6328;
 wire net6326;
 wire net6331;
 wire net6332;
 wire net6333;
 wire net6335;
 wire net6334;
 wire net6336;
 wire net6339;
 wire net6337;
 wire net6338;
 wire net6340;
 wire net6341;
 wire net6342;
 wire net6343;
 wire net6344;
 wire net6345;
 wire net6348;
 wire net6346;
 wire net6347;
 wire net6351;
 wire net6349;
 wire net6350;
 wire net6352;
 wire net6373;
 wire net6353;
 wire net6354;
 wire net6372;
 wire net6355;
 wire net6356;
 wire net6363;
 wire net6357;
 wire net6358;
 wire net6359;
 wire net6360;
 wire net6361;
 wire net6362;
 wire net6364;
 wire net6365;
 wire net6366;
 wire net6371;
 wire net6367;
 wire net6368;
 wire net6370;
 wire net6369;
 wire net6379;
 wire net6378;
 wire net6377;
 wire net6376;
 wire net6375;
 wire net6374;
 wire net6380;
 wire net6381;
 wire net6383;
 wire net6385;
 wire net6384;
 wire net6386;
 wire net6387;
 wire net6388;
 wire net6389;
 wire net6390;
 wire net6392;
 wire net6391;
 wire net6393;
 wire net6394;
 wire net6395;
 wire net6397;
 wire net6396;
 wire net6398;
 wire net6399;
 wire net6400;
 wire net6401;
 wire net6402;
 wire net6403;
 wire net6404;
 wire net6405;
 wire net6406;
 wire net6407;
 wire net6409;
 wire net6408;
 wire net6410;
 wire net6411;
 wire net6412;
 wire net6413;
 wire net6414;
 wire net6415;
 wire net6418;
 wire net6416;
 wire net6417;
 wire net6419;
 wire net6420;
 wire net6421;
 wire net6422;
 wire net6423;
 wire net6424;
 wire net6425;
 wire net6426;
 wire net6427;
 wire net6430;
 wire net6428;
 wire net6429;
 wire net6431;
 wire net6432;
 wire net6433;
 wire net6434;
 wire net6435;
 wire net6436;
 wire net6437;
 wire net6438;
 wire net6439;
 wire net6440;
 wire net6441;
 wire net6442;
 wire net6464;
 wire net6463;
 wire net6443;
 wire net6444;
 wire net6445;
 wire net6462;
 wire net6461;
 wire net6460;
 wire net6459;
 wire net6458;
 wire net6457;
 wire net6456;
 wire net6455;
 wire net6453;
 wire net6446;
 wire net6447;
 wire net6448;
 wire net6451;
 wire net6449;
 wire net6450;
 wire net6452;
 wire net6454;
 wire net6466;
 wire net6467;
 wire net6468;
 wire net6469;
 wire net6470;
 wire net6471;
 wire net6472;
 wire net6473;
 wire net6474;
 wire net6475;
 wire net6476;
 wire net6477;
 wire net6478;
 wire net6479;
 wire net6480;
 wire net6481;
 wire net6482;
 wire net6483;
 wire net6484;
 wire net6485;
 wire net6486;
 wire net6487;
 wire net6488;
 wire net6489;
 wire net6490;
 wire net6491;
 wire net6492;
 wire net6493;
 wire net6494;
 wire net6495;
 wire net6496;
 wire net6497;
 wire net6498;
 wire net6499;
 wire net6500;
 wire net6501;
 wire net6502;
 wire net6503;
 wire net6504;
 wire net6505;
 wire net6506;
 wire net6507;
 wire net6508;
 wire net6510;
 wire net6509;
 wire net6511;
 wire net6512;
 wire net6513;
 wire net6514;
 wire net6515;
 wire net6516;
 wire net6517;
 wire net6518;
 wire net6519;
 wire net6520;
 wire net6521;
 wire net6522;
 wire net6523;
 wire net6524;
 wire net6525;
 wire net6526;
 wire net6527;
 wire net6528;
 wire net6529;
 wire net6530;
 wire net6531;
 wire net6532;
 wire net6533;
 wire net6537;
 wire net6534;
 wire net6535;
 wire net6536;
 wire net6538;
 wire net6539;
 wire net6540;
 wire net6541;
 wire net6542;
 wire net6543;
 wire net6544;
 wire net6546;
 wire net6545;
 wire net6547;
 wire net6548;
 wire net6549;
 wire net6550;
 wire net6551;
 wire net6552;
 wire net6553;
 wire net6554;
 wire net6555;
 wire net6556;
 wire net6557;
 wire net6558;
 wire net6559;
 wire net6560;
 wire net6561;
 wire net6562;
 wire net6563;
 wire net6569;
 wire net6564;
 wire net6567;
 wire net6565;
 wire net6568;
 wire net6566;
 wire net6571;
 wire net6570;
 wire net6572;
 wire net6573;
 wire net6580;
 wire net6574;
 wire net6577;
 wire net6575;
 wire net6579;
 wire net6576;
 wire net6578;
 wire net6581;
 wire net6583;
 wire net6582;
 wire net6586;
 wire net6584;
 wire net6593;
 wire net6585;
 wire net6587;
 wire net6588;
 wire net6591;
 wire net6589;
 wire net6590;
 wire net6592;
 wire net6594;
 wire net6595;
 wire net6596;
 wire net6597;
 wire net6601;
 wire net6599;
 wire net6598;
 wire net6600;
 wire clknet_2_2_0_clk;
 wire clknet_2_3_0_clk;
 wire net6602;
 wire clknet_2_1_0_clk;
 wire net6606;
 wire net6605;
 wire net6603;
 wire net6604;
 wire clknet_0_clk;
 wire net6607;
 wire clknet_2_0_0_clk;
 wire clknet_leaf_34_clk;
 wire net6608;
 wire net6609;
 wire net6610;
 wire clknet_leaf_33_clk;
 wire net6611;
 wire net6613;
 wire net6612;
 wire net6614;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_31_clk;
 wire net6673;
 wire net6672;
 wire net6618;
 wire net6615;
 wire net6616;
 wire net6617;
 wire net6670;
 wire net6669;
 wire net6671;
 wire net6668;
 wire net6623;
 wire net6619;
 wire net6620;
 wire net6621;
 wire net6622;
 wire net6624;
 wire net6667;
 wire net6666;
 wire net6665;
 wire net6625;
 wire net6627;
 wire net6626;
 wire net6631;
 wire net6628;
 wire net6630;
 wire net6629;
 wire net6639;
 wire net6664;
 wire net6632;
 wire net6633;
 wire net6634;
 wire net6635;
 wire net6636;
 wire net6638;
 wire net6637;
 wire net6663;
 wire net6640;
 wire net6662;
 wire net6661;
 wire net6660;
 wire net6659;
 wire net6658;
 wire net6641;
 wire net6644;
 wire net6642;
 wire net6643;
 wire net6656;
 wire net6657;
 wire net6649;
 wire net6645;
 wire net6646;
 wire net6648;
 wire net6647;
 wire net6651;
 wire net6650;
 wire net6652;
 wire net6654;
 wire net6653;
 wire net6655;
 wire net6677;
 wire net6676;
 wire net6675;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_12_clk;
 wire net6679;
 wire net6678;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_27_clk;
 wire net6681;
 wire net6682;
 wire net6690;
 wire net6689;
 wire net6687;
 wire net6686;
 wire net6688;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_9_clk;
 wire net4454;
 wire net4457;

 XOR2x2_ASAP7_75t_R _15840_ (.A(net6548),
    .B(net6477),
    .Y(_00265_));
 XOR2x2_ASAP7_75t_R _15842_ (.A(net6545),
    .B(net6473),
    .Y(_00266_));
 XOR2x2_ASAP7_75t_R _15844_ (.A(net6544),
    .B(_00956_),
    .Y(_00267_));
 XOR2x2_ASAP7_75t_R _15845_ (.A(_00698_),
    .B(_00959_),
    .Y(_00268_));
 XOR2x2_ASAP7_75t_R _15846_ (.A(net6543),
    .B(_00960_),
    .Y(_00269_));
 XOR2x2_ASAP7_75t_R _15848_ (.A(_00700_),
    .B(_00961_),
    .Y(_00270_));
 XOR2x2_ASAP7_75t_R _15849_ (.A(_00701_),
    .B(_00962_),
    .Y(_00271_));
 XOR2x2_ASAP7_75t_R _15851_ (.A(net6542),
    .B(_00963_),
    .Y(_00272_));
 XOR2x2_ASAP7_75t_R _15854_ (.A(net6553),
    .B(net6492),
    .Y(_00217_));
 XOR2x2_ASAP7_75t_R _15857_ (.A(net6552),
    .B(net6487),
    .Y(_00218_));
 XOR2x2_ASAP7_75t_R _15859_ (.A(net6551),
    .B(net6480),
    .Y(_00219_));
 XOR2x2_ASAP7_75t_R _15860_ (.A(net6550),
    .B(_00927_),
    .Y(_00220_));
 XOR2x2_ASAP7_75t_R _15861_ (.A(_00691_),
    .B(_00928_),
    .Y(_00221_));
 XOR2x2_ASAP7_75t_R _15863_ (.A(_00692_),
    .B(_00929_),
    .Y(_00222_));
 XOR2x2_ASAP7_75t_R _15864_ (.A(_00693_),
    .B(_00930_),
    .Y(_00223_));
 XOR2x2_ASAP7_75t_R _15866_ (.A(net6549),
    .B(_00931_),
    .Y(_00224_));
 XOR2x2_ASAP7_75t_R _15868_ (.A(net6559),
    .B(net6512),
    .Y(_00249_));
 XOR2x2_ASAP7_75t_R _15871_ (.A(net6558),
    .B(net6505),
    .Y(_00250_));
 XOR2x2_ASAP7_75t_R _15873_ (.A(_00681_),
    .B(net6499),
    .Y(_00251_));
 XOR2x2_ASAP7_75t_R _15874_ (.A(_00682_),
    .B(net6498),
    .Y(_00252_));
 XOR2x2_ASAP7_75t_R _15875_ (.A(net6556),
    .B(net6497),
    .Y(_00253_));
 XOR2x2_ASAP7_75t_R _15876_ (.A(net6555),
    .B(net6496),
    .Y(_00254_));
 XOR2x2_ASAP7_75t_R _15877_ (.A(_00685_),
    .B(net6495),
    .Y(_00255_));
 XOR2x2_ASAP7_75t_R _15879_ (.A(net6554),
    .B(_00899_),
    .Y(_00256_));
 XOR2x2_ASAP7_75t_R _15882_ (.A(net6566),
    .B(net6539),
    .Y(_00161_));
 XOR2x2_ASAP7_75t_R _15884_ (.A(net6565),
    .B(net6529),
    .Y(_00162_));
 XOR2x2_ASAP7_75t_R _15887_ (.A(net6564),
    .B(net6522),
    .Y(_00163_));
 XOR2x2_ASAP7_75t_R _15888_ (.A(net6563),
    .B(net6519),
    .Y(_00164_));
 XOR2x2_ASAP7_75t_R _15889_ (.A(net6562),
    .B(net6518),
    .Y(_00165_));
 XOR2x2_ASAP7_75t_R _15891_ (.A(net6561),
    .B(net6517),
    .Y(_00166_));
 XOR2x2_ASAP7_75t_R _15892_ (.A(_00677_),
    .B(net6516),
    .Y(_00167_));
 XOR2x2_ASAP7_75t_R _15894_ (.A(net6560),
    .B(net6515),
    .Y(_00168_));
 XOR2x2_ASAP7_75t_R _15895_ (.A(net6576),
    .B(_00964_),
    .Y(_00193_));
 XOR2x2_ASAP7_75t_R _15897_ (.A(net6472),
    .B(net6575),
    .Y(_00194_));
 XOR2x2_ASAP7_75t_R _15900_ (.A(net6574),
    .B(net6476),
    .Y(_00195_));
 XOR2x2_ASAP7_75t_R _15902_ (.A(net6573),
    .B(_00936_),
    .Y(_00196_));
 XOR2x2_ASAP7_75t_R _15903_ (.A(net6572),
    .B(_00937_),
    .Y(_00197_));
 XOR2x2_ASAP7_75t_R _15904_ (.A(_00668_),
    .B(_00938_),
    .Y(_00198_));
 XOR2x2_ASAP7_75t_R _15905_ (.A(_00669_),
    .B(_00939_),
    .Y(_00199_));
 XOR2x2_ASAP7_75t_R _15907_ (.A(net6570),
    .B(_00940_),
    .Y(_00200_));
 XOR2x2_ASAP7_75t_R _15909_ (.A(net6586),
    .B(net6479),
    .Y(_00225_));
 XOR2x2_ASAP7_75t_R _15911_ (.A(net6584),
    .B(net6478),
    .Y(_00226_));
 XOR2x2_ASAP7_75t_R _15914_ (.A(net6582),
    .B(net6491),
    .Y(_00227_));
 XOR2x2_ASAP7_75t_R _15917_ (.A(net6581),
    .B(net6490),
    .Y(_00228_));
 XOR2x2_ASAP7_75t_R _15918_ (.A(_00659_),
    .B(_00905_),
    .Y(_00229_));
 XOR2x2_ASAP7_75t_R _15919_ (.A(_00660_),
    .B(_00906_),
    .Y(_00230_));
 XOR2x2_ASAP7_75t_R _15920_ (.A(_00661_),
    .B(_00907_),
    .Y(_00231_));
 XOR2x2_ASAP7_75t_R _15922_ (.A(net6578),
    .B(_00908_),
    .Y(_00232_));
 XOR2x2_ASAP7_75t_R _15924_ (.A(_00647_),
    .B(net6494),
    .Y(_00257_));
 XOR2x2_ASAP7_75t_R _15925_ (.A(net6590),
    .B(net6493),
    .Y(_00258_));
 XOR2x2_ASAP7_75t_R _15928_ (.A(net6589),
    .B(net6511),
    .Y(_00259_));
 XOR2x2_ASAP7_75t_R _15929_ (.A(_00650_),
    .B(net6510),
    .Y(_00260_));
 XOR2x2_ASAP7_75t_R _15930_ (.A(_00651_),
    .B(net6509),
    .Y(_00261_));
 XOR2x2_ASAP7_75t_R _15931_ (.A(net6588),
    .B(_00874_),
    .Y(_00262_));
 XOR2x2_ASAP7_75t_R _15932_ (.A(_00653_),
    .B(_00875_),
    .Y(_00263_));
 XOR2x2_ASAP7_75t_R _15934_ (.A(net6587),
    .B(_00876_),
    .Y(_00264_));
 XOR2x2_ASAP7_75t_R _15935_ (.A(net6599),
    .B(net6514),
    .Y(_00169_));
 XOR2x2_ASAP7_75t_R _15937_ (.A(net6597),
    .B(net6513),
    .Y(_00170_));
 XOR2x2_ASAP7_75t_R _15940_ (.A(net6596),
    .B(net6538),
    .Y(_00171_));
 XOR2x2_ASAP7_75t_R _15942_ (.A(net6595),
    .B(net6537),
    .Y(_00172_));
 XOR2x2_ASAP7_75t_R _15943_ (.A(_00643_),
    .B(net6536),
    .Y(_00173_));
 XOR2x2_ASAP7_75t_R _15944_ (.A(net6594),
    .B(net6535),
    .Y(_00174_));
 XOR2x2_ASAP7_75t_R _15945_ (.A(_00645_),
    .B(net6534),
    .Y(_00175_));
 XOR2x2_ASAP7_75t_R _15947_ (.A(net6593),
    .B(_00844_),
    .Y(_00176_));
 XOR2x2_ASAP7_75t_R _15948_ (.A(net6603),
    .B(net6475),
    .Y(_00201_));
 XOR2x2_ASAP7_75t_R _15949_ (.A(_00632_),
    .B(net6474),
    .Y(_00202_));
 XOR2x2_ASAP7_75t_R _15952_ (.A(net6602),
    .B(_00943_),
    .Y(_00203_));
 XOR2x2_ASAP7_75t_R _15953_ (.A(_00634_),
    .B(_00944_),
    .Y(_00204_));
 XOR2x2_ASAP7_75t_R _15954_ (.A(_00635_),
    .B(_00946_),
    .Y(_00205_));
 XOR2x2_ASAP7_75t_R _15955_ (.A(_00636_),
    .B(_00947_),
    .Y(_00206_));
 XOR2x2_ASAP7_75t_R _15956_ (.A(_00637_),
    .B(_00948_),
    .Y(_00207_));
 XOR2x2_ASAP7_75t_R _15958_ (.A(net6600),
    .B(_00949_),
    .Y(_00208_));
 XOR2x2_ASAP7_75t_R _15960_ (.A(net6612),
    .B(net6489),
    .Y(_00233_));
 XOR2x2_ASAP7_75t_R _15962_ (.A(net6611),
    .B(net6488),
    .Y(_00234_));
 XOR2x2_ASAP7_75t_R _15965_ (.A(net6610),
    .B(_00911_),
    .Y(_00235_));
 XOR2x2_ASAP7_75t_R _15968_ (.A(net6609),
    .B(_00912_),
    .Y(_00236_));
 XOR2x2_ASAP7_75t_R _15970_ (.A(net6608),
    .B(net6486),
    .Y(_00237_));
 XOR2x2_ASAP7_75t_R _15972_ (.A(_00628_),
    .B(_00915_),
    .Y(_00238_));
 XOR2x2_ASAP7_75t_R _15973_ (.A(net6607),
    .B(_00916_),
    .Y(_00239_));
 XOR2x2_ASAP7_75t_R _15975_ (.A(net6604),
    .B(net6485),
    .Y(_00240_));
 XOR2x2_ASAP7_75t_R _15976_ (.A(net6616),
    .B(net6508),
    .Y(_00273_));
 XOR2x2_ASAP7_75t_R _15977_ (.A(net6615),
    .B(net6507),
    .Y(_00274_));
 XOR2x2_ASAP7_75t_R _15980_ (.A(_00617_),
    .B(net6506),
    .Y(_00275_));
 XOR2x2_ASAP7_75t_R _15981_ (.A(_00618_),
    .B(_00880_),
    .Y(_00276_));
 XOR2x2_ASAP7_75t_R _15983_ (.A(_00619_),
    .B(_00882_),
    .Y(_00277_));
 XOR2x2_ASAP7_75t_R _15984_ (.A(_00620_),
    .B(_00883_),
    .Y(_00278_));
 XOR2x2_ASAP7_75t_R _15985_ (.A(_00621_),
    .B(_00884_),
    .Y(_00279_));
 XOR2x2_ASAP7_75t_R _15987_ (.A(net6614),
    .B(net6504),
    .Y(_00280_));
 XOR2x2_ASAP7_75t_R _15989_ (.A(net6622),
    .B(net6533),
    .Y(_00177_));
 XOR2x2_ASAP7_75t_R _15990_ (.A(net6621),
    .B(net6532),
    .Y(_00178_));
 XOR2x2_ASAP7_75t_R _15993_ (.A(_00609_),
    .B(net6531),
    .Y(_00179_));
 XOR2x2_ASAP7_75t_R _15994_ (.A(net6619),
    .B(net6530),
    .Y(_00180_));
 XOR2x2_ASAP7_75t_R _15995_ (.A(_00611_),
    .B(_00850_),
    .Y(_00181_));
 XOR2x2_ASAP7_75t_R _15996_ (.A(_00612_),
    .B(_00851_),
    .Y(_00182_));
 XOR2x2_ASAP7_75t_R _15997_ (.A(_00613_),
    .B(_00852_),
    .Y(_00183_));
 XOR2x2_ASAP7_75t_R _15999_ (.A(net6617),
    .B(_00853_),
    .Y(_00184_));
 XOR2x2_ASAP7_75t_R _16001_ (.A(net6628),
    .B(_00950_),
    .Y(_00209_));
 XOR2x2_ASAP7_75t_R _16003_ (.A(net6626),
    .B(_00951_),
    .Y(_00210_));
 XOR2x2_ASAP7_75t_R _16005_ (.A(net6625),
    .B(_00952_),
    .Y(_00211_));
 XOR2x2_ASAP7_75t_R _16006_ (.A(_00602_),
    .B(_00953_),
    .Y(_00212_));
 XOR2x2_ASAP7_75t_R _16007_ (.A(_00603_),
    .B(_00954_),
    .Y(_00213_));
 XOR2x2_ASAP7_75t_R _16008_ (.A(_00604_),
    .B(_00955_),
    .Y(_00214_));
 XOR2x2_ASAP7_75t_R _16009_ (.A(_00605_),
    .B(_00957_),
    .Y(_00215_));
 XOR2x2_ASAP7_75t_R _16011_ (.A(net6624),
    .B(_00958_),
    .Y(_00216_));
 XOR2x2_ASAP7_75t_R _16013_ (.A(net6637),
    .B(net6484),
    .Y(_00241_));
 XOR2x2_ASAP7_75t_R _16016_ (.A(net6635),
    .B(net6483),
    .Y(_00242_));
 XOR2x2_ASAP7_75t_R _16019_ (.A(net6634),
    .B(net6482),
    .Y(_00243_));
 XOR2x2_ASAP7_75t_R _16020_ (.A(net6633),
    .B(net6481),
    .Y(_00244_));
 XOR2x2_ASAP7_75t_R _16021_ (.A(_00595_),
    .B(_00922_),
    .Y(_00245_));
 XOR2x2_ASAP7_75t_R _16022_ (.A(net6632),
    .B(_00923_),
    .Y(_00246_));
 XOR2x2_ASAP7_75t_R _16023_ (.A(_00597_),
    .B(_00925_),
    .Y(_00247_));
 XOR2x2_ASAP7_75t_R _16025_ (.A(net6629),
    .B(_00926_),
    .Y(_00248_));
 XOR2x2_ASAP7_75t_R _16027_ (.A(net6642),
    .B(net6503),
    .Y(_00281_));
 XOR2x2_ASAP7_75t_R _16030_ (.A(_00584_),
    .B(net6502),
    .Y(_00282_));
 XOR2x2_ASAP7_75t_R _16033_ (.A(_00585_),
    .B(net6501),
    .Y(_00283_));
 XOR2x2_ASAP7_75t_R _16034_ (.A(_00586_),
    .B(net6500),
    .Y(_00284_));
 XOR2x2_ASAP7_75t_R _16035_ (.A(_00587_),
    .B(_00890_),
    .Y(_00285_));
 XOR2x2_ASAP7_75t_R _16036_ (.A(_00588_),
    .B(_00891_),
    .Y(_00286_));
 XOR2x2_ASAP7_75t_R _16037_ (.A(_00589_),
    .B(_00893_),
    .Y(_00287_));
 XOR2x2_ASAP7_75t_R _16039_ (.A(net6640),
    .B(_00894_),
    .Y(_00288_));
 XOR2x2_ASAP7_75t_R _16041_ (.A(net6652),
    .B(net6528),
    .Y(_00185_));
 XOR2x2_ASAP7_75t_R _16044_ (.A(net6648),
    .B(net6527),
    .Y(_00186_));
 XOR2x2_ASAP7_75t_R _16047_ (.A(_00577_),
    .B(net6526),
    .Y(_00187_));
 XOR2x2_ASAP7_75t_R _16048_ (.A(net6645),
    .B(net6525),
    .Y(_00188_));
 XOR2x2_ASAP7_75t_R _16049_ (.A(_00579_),
    .B(net6524),
    .Y(_00189_));
 XOR2x2_ASAP7_75t_R _16050_ (.A(_00580_),
    .B(net6523),
    .Y(_00190_));
 XOR2x2_ASAP7_75t_R _16051_ (.A(_00581_),
    .B(net6521),
    .Y(_00191_));
 XOR2x2_ASAP7_75t_R _16053_ (.A(net6643),
    .B(net6520),
    .Y(_00192_));
 INVx8_ASAP7_75t_R _16055_ (.A(net6685),
    .Y(_08030_));
 INVx1_ASAP7_75t_R _16060_ (.A(_00572_),
    .Y(_08035_));
 AND5x1_ASAP7_75t_R _16061_ (.A(_00411_),
    .B(net6678),
    .C(_08035_),
    .D(_00570_),
    .E(_00571_),
    .Y(_00160_));
 INVx1_ASAP7_75t_R _16062_ (.A(_00965_),
    .Y(\u0.r0.rcnt[1] ));
 INVx1_ASAP7_75t_R _16063_ (.A(\u0.r0.rcnt_next[0] ),
    .Y(\u0.r0.rcnt[0] ));
 XOR2x2_ASAP7_75t_R _16065_ (.A(_00439_),
    .B(_00912_),
    .Y(_08037_));
 INVx1_ASAP7_75t_R _16066_ (.A(_00944_),
    .Y(_08038_));
 XOR2x2_ASAP7_75t_R _16067_ (.A(_08037_),
    .B(_08038_),
    .Y(_08039_));
 XNOR2x2_ASAP7_75t_R _16068_ (.A(_00848_),
    .B(_00880_),
    .Y(_08040_));
 XOR2x2_ASAP7_75t_R _16069_ (.A(_08039_),
    .B(_08040_),
    .Y(_08041_));
 NOR2x1_ASAP7_75t_R _16070_ (.A(net39),
    .B(net6679),
    .Y(_08042_));
 AOI21x1_ASAP7_75t_R _16071_ (.A1(net6679),
    .A2(_08041_),
    .B(_08042_),
    .Y(_08043_));
 XOR2x2_ASAP7_75t_R _16074_ (.A(_00437_),
    .B(_00909_),
    .Y(_08045_));
 INVx1_ASAP7_75t_R _16075_ (.A(_00941_),
    .Y(_08046_));
 XOR2x2_ASAP7_75t_R _16076_ (.A(_08045_),
    .B(_08046_),
    .Y(_08047_));
 XNOR2x2_ASAP7_75t_R _16077_ (.A(_00845_),
    .B(_00877_),
    .Y(_08048_));
 XOR2x2_ASAP7_75t_R _16078_ (.A(_08047_),
    .B(_08048_),
    .Y(_08049_));
 NAND2x1_ASAP7_75t_R _16079_ (.A(_08030_),
    .B(_08049_),
    .Y(_08050_));
 OAI21x1_ASAP7_75t_R _16080_ (.A1(_08030_),
    .A2(net36),
    .B(_08050_),
    .Y(_08051_));
 XOR2x2_ASAP7_75t_R _16082_ (.A(_00412_),
    .B(_00847_),
    .Y(_08052_));
 XOR2x2_ASAP7_75t_R _16083_ (.A(_00879_),
    .B(_00911_),
    .Y(_08053_));
 XOR2x2_ASAP7_75t_R _16084_ (.A(_08052_),
    .B(_08053_),
    .Y(_08054_));
 XOR2x2_ASAP7_75t_R _16085_ (.A(_08054_),
    .B(_00943_),
    .Y(_08055_));
 AND2x2_ASAP7_75t_R _16086_ (.A(net6687),
    .B(net38),
    .Y(_08056_));
 INVx1_ASAP7_75t_R _16087_ (.A(_08056_),
    .Y(_08057_));
 OA21x2_ASAP7_75t_R _16088_ (.A1(_08055_),
    .A2(net6689),
    .B(_08057_),
    .Y(_08058_));
 INVx1_ASAP7_75t_R _16090_ (.A(_08058_),
    .Y(_08060_));
 XOR2x2_ASAP7_75t_R _16093_ (.A(_00438_),
    .B(_00910_),
    .Y(_08062_));
 INVx1_ASAP7_75t_R _16094_ (.A(_00942_),
    .Y(_08063_));
 XOR2x2_ASAP7_75t_R _16095_ (.A(_08062_),
    .B(_08063_),
    .Y(_08064_));
 XNOR2x2_ASAP7_75t_R _16096_ (.A(_00846_),
    .B(_00878_),
    .Y(_08065_));
 XOR2x2_ASAP7_75t_R _16097_ (.A(_08064_),
    .B(_08065_),
    .Y(_08066_));
 NAND2x1p5_ASAP7_75t_R _16098_ (.A(_08030_),
    .B(_08066_),
    .Y(_08067_));
 OAI21x1_ASAP7_75t_R _16099_ (.A1(net37),
    .A2(_08030_),
    .B(_08067_),
    .Y(_00980_));
 XOR2x2_ASAP7_75t_R _16100_ (.A(_00440_),
    .B(_00914_),
    .Y(_08068_));
 INVx1_ASAP7_75t_R _16101_ (.A(_00946_),
    .Y(_08069_));
 XOR2x2_ASAP7_75t_R _16102_ (.A(_08068_),
    .B(_08069_),
    .Y(_08070_));
 XNOR2x2_ASAP7_75t_R _16103_ (.A(_00850_),
    .B(_00882_),
    .Y(_08071_));
 XOR2x2_ASAP7_75t_R _16104_ (.A(_08070_),
    .B(_08071_),
    .Y(_08072_));
 NAND2x1_ASAP7_75t_R _16105_ (.A(net6677),
    .B(_08072_),
    .Y(_08073_));
 OA21x2_ASAP7_75t_R _16106_ (.A1(net6677),
    .A2(net41),
    .B(_08073_),
    .Y(_08074_));
 XOR2x2_ASAP7_75t_R _16110_ (.A(_00441_),
    .B(_00915_),
    .Y(_08077_));
 XNOR2x2_ASAP7_75t_R _16111_ (.A(_00947_),
    .B(_08077_),
    .Y(_08078_));
 XNOR2x2_ASAP7_75t_R _16112_ (.A(_00851_),
    .B(_00883_),
    .Y(_08079_));
 XOR2x2_ASAP7_75t_R _16113_ (.A(_08078_),
    .B(_08079_),
    .Y(_08080_));
 NAND2x1_ASAP7_75t_R _16114_ (.A(net6678),
    .B(_08080_),
    .Y(_08081_));
 OA21x2_ASAP7_75t_R _16115_ (.A1(net6678),
    .A2(net42),
    .B(_08081_),
    .Y(_08082_));
 XOR2x2_ASAP7_75t_R _16119_ (.A(_00442_),
    .B(_00916_),
    .Y(_08085_));
 XNOR2x2_ASAP7_75t_R _16120_ (.A(_00948_),
    .B(_08085_),
    .Y(_08086_));
 XNOR2x2_ASAP7_75t_R _16121_ (.A(_00852_),
    .B(_00884_),
    .Y(_08087_));
 XOR2x2_ASAP7_75t_R _16122_ (.A(_08086_),
    .B(_08087_),
    .Y(_08088_));
 NAND2x1_ASAP7_75t_R _16123_ (.A(net6677),
    .B(_08088_),
    .Y(_08089_));
 OA21x2_ASAP7_75t_R _16124_ (.A1(net6677),
    .A2(net43),
    .B(_08089_),
    .Y(_08090_));
 XOR2x2_ASAP7_75t_R _16127_ (.A(_00443_),
    .B(_00917_),
    .Y(_08092_));
 XNOR2x2_ASAP7_75t_R _16128_ (.A(_00949_),
    .B(_08092_),
    .Y(_08093_));
 XNOR2x2_ASAP7_75t_R _16129_ (.A(_00853_),
    .B(net6504),
    .Y(_08094_));
 XOR2x2_ASAP7_75t_R _16130_ (.A(_08093_),
    .B(_08094_),
    .Y(_08095_));
 NAND2x1_ASAP7_75t_R _16131_ (.A(net6678),
    .B(_08095_),
    .Y(_08096_));
 OA21x2_ASAP7_75t_R _16132_ (.A1(net6678),
    .A2(net44),
    .B(_08096_),
    .Y(_08097_));
 INVx3_ASAP7_75t_R _16134_ (.A(_00980_),
    .Y(_00972_));
 INVx2_ASAP7_75t_R _16137_ (.A(_08051_),
    .Y(_00973_));
 NOR2x1_ASAP7_75t_R _16138_ (.A(_00979_),
    .B(_08043_),
    .Y(_08099_));
 AND2x2_ASAP7_75t_R _16139_ (.A(_08099_),
    .B(net6372),
    .Y(_08100_));
 INVx1_ASAP7_75t_R _16140_ (.A(net4985),
    .Y(_08101_));
 NAND2x1_ASAP7_75t_R _16141_ (.A(net6378),
    .B(net6369),
    .Y(_08102_));
 NOR2x1_ASAP7_75t_R _16142_ (.A(net6340),
    .B(_08102_),
    .Y(_08103_));
 INVx1_ASAP7_75t_R _16143_ (.A(_00974_),
    .Y(_08104_));
 NOR2x1_ASAP7_75t_R _16144_ (.A(_08104_),
    .B(net6369),
    .Y(_08105_));
 AO21x1_ASAP7_75t_R _16146_ (.A1(_08105_),
    .A2(net6378),
    .B(net6336),
    .Y(_08107_));
 NOR2x1_ASAP7_75t_R _16147_ (.A(_08103_),
    .B(_08107_),
    .Y(_08108_));
 AOI21x1_ASAP7_75t_R _16149_ (.A1(_08101_),
    .A2(_08108_),
    .B(net6333),
    .Y(_08110_));
 INVx2_ASAP7_75t_R _16150_ (.A(_08043_),
    .Y(_08111_));
 INVx1_ASAP7_75t_R _16151_ (.A(_00975_),
    .Y(_08112_));
 NOR2x1p5_ASAP7_75t_R _16152_ (.A(net6369),
    .B(_08112_),
    .Y(_08113_));
 NOR2x1p5_ASAP7_75t_R _16153_ (.A(net6327),
    .B(_08113_),
    .Y(_08114_));
 NOR2x1_ASAP7_75t_R _16154_ (.A(_00982_),
    .B(net6369),
    .Y(_08115_));
 NAND2x1_ASAP7_75t_R _16155_ (.A(net6327),
    .B(net5251),
    .Y(_08116_));
 INVx2_ASAP7_75t_R _16156_ (.A(_08074_),
    .Y(_08117_));
 NOR2x1_ASAP7_75t_R _16157_ (.A(_08117_),
    .B(_08100_),
    .Y(_08118_));
 NAND2x1_ASAP7_75t_R _16158_ (.A(_08116_),
    .B(_08118_),
    .Y(_08119_));
 OR2x2_ASAP7_75t_R _16159_ (.A(_08114_),
    .B(_08119_),
    .Y(_08120_));
 INVx1_ASAP7_75t_R _16160_ (.A(_08090_),
    .Y(_08121_));
 AOI21x1_ASAP7_75t_R _16161_ (.A1(_08110_),
    .A2(_08120_),
    .B(net5975),
    .Y(_08122_));
 NAND2x1p5_ASAP7_75t_R _16163_ (.A(net6369),
    .B(net5029),
    .Y(_08124_));
 NOR2x1_ASAP7_75t_R _16166_ (.A(net6373),
    .B(net6337),
    .Y(_08127_));
 NOR2x1_ASAP7_75t_R _16167_ (.A(net6378),
    .B(_08127_),
    .Y(_08128_));
 NAND2x1_ASAP7_75t_R _16168_ (.A(net4790),
    .B(_08128_),
    .Y(_08129_));
 NOR2x1_ASAP7_75t_R _16169_ (.A(net6372),
    .B(net6340),
    .Y(_08130_));
 INVx1_ASAP7_75t_R _16170_ (.A(_08130_),
    .Y(_08131_));
 NAND2x1_ASAP7_75t_R _16171_ (.A(_00981_),
    .B(net6369),
    .Y(_08132_));
 AO21x1_ASAP7_75t_R _16173_ (.A1(_08131_),
    .A2(net5250),
    .B(net6329),
    .Y(_08134_));
 AOI21x1_ASAP7_75t_R _16175_ (.A1(_08129_),
    .A2(_08134_),
    .B(net6335),
    .Y(_08136_));
 NOR2x1_ASAP7_75t_R _16176_ (.A(_00984_),
    .B(net6373),
    .Y(_08137_));
 INVx1_ASAP7_75t_R _16177_ (.A(_08137_),
    .Y(_08138_));
 NAND2x1_ASAP7_75t_R _16178_ (.A(_00983_),
    .B(net6373),
    .Y(_08139_));
 AO21x1_ASAP7_75t_R _16179_ (.A1(_08138_),
    .A2(_08139_),
    .B(net6376),
    .Y(_08140_));
 INVx1_ASAP7_75t_R _16180_ (.A(_08140_),
    .Y(_08141_));
 INVx1_ASAP7_75t_R _16182_ (.A(_00979_),
    .Y(_08143_));
 OA21x2_ASAP7_75t_R _16183_ (.A1(net6371),
    .A2(net5249),
    .B(net6378),
    .Y(_08144_));
 OA21x2_ASAP7_75t_R _16184_ (.A1(_08141_),
    .A2(_08144_),
    .B(net6335),
    .Y(_08145_));
 OAI21x1_ASAP7_75t_R _16186_ (.A1(_08136_),
    .A2(_08145_),
    .B(net6333),
    .Y(_08147_));
 NAND2x1_ASAP7_75t_R _16187_ (.A(_08122_),
    .B(_08147_),
    .Y(_08148_));
 NAND2x1_ASAP7_75t_R _16189_ (.A(net6376),
    .B(net5561),
    .Y(_08150_));
 NAND2x1_ASAP7_75t_R _16190_ (.A(net5321),
    .B(net6339),
    .Y(_08151_));
 AO21x1_ASAP7_75t_R _16192_ (.A1(net5248),
    .A2(net5250),
    .B(net6376),
    .Y(_08153_));
 AOI21x1_ASAP7_75t_R _16195_ (.A1(_08150_),
    .A2(_08153_),
    .B(net5980),
    .Y(_08156_));
 NOR2x1_ASAP7_75t_R _16196_ (.A(net5321),
    .B(net6372),
    .Y(_08157_));
 AO21x1_ASAP7_75t_R _16197_ (.A1(net6373),
    .A2(_00982_),
    .B(net6330),
    .Y(_08158_));
 NOR2x1_ASAP7_75t_R _16198_ (.A(net5247),
    .B(_08158_),
    .Y(_08159_));
 NOR2x1_ASAP7_75t_R _16200_ (.A(net6376),
    .B(_08138_),
    .Y(_08161_));
 OA21x2_ASAP7_75t_R _16202_ (.A1(_08159_),
    .A2(_08161_),
    .B(net5980),
    .Y(_08163_));
 OAI21x1_ASAP7_75t_R _16203_ (.A1(_08156_),
    .A2(_08163_),
    .B(net6333),
    .Y(_08164_));
 NOR2x1_ASAP7_75t_R _16204_ (.A(net6374),
    .B(net4790),
    .Y(_08165_));
 OAI21x1_ASAP7_75t_R _16207_ (.A1(_00991_),
    .A2(net6327),
    .B(net6336),
    .Y(_08168_));
 INVx1_ASAP7_75t_R _16208_ (.A(_08082_),
    .Y(_08169_));
 OA21x2_ASAP7_75t_R _16210_ (.A1(_08165_),
    .A2(_08168_),
    .B(net5972),
    .Y(_08171_));
 NOR2x1_ASAP7_75t_R _16211_ (.A(net6340),
    .B(_08060_),
    .Y(_08172_));
 INVx1_ASAP7_75t_R _16212_ (.A(_08172_),
    .Y(_08173_));
 INVx1_ASAP7_75t_R _16213_ (.A(_00983_),
    .Y(_08174_));
 NOR2x1_ASAP7_75t_R _16214_ (.A(_08174_),
    .B(net6369),
    .Y(_08175_));
 INVx1_ASAP7_75t_R _16215_ (.A(_08175_),
    .Y(_08176_));
 AO21x1_ASAP7_75t_R _16216_ (.A1(_08173_),
    .A2(net4982),
    .B(net6330),
    .Y(_08177_));
 NAND2x1_ASAP7_75t_R _16217_ (.A(net6369),
    .B(net6340),
    .Y(_08178_));
 AO21x1_ASAP7_75t_R _16218_ (.A1(net5248),
    .A2(_08178_),
    .B(net6375),
    .Y(_08179_));
 NAND3x1_ASAP7_75t_R _16219_ (.A(_08177_),
    .B(net5980),
    .C(_08179_),
    .Y(_08180_));
 AOI21x1_ASAP7_75t_R _16220_ (.A1(_08171_),
    .A2(_08180_),
    .B(net6332),
    .Y(_08181_));
 INVx1_ASAP7_75t_R _16221_ (.A(_08097_),
    .Y(_08182_));
 AOI21x1_ASAP7_75t_R _16222_ (.A1(_08164_),
    .A2(_08181_),
    .B(_08182_),
    .Y(_08183_));
 NAND2x1_ASAP7_75t_R _16223_ (.A(_08148_),
    .B(_08183_),
    .Y(_08184_));
 NAND2x1_ASAP7_75t_R _16224_ (.A(_08174_),
    .B(net6369),
    .Y(_08185_));
 NAND2x1_ASAP7_75t_R _16225_ (.A(net5246),
    .B(_08114_),
    .Y(_08186_));
 AO21x1_ASAP7_75t_R _16227_ (.A1(net4982),
    .A2(net5250),
    .B(net6374),
    .Y(_08188_));
 AOI21x1_ASAP7_75t_R _16228_ (.A1(_08186_),
    .A2(_08188_),
    .B(net6336),
    .Y(_08189_));
 AO21x1_ASAP7_75t_R _16229_ (.A1(net6369),
    .A2(net5261),
    .B(net6327),
    .Y(_08190_));
 AND2x2_ASAP7_75t_R _16230_ (.A(_08190_),
    .B(net6336),
    .Y(_08191_));
 INVx3_ASAP7_75t_R _16231_ (.A(net4792),
    .Y(_08192_));
 NAND2x1_ASAP7_75t_R _16232_ (.A(net6373),
    .B(net6337),
    .Y(_08193_));
 AO21x1_ASAP7_75t_R _16234_ (.A1(_08192_),
    .A2(net5970),
    .B(net6374),
    .Y(_08195_));
 AND2x2_ASAP7_75t_R _16235_ (.A(_08191_),
    .B(_08195_),
    .Y(_08196_));
 OAI21x1_ASAP7_75t_R _16237_ (.A1(_08189_),
    .A2(_08196_),
    .B(net5972),
    .Y(_08198_));
 NAND2x1_ASAP7_75t_R _16238_ (.A(_08104_),
    .B(net6370),
    .Y(_08199_));
 NOR2x1p5_ASAP7_75t_R _16239_ (.A(net6378),
    .B(net4792),
    .Y(_08200_));
 NAND2x1_ASAP7_75t_R _16240_ (.A(_08199_),
    .B(_08200_),
    .Y(_08201_));
 NAND2x1_ASAP7_75t_R _16241_ (.A(_00981_),
    .B(net6338),
    .Y(_08202_));
 AO21x1_ASAP7_75t_R _16243_ (.A1(_08202_),
    .A2(_08139_),
    .B(net6327),
    .Y(_08204_));
 AOI21x1_ASAP7_75t_R _16245_ (.A1(_08201_),
    .A2(_08204_),
    .B(net6335),
    .Y(_08206_));
 NAND2x1_ASAP7_75t_R _16246_ (.A(net6340),
    .B(net6337),
    .Y(_08207_));
 NOR2x1_ASAP7_75t_R _16247_ (.A(net6378),
    .B(_08130_),
    .Y(_08208_));
 NAND2x1_ASAP7_75t_R _16248_ (.A(_08207_),
    .B(_08208_),
    .Y(_08209_));
 AO21x1_ASAP7_75t_R _16249_ (.A1(_08131_),
    .A2(_08207_),
    .B(net6330),
    .Y(_08210_));
 AOI21x1_ASAP7_75t_R _16251_ (.A1(_08209_),
    .A2(_08210_),
    .B(net5980),
    .Y(_08212_));
 OAI21x1_ASAP7_75t_R _16252_ (.A1(_08206_),
    .A2(_08212_),
    .B(net6333),
    .Y(_08213_));
 AOI21x1_ASAP7_75t_R _16253_ (.A1(_08198_),
    .A2(_08213_),
    .B(net6332),
    .Y(_08214_));
 NAND2x1_ASAP7_75t_R _16254_ (.A(net6340),
    .B(net6338),
    .Y(_08215_));
 INVx1_ASAP7_75t_R _16255_ (.A(_00978_),
    .Y(_08216_));
 AO21x1_ASAP7_75t_R _16256_ (.A1(net6372),
    .A2(_08216_),
    .B(net6380),
    .Y(_08217_));
 INVx1_ASAP7_75t_R _16257_ (.A(_08217_),
    .Y(_08218_));
 NAND2x1_ASAP7_75t_R _16258_ (.A(net5968),
    .B(_08218_),
    .Y(_08219_));
 AO21x1_ASAP7_75t_R _16260_ (.A1(net6372),
    .A2(net5322),
    .B(net6327),
    .Y(_08221_));
 OA21x2_ASAP7_75t_R _16261_ (.A1(_08221_),
    .A2(net4792),
    .B(net6334),
    .Y(_08222_));
 AO21x1_ASAP7_75t_R _16262_ (.A1(net6340),
    .A2(net6369),
    .B(net6378),
    .Y(_08223_));
 NAND2x1_ASAP7_75t_R _16263_ (.A(net5977),
    .B(_08223_),
    .Y(_08224_));
 NAND2x1_ASAP7_75t_R _16264_ (.A(net5321),
    .B(net6372),
    .Y(_08225_));
 INVx1_ASAP7_75t_R _16265_ (.A(_08225_),
    .Y(_08226_));
 NOR2x1_ASAP7_75t_R _16266_ (.A(_00979_),
    .B(net6372),
    .Y(_08227_));
 OA21x2_ASAP7_75t_R _16267_ (.A1(_08226_),
    .A2(_08227_),
    .B(net6380),
    .Y(_08228_));
 OAI21x1_ASAP7_75t_R _16268_ (.A1(_08224_),
    .A2(_08228_),
    .B(net6333),
    .Y(_08229_));
 AO21x1_ASAP7_75t_R _16269_ (.A1(_08219_),
    .A2(_08222_),
    .B(_08229_),
    .Y(_08230_));
 NOR2x1_ASAP7_75t_R _16270_ (.A(net5322),
    .B(net6371),
    .Y(_08231_));
 OA21x2_ASAP7_75t_R _16271_ (.A1(net5971),
    .A2(_08231_),
    .B(net6379),
    .Y(_08232_));
 NAND2x1_ASAP7_75t_R _16272_ (.A(net6337),
    .B(_08060_),
    .Y(_08233_));
 AO21x1_ASAP7_75t_R _16273_ (.A1(_08218_),
    .A2(net5967),
    .B(net5979),
    .Y(_08234_));
 AO21x1_ASAP7_75t_R _16274_ (.A1(_08138_),
    .A2(net5969),
    .B(net6377),
    .Y(_08235_));
 AOI21x1_ASAP7_75t_R _16275_ (.A1(_08235_),
    .A2(_08108_),
    .B(net6333),
    .Y(_08236_));
 OAI21x1_ASAP7_75t_R _16276_ (.A1(_08232_),
    .A2(_08234_),
    .B(_08236_),
    .Y(_08237_));
 AOI21x1_ASAP7_75t_R _16278_ (.A1(_08230_),
    .A2(_08237_),
    .B(_08121_),
    .Y(_08239_));
 OAI21x1_ASAP7_75t_R _16279_ (.A1(_08214_),
    .A2(_08239_),
    .B(_08182_),
    .Y(_08240_));
 NAND2x1_ASAP7_75t_R _16280_ (.A(_08184_),
    .B(_08240_),
    .Y(_00000_));
 AO21x1_ASAP7_75t_R _16282_ (.A1(net5968),
    .A2(net5969),
    .B(net6376),
    .Y(_08242_));
 NAND2x1_ASAP7_75t_R _16283_ (.A(net5969),
    .B(_08144_),
    .Y(_08243_));
 AND3x1_ASAP7_75t_R _16284_ (.A(_08242_),
    .B(net5972),
    .C(_08243_),
    .Y(_08244_));
 AO21x1_ASAP7_75t_R _16285_ (.A1(net6338),
    .A2(net6340),
    .B(net6378),
    .Y(_08245_));
 INVx1_ASAP7_75t_R _16286_ (.A(_08185_),
    .Y(_08246_));
 NAND2x1_ASAP7_75t_R _16287_ (.A(net6379),
    .B(_08226_),
    .Y(_08247_));
 OA21x2_ASAP7_75t_R _16288_ (.A1(_08245_),
    .A2(_08246_),
    .B(_08247_),
    .Y(_08248_));
 NAND2x1_ASAP7_75t_R _16289_ (.A(net6378),
    .B(net4984),
    .Y(_08249_));
 AND2x2_ASAP7_75t_R _16290_ (.A(_08249_),
    .B(net6333),
    .Y(_08250_));
 AO21x1_ASAP7_75t_R _16292_ (.A1(_08248_),
    .A2(_08250_),
    .B(net5980),
    .Y(_08252_));
 INVx1_ASAP7_75t_R _16293_ (.A(_00992_),
    .Y(_08253_));
 OR3x1_ASAP7_75t_R _16294_ (.A(net6333),
    .B(_08253_),
    .C(net6329),
    .Y(_08254_));
 INVx1_ASAP7_75t_R _16295_ (.A(_08105_),
    .Y(_08255_));
 AO21x1_ASAP7_75t_R _16296_ (.A1(_08255_),
    .A2(_08132_),
    .B(net6377),
    .Y(_08256_));
 AO21x1_ASAP7_75t_R _16298_ (.A1(_08254_),
    .A2(_08256_),
    .B(net6335),
    .Y(_08258_));
 OAI21x1_ASAP7_75t_R _16299_ (.A1(_08244_),
    .A2(_08252_),
    .B(_08258_),
    .Y(_08259_));
 NOR2x1_ASAP7_75t_R _16300_ (.A(net6332),
    .B(_08259_),
    .Y(_08260_));
 INVx1_ASAP7_75t_R _16301_ (.A(net5572),
    .Y(_08261_));
 NAND2x1_ASAP7_75t_R _16302_ (.A(_08261_),
    .B(net6372),
    .Y(_08262_));
 INVx1_ASAP7_75t_R _16303_ (.A(_08231_),
    .Y(_08263_));
 NAND2x1_ASAP7_75t_R _16304_ (.A(_08262_),
    .B(_08263_),
    .Y(_08264_));
 NOR2x1_ASAP7_75t_R _16306_ (.A(net5261),
    .B(net6372),
    .Y(_08266_));
 AO21x1_ASAP7_75t_R _16307_ (.A1(net6372),
    .A2(_08104_),
    .B(net6327),
    .Y(_08267_));
 NOR2x1_ASAP7_75t_R _16308_ (.A(net5028),
    .B(_08267_),
    .Y(_08268_));
 AOI211x1_ASAP7_75t_R _16309_ (.A1(_08264_),
    .A2(net6326),
    .B(_08268_),
    .C(net5979),
    .Y(_08269_));
 OA21x2_ASAP7_75t_R _16310_ (.A1(net4716),
    .A2(net6378),
    .B(_08117_),
    .Y(_08270_));
 NOR2x1_ASAP7_75t_R _16311_ (.A(net5971),
    .B(net4602),
    .Y(_08271_));
 AO21x1_ASAP7_75t_R _16312_ (.A1(_08270_),
    .A2(_08271_),
    .B(net6333),
    .Y(_08272_));
 OAI21x1_ASAP7_75t_R _16313_ (.A1(_08269_),
    .A2(_08272_),
    .B(net6332),
    .Y(_08273_));
 AO21x1_ASAP7_75t_R _16315_ (.A1(net5968),
    .A2(_08139_),
    .B(net6376),
    .Y(_08275_));
 AO21x1_ASAP7_75t_R _16316_ (.A1(_08275_),
    .A2(_08243_),
    .B(net6335),
    .Y(_08276_));
 AO21x1_ASAP7_75t_R _16317_ (.A1(_08173_),
    .A2(_08138_),
    .B(net6377),
    .Y(_08277_));
 AO21x1_ASAP7_75t_R _16318_ (.A1(net4982),
    .A2(net4791),
    .B(net6326),
    .Y(_08278_));
 AO21x1_ASAP7_75t_R _16319_ (.A1(_08277_),
    .A2(_08278_),
    .B(net5978),
    .Y(_08279_));
 AOI21x1_ASAP7_75t_R _16321_ (.A1(_08276_),
    .A2(_08279_),
    .B(net5972),
    .Y(_08281_));
 OAI21x1_ASAP7_75t_R _16322_ (.A1(_08273_),
    .A2(_08281_),
    .B(_08182_),
    .Y(_08282_));
 AO21x1_ASAP7_75t_R _16323_ (.A1(net6339),
    .A2(net5252),
    .B(net6334),
    .Y(_08283_));
 OA21x2_ASAP7_75t_R _16324_ (.A1(_08268_),
    .A2(_08283_),
    .B(net6333),
    .Y(_08284_));
 INVx1_ASAP7_75t_R _16325_ (.A(_08233_),
    .Y(_08285_));
 OA21x2_ASAP7_75t_R _16326_ (.A1(_08221_),
    .A2(_08285_),
    .B(net6334),
    .Y(_08286_));
 OAI21x1_ASAP7_75t_R _16327_ (.A1(net6379),
    .A2(net4715),
    .B(_08286_),
    .Y(_08287_));
 AOI21x1_ASAP7_75t_R _16328_ (.A1(_08284_),
    .A2(_08287_),
    .B(_08121_),
    .Y(_08288_));
 NAND2x1_ASAP7_75t_R _16329_ (.A(_08143_),
    .B(net6372),
    .Y(_08289_));
 AO21x1_ASAP7_75t_R _16331_ (.A1(_08192_),
    .A2(_08289_),
    .B(net6326),
    .Y(_08291_));
 AO21x1_ASAP7_75t_R _16332_ (.A1(_08173_),
    .A2(net4982),
    .B(net6379),
    .Y(_08292_));
 AOI21x1_ASAP7_75t_R _16333_ (.A1(_08291_),
    .A2(_08292_),
    .B(net5979),
    .Y(_08293_));
 NAND2x1_ASAP7_75t_R _16334_ (.A(net5981),
    .B(_00972_),
    .Y(_08294_));
 AO21x1_ASAP7_75t_R _16335_ (.A1(_08294_),
    .A2(net5968),
    .B(net6328),
    .Y(_08295_));
 NOR2x1_ASAP7_75t_R _16336_ (.A(net6339),
    .B(net5029),
    .Y(_08296_));
 INVx1_ASAP7_75t_R _16337_ (.A(_08296_),
    .Y(_08297_));
 AO21x1_ASAP7_75t_R _16338_ (.A1(_08297_),
    .A2(_08131_),
    .B(net6375),
    .Y(_08298_));
 AOI21x1_ASAP7_75t_R _16339_ (.A1(_08295_),
    .A2(_08298_),
    .B(net6334),
    .Y(_08299_));
 OAI21x1_ASAP7_75t_R _16340_ (.A1(_08293_),
    .A2(_08299_),
    .B(net5972),
    .Y(_08300_));
 AOI21x1_ASAP7_75t_R _16341_ (.A1(_08288_),
    .A2(_08300_),
    .B(_08182_),
    .Y(_08301_));
 NAND2x1_ASAP7_75t_R _16342_ (.A(_00986_),
    .B(net6380),
    .Y(_08302_));
 AND2x2_ASAP7_75t_R _16343_ (.A(net6334),
    .B(_08302_),
    .Y(_08303_));
 AO21x1_ASAP7_75t_R _16344_ (.A1(net5967),
    .A2(_08289_),
    .B(net6379),
    .Y(_08304_));
 AOI21x1_ASAP7_75t_R _16345_ (.A1(_08303_),
    .A2(_08304_),
    .B(net6333),
    .Y(_08305_));
 AO21x1_ASAP7_75t_R _16346_ (.A1(_08263_),
    .A2(net4791),
    .B(net6326),
    .Y(_08306_));
 AO21x1_ASAP7_75t_R _16347_ (.A1(net5248),
    .A2(_08289_),
    .B(net6379),
    .Y(_08307_));
 NAND3x1_ASAP7_75t_R _16348_ (.A(_08306_),
    .B(_08307_),
    .C(net5978),
    .Y(_08308_));
 AOI21x1_ASAP7_75t_R _16349_ (.A1(_08305_),
    .A2(_08308_),
    .B(net6332),
    .Y(_08309_));
 NAND2x1_ASAP7_75t_R _16350_ (.A(_08207_),
    .B(_08128_),
    .Y(_08310_));
 AOI21x1_ASAP7_75t_R _16351_ (.A1(_08247_),
    .A2(_08310_),
    .B(net6335),
    .Y(_08311_));
 AND2x2_ASAP7_75t_R _16352_ (.A(_08178_),
    .B(_08114_),
    .Y(_08312_));
 OA21x2_ASAP7_75t_R _16353_ (.A1(net6371),
    .A2(net5249),
    .B(net6330),
    .Y(_08313_));
 AND2x2_ASAP7_75t_R _16354_ (.A(_08313_),
    .B(_08173_),
    .Y(_08314_));
 OA21x2_ASAP7_75t_R _16355_ (.A1(_08312_),
    .A2(_08314_),
    .B(net6335),
    .Y(_08315_));
 OAI21x1_ASAP7_75t_R _16356_ (.A1(_08311_),
    .A2(_08315_),
    .B(net6333),
    .Y(_08316_));
 NAND2x1_ASAP7_75t_R _16357_ (.A(_08316_),
    .B(_08309_),
    .Y(_08317_));
 NAND2x1_ASAP7_75t_R _16358_ (.A(_08301_),
    .B(_08317_),
    .Y(_08318_));
 OAI21x1_ASAP7_75t_R _16359_ (.A1(_08260_),
    .A2(_08282_),
    .B(_08318_),
    .Y(_00001_));
 NAND2x1_ASAP7_75t_R _16360_ (.A(net6378),
    .B(net5981),
    .Y(_08319_));
 INVx1_ASAP7_75t_R _16361_ (.A(net5970),
    .Y(_08320_));
 AO21x1_ASAP7_75t_R _16362_ (.A1(_08319_),
    .A2(net6331),
    .B(_08320_),
    .Y(_08321_));
 AND3x1_ASAP7_75t_R _16363_ (.A(_08321_),
    .B(net6335),
    .C(_08129_),
    .Y(_08322_));
 OA22x2_ASAP7_75t_R _16364_ (.A1(_00991_),
    .A2(net6374),
    .B1(_08190_),
    .B2(net5247),
    .Y(_08323_));
 AO21x1_ASAP7_75t_R _16365_ (.A1(_08323_),
    .A2(_08117_),
    .B(net5972),
    .Y(_08324_));
 NOR2x1_ASAP7_75t_R _16366_ (.A(_08322_),
    .B(_08324_),
    .Y(_08325_));
 AND3x1_ASAP7_75t_R _16367_ (.A(_08202_),
    .B(net6374),
    .C(net4790),
    .Y(_08326_));
 AND2x2_ASAP7_75t_R _16368_ (.A(_08128_),
    .B(_08139_),
    .Y(_08327_));
 OAI21x1_ASAP7_75t_R _16369_ (.A1(_08326_),
    .A2(_08327_),
    .B(net6335),
    .Y(_08328_));
 NAND2x1_ASAP7_75t_R _16370_ (.A(_00992_),
    .B(net6329),
    .Y(_08329_));
 NOR2x1_ASAP7_75t_R _16371_ (.A(net6329),
    .B(_08127_),
    .Y(_08330_));
 AOI21x1_ASAP7_75t_R _16372_ (.A1(_08207_),
    .A2(_08330_),
    .B(net6335),
    .Y(_08331_));
 AOI21x1_ASAP7_75t_R _16373_ (.A1(_08329_),
    .A2(_08331_),
    .B(net6333),
    .Y(_08332_));
 AO21x1_ASAP7_75t_R _16374_ (.A1(_08328_),
    .A2(_08332_),
    .B(net5975),
    .Y(_08333_));
 AO21x1_ASAP7_75t_R _16375_ (.A1(_08233_),
    .A2(net5245),
    .B(net6326),
    .Y(_08334_));
 OA21x2_ASAP7_75t_R _16376_ (.A1(net6380),
    .A2(_00988_),
    .B(net6334),
    .Y(_08335_));
 NOR2x1_ASAP7_75t_R _16377_ (.A(net6334),
    .B(_08218_),
    .Y(_08336_));
 NAND2x1_ASAP7_75t_R _16378_ (.A(_00990_),
    .B(net6380),
    .Y(_08337_));
 AOI22x1_ASAP7_75t_R _16379_ (.A1(_08334_),
    .A2(_08335_),
    .B1(_08336_),
    .B2(_08337_),
    .Y(_08338_));
 NAND2x1_ASAP7_75t_R _16380_ (.A(net5972),
    .B(_08338_),
    .Y(_08339_));
 INVx1_ASAP7_75t_R _16381_ (.A(_08266_),
    .Y(_08340_));
 AO21x1_ASAP7_75t_R _16382_ (.A1(_08340_),
    .A2(_08289_),
    .B(net6326),
    .Y(_08341_));
 OA21x2_ASAP7_75t_R _16383_ (.A1(net4982),
    .A2(net6379),
    .B(net5980),
    .Y(_08342_));
 AOI21x1_ASAP7_75t_R _16384_ (.A1(_08341_),
    .A2(_08342_),
    .B(net5972),
    .Y(_08343_));
 NAND2x1_ASAP7_75t_R _16385_ (.A(net5323),
    .B(net6371),
    .Y(_08344_));
 AO21x1_ASAP7_75t_R _16386_ (.A1(net5968),
    .A2(_08344_),
    .B(net6326),
    .Y(_08345_));
 NAND3x1_ASAP7_75t_R _16387_ (.A(_08256_),
    .B(_08345_),
    .C(net6334),
    .Y(_08346_));
 AOI21x1_ASAP7_75t_R _16388_ (.A1(_08343_),
    .A2(_08346_),
    .B(net6332),
    .Y(_08347_));
 AOI21x1_ASAP7_75t_R _16389_ (.A1(_08339_),
    .A2(_08347_),
    .B(_08182_),
    .Y(_08348_));
 OAI21x1_ASAP7_75t_R _16390_ (.A1(_08325_),
    .A2(_08333_),
    .B(_08348_),
    .Y(_08349_));
 INVx1_ASAP7_75t_R _16391_ (.A(_00982_),
    .Y(_08350_));
 AO21x1_ASAP7_75t_R _16392_ (.A1(net6338),
    .A2(_08350_),
    .B(net6327),
    .Y(_08351_));
 INVx1_ASAP7_75t_R _16393_ (.A(net5322),
    .Y(_08352_));
 NAND2x1_ASAP7_75t_R _16394_ (.A(_08352_),
    .B(net6370),
    .Y(_08353_));
 AOI21x1_ASAP7_75t_R _16395_ (.A1(net4979),
    .A2(_08208_),
    .B(net5980),
    .Y(_08354_));
 OA21x2_ASAP7_75t_R _16396_ (.A1(_08320_),
    .A2(_08351_),
    .B(_08354_),
    .Y(_08355_));
 NAND2x1p5_ASAP7_75t_R _16397_ (.A(net4603),
    .B(net4790),
    .Y(_08356_));
 NAND2x1_ASAP7_75t_R _16398_ (.A(_08350_),
    .B(net6369),
    .Y(_08357_));
 AO21x1_ASAP7_75t_R _16399_ (.A1(_08131_),
    .A2(_08357_),
    .B(net6375),
    .Y(_08358_));
 AOI21x1_ASAP7_75t_R _16400_ (.A1(_08358_),
    .A2(_08356_),
    .B(net6335),
    .Y(_08359_));
 OA21x2_ASAP7_75t_R _16401_ (.A1(_08359_),
    .A2(_08355_),
    .B(net6333),
    .Y(_08360_));
 AO21x1_ASAP7_75t_R _16403_ (.A1(_08131_),
    .A2(net4980),
    .B(net6328),
    .Y(_08362_));
 NOR2x1_ASAP7_75t_R _16404_ (.A(net6378),
    .B(_08353_),
    .Y(_08363_));
 NOR2x1_ASAP7_75t_R _16405_ (.A(_08117_),
    .B(_08363_),
    .Y(_08364_));
 NAND3x1_ASAP7_75t_R _16406_ (.A(_08362_),
    .B(net4983),
    .C(_08364_),
    .Y(_08365_));
 INVx1_ASAP7_75t_R _16407_ (.A(_08127_),
    .Y(_08366_));
 AO21x1_ASAP7_75t_R _16408_ (.A1(_08366_),
    .A2(net4980),
    .B(net6328),
    .Y(_08367_));
 AOI211x1_ASAP7_75t_R _16409_ (.A1(net6327),
    .A2(net5251),
    .B(net4985),
    .C(net6334),
    .Y(_08368_));
 AOI21x1_ASAP7_75t_R _16410_ (.A1(_08367_),
    .A2(_08368_),
    .B(net6333),
    .Y(_08369_));
 AO21x1_ASAP7_75t_R _16411_ (.A1(_08365_),
    .A2(_08369_),
    .B(net5975),
    .Y(_08370_));
 NAND2x1_ASAP7_75t_R _16412_ (.A(net5322),
    .B(net6371),
    .Y(_08371_));
 NAND2x1_ASAP7_75t_R _16413_ (.A(_08371_),
    .B(_08313_),
    .Y(_08372_));
 AOI21x1_ASAP7_75t_R _16414_ (.A1(_08372_),
    .A2(_08334_),
    .B(net5979),
    .Y(_08373_));
 AO21x1_ASAP7_75t_R _16415_ (.A1(net5248),
    .A2(_08289_),
    .B(net6326),
    .Y(_08374_));
 AO21x1_ASAP7_75t_R _16416_ (.A1(_08366_),
    .A2(net4791),
    .B(net6379),
    .Y(_08375_));
 AOI21x1_ASAP7_75t_R _16417_ (.A1(_08374_),
    .A2(_08375_),
    .B(net6334),
    .Y(_08376_));
 OAI21x1_ASAP7_75t_R _16418_ (.A1(_08373_),
    .A2(_08376_),
    .B(net5972),
    .Y(_08377_));
 AO21x1_ASAP7_75t_R _16419_ (.A1(_08263_),
    .A2(_08344_),
    .B(net6326),
    .Y(_08378_));
 AOI21x1_ASAP7_75t_R _16420_ (.A1(_08378_),
    .A2(_08336_),
    .B(net5972),
    .Y(_08379_));
 NOR2x1_ASAP7_75t_R _16421_ (.A(net6330),
    .B(_08130_),
    .Y(_08380_));
 NAND2x1_ASAP7_75t_R _16422_ (.A(_08262_),
    .B(_08380_),
    .Y(_08381_));
 AOI21x1_ASAP7_75t_R _16423_ (.A1(net6372),
    .A2(net6337),
    .B(net6378),
    .Y(_08382_));
 NAND2x1_ASAP7_75t_R _16424_ (.A(_08340_),
    .B(_08382_),
    .Y(_08383_));
 AO21x1_ASAP7_75t_R _16425_ (.A1(_08381_),
    .A2(_08383_),
    .B(net5976),
    .Y(_08384_));
 AOI21x1_ASAP7_75t_R _16426_ (.A1(_08379_),
    .A2(_08384_),
    .B(net6332),
    .Y(_08385_));
 AOI21x1_ASAP7_75t_R _16427_ (.A1(_08377_),
    .A2(_08385_),
    .B(_08097_),
    .Y(_08386_));
 OAI21x1_ASAP7_75t_R _16428_ (.A1(_08370_),
    .A2(_08360_),
    .B(_08386_),
    .Y(_08387_));
 NAND2x1_ASAP7_75t_R _16429_ (.A(_08349_),
    .B(_08387_),
    .Y(_00002_));
 AO21x1_ASAP7_75t_R _16430_ (.A1(_08173_),
    .A2(_08340_),
    .B(net6379),
    .Y(_08388_));
 OAI21x1_ASAP7_75t_R _16431_ (.A1(net5973),
    .A2(_08221_),
    .B(_08388_),
    .Y(_08389_));
 INVx1_ASAP7_75t_R _16432_ (.A(_08115_),
    .Y(_08390_));
 OA21x2_ASAP7_75t_R _16433_ (.A1(_08390_),
    .A2(net6330),
    .B(net6333),
    .Y(_08391_));
 NAND2x1_ASAP7_75t_R _16434_ (.A(_08391_),
    .B(_08358_),
    .Y(_08392_));
 OAI21x1_ASAP7_75t_R _16435_ (.A1(net6333),
    .A2(_08389_),
    .B(_08392_),
    .Y(_08393_));
 NOR2x1p5_ASAP7_75t_R _16436_ (.A(net6374),
    .B(_08192_),
    .Y(_08394_));
 AO21x1_ASAP7_75t_R _16437_ (.A1(net5561),
    .A2(net6376),
    .B(net5980),
    .Y(_08395_));
 AO21x1_ASAP7_75t_R _16438_ (.A1(_08394_),
    .A2(net6333),
    .B(_08395_),
    .Y(_08396_));
 INVx1_ASAP7_75t_R _16439_ (.A(_00981_),
    .Y(_08397_));
 AO21x1_ASAP7_75t_R _16440_ (.A1(net6369),
    .A2(_08397_),
    .B(net6378),
    .Y(_08398_));
 NOR2x1_ASAP7_75t_R _16441_ (.A(net5974),
    .B(_08398_),
    .Y(_08399_));
 NOR2x1_ASAP7_75t_R _16442_ (.A(net5029),
    .B(net6331),
    .Y(_08400_));
 OA21x2_ASAP7_75t_R _16443_ (.A1(_08399_),
    .A2(_08400_),
    .B(net5972),
    .Y(_08401_));
 OAI21x1_ASAP7_75t_R _16444_ (.A1(_08396_),
    .A2(_08401_),
    .B(net5975),
    .Y(_08402_));
 AOI21x1_ASAP7_75t_R _16445_ (.A1(net5980),
    .A2(_08393_),
    .B(_08402_),
    .Y(_08403_));
 AO21x1_ASAP7_75t_R _16446_ (.A1(net5968),
    .A2(_08357_),
    .B(net6326),
    .Y(_08404_));
 AOI21x1_ASAP7_75t_R _16447_ (.A1(_08404_),
    .A2(_08256_),
    .B(net6335),
    .Y(_08405_));
 OAI21x1_ASAP7_75t_R _16448_ (.A1(_08354_),
    .A2(_08405_),
    .B(net5972),
    .Y(_08406_));
 NAND2x1_ASAP7_75t_R _16449_ (.A(_08371_),
    .B(_08200_),
    .Y(_08407_));
 AO21x1_ASAP7_75t_R _16450_ (.A1(_08390_),
    .A2(_08178_),
    .B(net6330),
    .Y(_08408_));
 AOI21x1_ASAP7_75t_R _16451_ (.A1(_08407_),
    .A2(_08408_),
    .B(net5980),
    .Y(_08409_));
 AOI21x1_ASAP7_75t_R _16452_ (.A1(_08310_),
    .A2(_08177_),
    .B(net6335),
    .Y(_08410_));
 OAI21x1_ASAP7_75t_R _16453_ (.A1(_08409_),
    .A2(_08410_),
    .B(net6333),
    .Y(_08411_));
 AOI21x1_ASAP7_75t_R _16454_ (.A1(_08406_),
    .A2(_08411_),
    .B(net5975),
    .Y(_08412_));
 OAI21x1_ASAP7_75t_R _16455_ (.A1(_08403_),
    .A2(_08412_),
    .B(_08182_),
    .Y(_08413_));
 AO21x1_ASAP7_75t_R _16456_ (.A1(net5971),
    .A2(net6330),
    .B(_08117_),
    .Y(_08414_));
 AO21x1_ASAP7_75t_R _16457_ (.A1(_08297_),
    .A2(net4982),
    .B(net6327),
    .Y(_08415_));
 OAI21x1_ASAP7_75t_R _16458_ (.A1(net6378),
    .A2(_08202_),
    .B(_08415_),
    .Y(_08416_));
 AOI21x1_ASAP7_75t_R _16459_ (.A1(net4789),
    .A2(_08382_),
    .B(net6334),
    .Y(_08417_));
 AO21x1_ASAP7_75t_R _16460_ (.A1(_08263_),
    .A2(_08289_),
    .B(net6330),
    .Y(_08418_));
 AOI21x1_ASAP7_75t_R _16461_ (.A1(_08417_),
    .A2(_08418_),
    .B(net5972),
    .Y(_08419_));
 OAI21x1_ASAP7_75t_R _16462_ (.A1(net5559),
    .A2(_08416_),
    .B(_08419_),
    .Y(_08420_));
 INVx1_ASAP7_75t_R _16463_ (.A(net4602),
    .Y(_08421_));
 AO21x1_ASAP7_75t_R _16464_ (.A1(_08173_),
    .A2(_08207_),
    .B(net6375),
    .Y(_08422_));
 OAI21x1_ASAP7_75t_R _16465_ (.A1(_08421_),
    .A2(net5560),
    .B(_08422_),
    .Y(_08423_));
 NAND2x1_ASAP7_75t_R _16466_ (.A(net5968),
    .B(_08382_),
    .Y(_08424_));
 AOI21x1_ASAP7_75t_R _16467_ (.A1(_08424_),
    .A2(_08191_),
    .B(net6333),
    .Y(_08425_));
 OAI21x1_ASAP7_75t_R _16468_ (.A1(net6334),
    .A2(_08423_),
    .B(_08425_),
    .Y(_08426_));
 AOI21x1_ASAP7_75t_R _16469_ (.A1(_08420_),
    .A2(_08426_),
    .B(net6332),
    .Y(_08427_));
 AO21x1_ASAP7_75t_R _16470_ (.A1(_08202_),
    .A2(net5245),
    .B(net6327),
    .Y(_08428_));
 AO21x1_ASAP7_75t_R _16471_ (.A1(net4716),
    .A2(net4791),
    .B(net6378),
    .Y(_08429_));
 AOI21x1_ASAP7_75t_R _16472_ (.A1(_08428_),
    .A2(_08429_),
    .B(net6334),
    .Y(_08430_));
 AO21x1_ASAP7_75t_R _16473_ (.A1(_08192_),
    .A2(net5250),
    .B(net6378),
    .Y(_08431_));
 NAND2x1_ASAP7_75t_R _16474_ (.A(net6340),
    .B(net5982),
    .Y(_08432_));
 INVx1_ASAP7_75t_R _16475_ (.A(_08432_),
    .Y(_08433_));
 OAI21x1_ASAP7_75t_R _16476_ (.A1(net5971),
    .A2(_08433_),
    .B(net6378),
    .Y(_08434_));
 AOI21x1_ASAP7_75t_R _16477_ (.A1(_08431_),
    .A2(_08434_),
    .B(net5977),
    .Y(_08435_));
 OAI21x1_ASAP7_75t_R _16478_ (.A1(_08430_),
    .A2(_08435_),
    .B(net6333),
    .Y(_08436_));
 AO21x1_ASAP7_75t_R _16479_ (.A1(_08192_),
    .A2(_08357_),
    .B(net6379),
    .Y(_08437_));
 AO21x1_ASAP7_75t_R _16480_ (.A1(_08366_),
    .A2(_08353_),
    .B(net6330),
    .Y(_08438_));
 AOI21x1_ASAP7_75t_R _16481_ (.A1(_08437_),
    .A2(_08438_),
    .B(net5976),
    .Y(_08439_));
 AO21x1_ASAP7_75t_R _16482_ (.A1(net6372),
    .A2(_08216_),
    .B(net6326),
    .Y(_08440_));
 AOI21x1_ASAP7_75t_R _16483_ (.A1(_08440_),
    .A2(_08422_),
    .B(net6334),
    .Y(_08441_));
 OAI21x1_ASAP7_75t_R _16484_ (.A1(_08439_),
    .A2(_08441_),
    .B(net5972),
    .Y(_08442_));
 AOI21x1_ASAP7_75t_R _16485_ (.A1(_08436_),
    .A2(_08442_),
    .B(net5975),
    .Y(_08443_));
 OAI21x1_ASAP7_75t_R _16486_ (.A1(_08427_),
    .A2(_08443_),
    .B(_08097_),
    .Y(_08444_));
 NAND2x1_ASAP7_75t_R _16487_ (.A(_08413_),
    .B(_08444_),
    .Y(_00003_));
 NAND2x1_ASAP7_75t_R _16488_ (.A(net4790),
    .B(_08313_),
    .Y(_08445_));
 AO21x1_ASAP7_75t_R _16489_ (.A1(net6372),
    .A2(net5572),
    .B(net6380),
    .Y(_08446_));
 AND3x1_ASAP7_75t_R _16490_ (.A(_08267_),
    .B(_08446_),
    .C(net6334),
    .Y(_08447_));
 AOI211x1_ASAP7_75t_R _16491_ (.A1(net4532),
    .A2(_08445_),
    .B(_08447_),
    .C(net5972),
    .Y(_08448_));
 AO21x1_ASAP7_75t_R _16492_ (.A1(_08320_),
    .A2(net6326),
    .B(net5978),
    .Y(_08449_));
 OAI21x1_ASAP7_75t_R _16493_ (.A1(net6377),
    .A2(net4982),
    .B(_08243_),
    .Y(_08450_));
 NAND2x1_ASAP7_75t_R _16494_ (.A(net6331),
    .B(net5980),
    .Y(_08451_));
 AO21x1_ASAP7_75t_R _16495_ (.A1(_08208_),
    .A2(_08371_),
    .B(_08451_),
    .Y(_08452_));
 OAI21x1_ASAP7_75t_R _16496_ (.A1(_08449_),
    .A2(_08450_),
    .B(_08452_),
    .Y(_08453_));
 OAI21x1_ASAP7_75t_R _16497_ (.A1(net6333),
    .A2(_08453_),
    .B(_08182_),
    .Y(_08454_));
 OAI21x1_ASAP7_75t_R _16498_ (.A1(_08448_),
    .A2(_08454_),
    .B(net6332),
    .Y(_08455_));
 NOR2x1_ASAP7_75t_R _16499_ (.A(net5561),
    .B(net5980),
    .Y(_08456_));
 AO21x1_ASAP7_75t_R _16500_ (.A1(_08456_),
    .A2(_08158_),
    .B(net5972),
    .Y(_08457_));
 OAI21x1_ASAP7_75t_R _16501_ (.A1(_08246_),
    .A2(_08245_),
    .B(net5980),
    .Y(_08458_));
 NAND2x1_ASAP7_75t_R _16502_ (.A(net6373),
    .B(net5983),
    .Y(_08459_));
 AND3x1_ASAP7_75t_R _16503_ (.A(_08459_),
    .B(net6376),
    .C(net5968),
    .Y(_08460_));
 NOR2x1_ASAP7_75t_R _16504_ (.A(_08458_),
    .B(_08460_),
    .Y(_08461_));
 OAI21x1_ASAP7_75t_R _16505_ (.A1(_08457_),
    .A2(_08461_),
    .B(_08097_),
    .Y(_08462_));
 NAND2x1_ASAP7_75t_R _16506_ (.A(net5246),
    .B(_08233_),
    .Y(_08463_));
 AND3x1_ASAP7_75t_R _16507_ (.A(_08432_),
    .B(net6330),
    .C(net5970),
    .Y(_08464_));
 AO21x1_ASAP7_75t_R _16508_ (.A1(net6376),
    .A2(_08463_),
    .B(_08464_),
    .Y(_08465_));
 AO21x1_ASAP7_75t_R _16509_ (.A1(_08331_),
    .A2(_08242_),
    .B(net6333),
    .Y(_08466_));
 AOI21x1_ASAP7_75t_R _16510_ (.A1(net6335),
    .A2(_08465_),
    .B(_08466_),
    .Y(_08467_));
 NOR2x1_ASAP7_75t_R _16511_ (.A(_08462_),
    .B(_08467_),
    .Y(_08468_));
 OAI22x1_ASAP7_75t_R _16512_ (.A1(net6331),
    .A2(net5261),
    .B1(net5323),
    .B2(net6378),
    .Y(_08469_));
 AO21x1_ASAP7_75t_R _16513_ (.A1(_08469_),
    .A2(net5978),
    .B(net5972),
    .Y(_08470_));
 AO21x1_ASAP7_75t_R _16514_ (.A1(_08366_),
    .A2(_08357_),
    .B(net6326),
    .Y(_08471_));
 OA21x2_ASAP7_75t_R _16515_ (.A1(net5248),
    .A2(net6377),
    .B(net6335),
    .Y(_08472_));
 AND2x2_ASAP7_75t_R _16516_ (.A(_08471_),
    .B(_08472_),
    .Y(_08473_));
 OAI21x1_ASAP7_75t_R _16517_ (.A1(_08470_),
    .A2(_08473_),
    .B(_08182_),
    .Y(_08474_));
 INVx1_ASAP7_75t_R _16518_ (.A(_08404_),
    .Y(_08475_));
 OAI21x1_ASAP7_75t_R _16519_ (.A1(_08475_),
    .A2(_08464_),
    .B(net6335),
    .Y(_08476_));
 AO21x1_ASAP7_75t_R _16520_ (.A1(_08210_),
    .A2(_08140_),
    .B(net6335),
    .Y(_08477_));
 AOI21x1_ASAP7_75t_R _16521_ (.A1(_08476_),
    .A2(_08477_),
    .B(net6333),
    .Y(_08478_));
 OAI21x1_ASAP7_75t_R _16522_ (.A1(_08474_),
    .A2(_08478_),
    .B(net5975),
    .Y(_08479_));
 OA21x2_ASAP7_75t_R _16523_ (.A1(net6370),
    .A2(_08352_),
    .B(net6328),
    .Y(_08480_));
 AOI211x1_ASAP7_75t_R _16524_ (.A1(net4601),
    .A2(_08480_),
    .B(_08159_),
    .C(net6334),
    .Y(_08481_));
 AOI21x1_ASAP7_75t_R _16525_ (.A1(net4790),
    .A2(_08390_),
    .B(net6330),
    .Y(_08482_));
 OAI21x1_ASAP7_75t_R _16526_ (.A1(net4531),
    .A2(_08482_),
    .B(net6333),
    .Y(_08483_));
 OAI21x1_ASAP7_75t_R _16527_ (.A1(_08483_),
    .A2(_08481_),
    .B(_08097_),
    .Y(_08484_));
 NOR2x1_ASAP7_75t_R _16528_ (.A(net6326),
    .B(_08157_),
    .Y(_08485_));
 NAND2x1_ASAP7_75t_R _16529_ (.A(net5969),
    .B(_08485_),
    .Y(_08486_));
 AO21x1_ASAP7_75t_R _16530_ (.A1(_08486_),
    .A2(_08372_),
    .B(net5978),
    .Y(_08487_));
 AO21x1_ASAP7_75t_R _16531_ (.A1(_08459_),
    .A2(net4982),
    .B(net6326),
    .Y(_08488_));
 AO21x1_ASAP7_75t_R _16532_ (.A1(_08488_),
    .A2(_08307_),
    .B(net6335),
    .Y(_08489_));
 AOI21x1_ASAP7_75t_R _16533_ (.A1(_08487_),
    .A2(_08489_),
    .B(net6333),
    .Y(_08490_));
 NOR2x1_ASAP7_75t_R _16534_ (.A(_08490_),
    .B(_08484_),
    .Y(_08491_));
 OAI22x1_ASAP7_75t_R _16535_ (.A1(_08455_),
    .A2(_08468_),
    .B1(_08491_),
    .B2(_08479_),
    .Y(_00004_));
 OA21x2_ASAP7_75t_R _16536_ (.A1(net6331),
    .A2(net5242),
    .B(net6334),
    .Y(_08492_));
 AO21x1_ASAP7_75t_R _16537_ (.A1(net4715),
    .A2(_08353_),
    .B(net6378),
    .Y(_08493_));
 NAND2x1_ASAP7_75t_R _16538_ (.A(_08492_),
    .B(_08493_),
    .Y(_08494_));
 AO21x1_ASAP7_75t_R _16539_ (.A1(_08131_),
    .A2(net4980),
    .B(net6375),
    .Y(_08495_));
 AOI21x1_ASAP7_75t_R _16540_ (.A1(_08495_),
    .A2(net4532),
    .B(net5975),
    .Y(_08496_));
 AO21x1_ASAP7_75t_R _16541_ (.A1(net4789),
    .A2(net5250),
    .B(net6328),
    .Y(_08497_));
 OA21x2_ASAP7_75t_R _16542_ (.A1(net6375),
    .A2(_08192_),
    .B(_08364_),
    .Y(_08498_));
 NOR2x1_ASAP7_75t_R _16543_ (.A(net5323),
    .B(net6378),
    .Y(_08499_));
 AO22x1_ASAP7_75t_R _16544_ (.A1(net5242),
    .A2(net6378),
    .B1(_08499_),
    .B2(net6339),
    .Y(_08500_));
 AO21x1_ASAP7_75t_R _16545_ (.A1(_08500_),
    .A2(_08117_),
    .B(net6332),
    .Y(_08501_));
 AOI21x1_ASAP7_75t_R _16546_ (.A1(_08497_),
    .A2(_08498_),
    .B(_08501_),
    .Y(_08502_));
 AOI211x1_ASAP7_75t_R _16547_ (.A1(_08494_),
    .A2(_08496_),
    .B(_08502_),
    .C(net6333),
    .Y(_08503_));
 NOR2x1_ASAP7_75t_R _16548_ (.A(net4981),
    .B(_08380_),
    .Y(_08504_));
 AND2x2_ASAP7_75t_R _16549_ (.A(_08504_),
    .B(_08270_),
    .Y(_08505_));
 AO21x1_ASAP7_75t_R _16550_ (.A1(_08118_),
    .A2(_08221_),
    .B(net6332),
    .Y(_08506_));
 OA21x2_ASAP7_75t_R _16551_ (.A1(_08505_),
    .A2(_08506_),
    .B(net6333),
    .Y(_08507_));
 AOI21x1_ASAP7_75t_R _16552_ (.A1(_08319_),
    .A2(_08209_),
    .B(net6335),
    .Y(_08508_));
 AO21x1_ASAP7_75t_R _16553_ (.A1(_08340_),
    .A2(net5244),
    .B(net6326),
    .Y(_08509_));
 AO21x1_ASAP7_75t_R _16554_ (.A1(_08366_),
    .A2(_08357_),
    .B(net6379),
    .Y(_08510_));
 AOI21x1_ASAP7_75t_R _16555_ (.A1(_08509_),
    .A2(_08510_),
    .B(net5979),
    .Y(_08511_));
 OAI21x1_ASAP7_75t_R _16556_ (.A1(_08508_),
    .A2(_08511_),
    .B(net6332),
    .Y(_08512_));
 AO21x1_ASAP7_75t_R _16557_ (.A1(_08507_),
    .A2(_08512_),
    .B(_08097_),
    .Y(_08513_));
 NAND2x1_ASAP7_75t_R _16558_ (.A(_08371_),
    .B(_08144_),
    .Y(_08514_));
 AOI21x1_ASAP7_75t_R _16559_ (.A1(_08514_),
    .A2(_08235_),
    .B(net6334),
    .Y(_08515_));
 AO21x1_ASAP7_75t_R _16560_ (.A1(net5248),
    .A2(_08357_),
    .B(net6379),
    .Y(_08516_));
 AO21x1_ASAP7_75t_R _16561_ (.A1(net5968),
    .A2(_08289_),
    .B(net6326),
    .Y(_08517_));
 AOI21x1_ASAP7_75t_R _16562_ (.A1(_08516_),
    .A2(_08517_),
    .B(net5978),
    .Y(_08518_));
 OAI21x1_ASAP7_75t_R _16563_ (.A1(_08515_),
    .A2(_08518_),
    .B(net6332),
    .Y(_08519_));
 NAND2x1_ASAP7_75t_R _16564_ (.A(net6333),
    .B(_08519_),
    .Y(_08520_));
 AO21x1_ASAP7_75t_R _16565_ (.A1(_08294_),
    .A2(_08178_),
    .B(net6375),
    .Y(_08521_));
 NAND3x1_ASAP7_75t_R _16566_ (.A(_08521_),
    .B(net4717),
    .C(_08492_),
    .Y(_08522_));
 NOR2x1_ASAP7_75t_R _16567_ (.A(net6329),
    .B(net5983),
    .Y(_08523_));
 OAI21x1_ASAP7_75t_R _16568_ (.A1(_08523_),
    .A2(_08464_),
    .B(net5980),
    .Y(_08524_));
 AND3x1_ASAP7_75t_R _16569_ (.A(_08522_),
    .B(net5975),
    .C(_08524_),
    .Y(_08525_));
 NAND2x1_ASAP7_75t_R _16570_ (.A(net6334),
    .B(net5244),
    .Y(_08526_));
 OA21x2_ASAP7_75t_R _16571_ (.A1(_08526_),
    .A2(_08313_),
    .B(net6332),
    .Y(_08527_));
 NOR2x1_ASAP7_75t_R _16572_ (.A(net6334),
    .B(_08200_),
    .Y(_08528_));
 NAND2x1_ASAP7_75t_R _16573_ (.A(_08408_),
    .B(_08528_),
    .Y(_08529_));
 AOI21x1_ASAP7_75t_R _16574_ (.A1(_08527_),
    .A2(_08529_),
    .B(net6333),
    .Y(_08530_));
 NOR2x1_ASAP7_75t_R _16575_ (.A(net6330),
    .B(net5028),
    .Y(_08531_));
 AO21x1_ASAP7_75t_R _16576_ (.A1(_08531_),
    .A2(net5246),
    .B(_08363_),
    .Y(_08532_));
 OA21x2_ASAP7_75t_R _16577_ (.A1(net4791),
    .A2(net6326),
    .B(net6334),
    .Y(_08533_));
 AO21x1_ASAP7_75t_R _16578_ (.A1(net5967),
    .A2(_08262_),
    .B(net6379),
    .Y(_08534_));
 AOI21x1_ASAP7_75t_R _16579_ (.A1(_08533_),
    .A2(_08534_),
    .B(net6332),
    .Y(_08535_));
 OAI21x1_ASAP7_75t_R _16580_ (.A1(net6334),
    .A2(_08532_),
    .B(_08535_),
    .Y(_08536_));
 AOI21x1_ASAP7_75t_R _16581_ (.A1(_08530_),
    .A2(_08536_),
    .B(_08182_),
    .Y(_08537_));
 OAI21x1_ASAP7_75t_R _16582_ (.A1(_08520_),
    .A2(_08525_),
    .B(_08537_),
    .Y(_08538_));
 OAI21x1_ASAP7_75t_R _16583_ (.A1(_08503_),
    .A2(_08513_),
    .B(_08538_),
    .Y(_00005_));
 AND3x1_ASAP7_75t_R _16584_ (.A(_08432_),
    .B(net6380),
    .C(net5970),
    .Y(_08539_));
 AO21x1_ASAP7_75t_R _16585_ (.A1(_00993_),
    .A2(_00994_),
    .B(net6378),
    .Y(_08540_));
 NAND2x1_ASAP7_75t_R _16586_ (.A(net5977),
    .B(_08540_),
    .Y(_08541_));
 AO21x1_ASAP7_75t_R _16587_ (.A1(net4978),
    .A2(_08262_),
    .B(net6326),
    .Y(_08542_));
 OA21x2_ASAP7_75t_R _16588_ (.A1(net4982),
    .A2(net6380),
    .B(net6334),
    .Y(_08543_));
 AOI21x1_ASAP7_75t_R _16589_ (.A1(_08542_),
    .A2(_08543_),
    .B(net5972),
    .Y(_08544_));
 OAI21x1_ASAP7_75t_R _16590_ (.A1(_08539_),
    .A2(_08541_),
    .B(_08544_),
    .Y(_08545_));
 AO21x1_ASAP7_75t_R _16591_ (.A1(_08263_),
    .A2(_08357_),
    .B(net6379),
    .Y(_08546_));
 AO21x1_ASAP7_75t_R _16592_ (.A1(_08138_),
    .A2(_08344_),
    .B(net6326),
    .Y(_08547_));
 AOI21x1_ASAP7_75t_R _16593_ (.A1(_08546_),
    .A2(_08547_),
    .B(net6335),
    .Y(_08548_));
 NAND2x1p5_ASAP7_75t_R _16594_ (.A(net4791),
    .B(_08208_),
    .Y(_08549_));
 AOI21x1_ASAP7_75t_R _16595_ (.A1(_08408_),
    .A2(_08549_),
    .B(net5979),
    .Y(_08550_));
 OAI21x1_ASAP7_75t_R _16596_ (.A1(_08550_),
    .A2(_08548_),
    .B(net5972),
    .Y(_08551_));
 AOI21x1_ASAP7_75t_R _16597_ (.A1(_08551_),
    .A2(_08545_),
    .B(_08121_),
    .Y(_08552_));
 OR3x1_ASAP7_75t_R _16598_ (.A(net6339),
    .B(net5242),
    .C(net6379),
    .Y(_08553_));
 AO21x1_ASAP7_75t_R _16599_ (.A1(net5248),
    .A2(net5970),
    .B(net6326),
    .Y(_08554_));
 AOI21x1_ASAP7_75t_R _16600_ (.A1(_08553_),
    .A2(_08554_),
    .B(net5979),
    .Y(_08555_));
 NAND2x1_ASAP7_75t_R _16601_ (.A(_08173_),
    .B(_08485_),
    .Y(_08556_));
 AOI21x1_ASAP7_75t_R _16602_ (.A1(_08549_),
    .A2(_08556_),
    .B(net6334),
    .Y(_08557_));
 OAI21x1_ASAP7_75t_R _16603_ (.A1(_08555_),
    .A2(_08557_),
    .B(net5972),
    .Y(_08558_));
 NAND2x1_ASAP7_75t_R _16604_ (.A(_08192_),
    .B(net4718),
    .Y(_08559_));
 AOI21x1_ASAP7_75t_R _16605_ (.A1(_08337_),
    .A2(_08559_),
    .B(net5976),
    .Y(_08560_));
 NOR2x1_ASAP7_75t_R _16606_ (.A(_08285_),
    .B(_08440_),
    .Y(_08561_));
 NOR2x1_ASAP7_75t_R _16607_ (.A(net5028),
    .B(_08446_),
    .Y(_08562_));
 OA21x2_ASAP7_75t_R _16608_ (.A1(_08561_),
    .A2(_08562_),
    .B(net5976),
    .Y(_08563_));
 OAI21x1_ASAP7_75t_R _16609_ (.A1(_08560_),
    .A2(_08563_),
    .B(net6333),
    .Y(_08564_));
 AOI21x1_ASAP7_75t_R _16610_ (.A1(_08558_),
    .A2(_08564_),
    .B(net6332),
    .Y(_08565_));
 OAI21x1_ASAP7_75t_R _16611_ (.A1(_08552_),
    .A2(_08565_),
    .B(_08097_),
    .Y(_08566_));
 AOI21x1_ASAP7_75t_R _16612_ (.A1(_08398_),
    .A2(_08471_),
    .B(net5978),
    .Y(_08567_));
 AND3x1_ASAP7_75t_R _16613_ (.A(net5248),
    .B(net6379),
    .C(_08289_),
    .Y(_08568_));
 OAI21x1_ASAP7_75t_R _16614_ (.A1(net6335),
    .A2(_08568_),
    .B(net5972),
    .Y(_08569_));
 OAI21x1_ASAP7_75t_R _16615_ (.A1(_08567_),
    .A2(_08569_),
    .B(_08121_),
    .Y(_08570_));
 AOI21x1_ASAP7_75t_R _16616_ (.A1(_00987_),
    .A2(net6380),
    .B(net6334),
    .Y(_08571_));
 NAND2x1_ASAP7_75t_R _16617_ (.A(_08571_),
    .B(_08510_),
    .Y(_08572_));
 AO21x1_ASAP7_75t_R _16618_ (.A1(_08371_),
    .A2(_08531_),
    .B(_08414_),
    .Y(_08573_));
 AOI21x1_ASAP7_75t_R _16619_ (.A1(_08572_),
    .A2(_08573_),
    .B(net5972),
    .Y(_08574_));
 NOR2x1_ASAP7_75t_R _16620_ (.A(_08570_),
    .B(_08574_),
    .Y(_08575_));
 AOI21x1_ASAP7_75t_R _16621_ (.A1(net5243),
    .A2(_08219_),
    .B(net5979),
    .Y(_08576_));
 NAND2x1_ASAP7_75t_R _16622_ (.A(net6330),
    .B(net5028),
    .Y(_08577_));
 AOI21x1_ASAP7_75t_R _16623_ (.A1(_08577_),
    .A2(_08408_),
    .B(net6334),
    .Y(_08578_));
 OAI21x1_ASAP7_75t_R _16624_ (.A1(_08576_),
    .A2(_08578_),
    .B(net5972),
    .Y(_08579_));
 AO21x1_ASAP7_75t_R _16625_ (.A1(net6339),
    .A2(net5322),
    .B(net6379),
    .Y(_08580_));
 AO21x1_ASAP7_75t_R _16626_ (.A1(_08131_),
    .A2(_08432_),
    .B(net6330),
    .Y(_08581_));
 AOI21x1_ASAP7_75t_R _16627_ (.A1(_08580_),
    .A2(_08581_),
    .B(_08414_),
    .Y(_08582_));
 AO21x1_ASAP7_75t_R _16628_ (.A1(_08233_),
    .A2(net5245),
    .B(net6379),
    .Y(_08583_));
 AO21x1_ASAP7_75t_R _16629_ (.A1(_08173_),
    .A2(_08207_),
    .B(net6330),
    .Y(_08584_));
 AOI21x1_ASAP7_75t_R _16630_ (.A1(_08583_),
    .A2(_08584_),
    .B(net6334),
    .Y(_08585_));
 OAI21x1_ASAP7_75t_R _16631_ (.A1(_08582_),
    .A2(_08585_),
    .B(net6333),
    .Y(_08586_));
 AOI21x1_ASAP7_75t_R _16632_ (.A1(_08579_),
    .A2(_08586_),
    .B(_08121_),
    .Y(_08587_));
 OAI21x1_ASAP7_75t_R _16633_ (.A1(_08575_),
    .A2(_08587_),
    .B(_08182_),
    .Y(_08588_));
 NAND2x1_ASAP7_75t_R _16634_ (.A(_08588_),
    .B(_08566_),
    .Y(_00006_));
 AO21x1_ASAP7_75t_R _16635_ (.A1(net4982),
    .A2(net5970),
    .B(net6326),
    .Y(_08589_));
 AO21x1_ASAP7_75t_R _16636_ (.A1(net4982),
    .A2(_08262_),
    .B(net6380),
    .Y(_08590_));
 AO21x1_ASAP7_75t_R _16637_ (.A1(_08589_),
    .A2(_08590_),
    .B(net6334),
    .Y(_08591_));
 OAI21x1_ASAP7_75t_R _16638_ (.A1(net5252),
    .A2(_08539_),
    .B(net6334),
    .Y(_08592_));
 NAND2x1_ASAP7_75t_R _16639_ (.A(_08591_),
    .B(_08592_),
    .Y(_08593_));
 AO21x1_ASAP7_75t_R _16640_ (.A1(net5967),
    .A2(_08344_),
    .B(net6379),
    .Y(_08594_));
 AO21x1_ASAP7_75t_R _16641_ (.A1(_08404_),
    .A2(_08594_),
    .B(net5978),
    .Y(_08595_));
 AO21x1_ASAP7_75t_R _16642_ (.A1(_08192_),
    .A2(net5250),
    .B(net6326),
    .Y(_08596_));
 AO21x1_ASAP7_75t_R _16643_ (.A1(net4982),
    .A2(_08344_),
    .B(net6377),
    .Y(_08597_));
 AO21x1_ASAP7_75t_R _16644_ (.A1(_08596_),
    .A2(_08597_),
    .B(net6335),
    .Y(_08598_));
 AOI21x1_ASAP7_75t_R _16645_ (.A1(_08595_),
    .A2(_08598_),
    .B(net5972),
    .Y(_08599_));
 AOI211x1_ASAP7_75t_R _16646_ (.A1(_08593_),
    .A2(net5972),
    .B(_08599_),
    .C(_08121_),
    .Y(_08600_));
 NAND2x1_ASAP7_75t_R _16647_ (.A(net6327),
    .B(_08296_),
    .Y(_08601_));
 OA21x2_ASAP7_75t_R _16648_ (.A1(net6327),
    .A2(_00993_),
    .B(_08117_),
    .Y(_08602_));
 AO31x2_ASAP7_75t_R _16649_ (.A1(_08601_),
    .A2(net4983),
    .A3(_08602_),
    .B(net6333),
    .Y(_08603_));
 INVx1_ASAP7_75t_R _16650_ (.A(_00991_),
    .Y(_08604_));
 AOI221x1_ASAP7_75t_R _16651_ (.A1(_08604_),
    .A2(net6328),
    .B1(net4601),
    .B2(_08531_),
    .C(_08414_),
    .Y(_08605_));
 AO21x1_ASAP7_75t_R _16652_ (.A1(net5248),
    .A2(net5969),
    .B(net6377),
    .Y(_08606_));
 NAND2x1_ASAP7_75t_R _16653_ (.A(_08243_),
    .B(_08606_),
    .Y(_08607_));
 NAND2x1_ASAP7_75t_R _16654_ (.A(net5323),
    .B(net6380),
    .Y(_08608_));
 OA21x2_ASAP7_75t_R _16655_ (.A1(_08262_),
    .A2(net6380),
    .B(_08608_),
    .Y(_08609_));
 AOI21x1_ASAP7_75t_R _16656_ (.A1(net5976),
    .A2(_08609_),
    .B(net5972),
    .Y(_08610_));
 OAI21x1_ASAP7_75t_R _16657_ (.A1(net5980),
    .A2(_08607_),
    .B(_08610_),
    .Y(_08611_));
 OAI21x1_ASAP7_75t_R _16658_ (.A1(_08603_),
    .A2(_08605_),
    .B(_08611_),
    .Y(_08612_));
 OAI21x1_ASAP7_75t_R _16659_ (.A1(net6332),
    .A2(_08612_),
    .B(_08097_),
    .Y(_08613_));
 AO21x1_ASAP7_75t_R _16660_ (.A1(_08321_),
    .A2(_08546_),
    .B(net6335),
    .Y(_08614_));
 AO21x1_ASAP7_75t_R _16661_ (.A1(_08388_),
    .A2(_08306_),
    .B(net5978),
    .Y(_08615_));
 AOI21x1_ASAP7_75t_R _16662_ (.A1(_08614_),
    .A2(_08615_),
    .B(net6333),
    .Y(_08616_));
 NOR2x1_ASAP7_75t_R _16663_ (.A(net6335),
    .B(_08480_),
    .Y(_08617_));
 AO21x1_ASAP7_75t_R _16664_ (.A1(_08471_),
    .A2(_08617_),
    .B(net5972),
    .Y(_08618_));
 OA22x2_ASAP7_75t_R _16665_ (.A1(net6327),
    .A2(net4982),
    .B1(_08223_),
    .B2(net5247),
    .Y(_08619_));
 OA21x2_ASAP7_75t_R _16666_ (.A1(net6331),
    .A2(_08104_),
    .B(net6336),
    .Y(_08620_));
 AND2x2_ASAP7_75t_R _16667_ (.A(_08619_),
    .B(_08620_),
    .Y(_08621_));
 OAI21x1_ASAP7_75t_R _16668_ (.A1(_08618_),
    .A2(_08621_),
    .B(net6332),
    .Y(_08622_));
 NOR2x1_ASAP7_75t_R _16669_ (.A(net5978),
    .B(_08485_),
    .Y(_08623_));
 AO21x1_ASAP7_75t_R _16670_ (.A1(_08192_),
    .A2(_08344_),
    .B(net6377),
    .Y(_08624_));
 NAND2x1_ASAP7_75t_R _16671_ (.A(_08624_),
    .B(_08623_),
    .Y(_08625_));
 OA21x2_ASAP7_75t_R _16672_ (.A1(net4719),
    .A2(_08394_),
    .B(net5972),
    .Y(_08626_));
 AOI21x1_ASAP7_75t_R _16673_ (.A1(_08626_),
    .A2(_08625_),
    .B(net6332),
    .Y(_08627_));
 AO21x1_ASAP7_75t_R _16674_ (.A1(_08366_),
    .A2(_08344_),
    .B(net6377),
    .Y(_08628_));
 AOI21x1_ASAP7_75t_R _16675_ (.A1(_08628_),
    .A2(_08331_),
    .B(net5972),
    .Y(_08629_));
 NOR2x1_ASAP7_75t_R _16676_ (.A(net6376),
    .B(net5981),
    .Y(_08630_));
 OAI21x1_ASAP7_75t_R _16677_ (.A1(_08630_),
    .A2(_08460_),
    .B(net6335),
    .Y(_08631_));
 NAND2x1_ASAP7_75t_R _16678_ (.A(_08629_),
    .B(_08631_),
    .Y(_08632_));
 AOI21x1_ASAP7_75t_R _16679_ (.A1(_08632_),
    .A2(_08627_),
    .B(_08097_),
    .Y(_08633_));
 OAI21x1_ASAP7_75t_R _16680_ (.A1(_08616_),
    .A2(_08622_),
    .B(_08633_),
    .Y(_08634_));
 OAI21x1_ASAP7_75t_R _16681_ (.A1(_08600_),
    .A2(_08613_),
    .B(_08634_),
    .Y(_00007_));
 XOR2x2_ASAP7_75t_R _16682_ (.A(net6540),
    .B(net6539),
    .Y(_08635_));
 AND2x2_ASAP7_75t_R _16687_ (.A(net6684),
    .B(net124),
    .Y(_08640_));
 AO21x1_ASAP7_75t_R _16688_ (.A1(_08635_),
    .A2(net6675),
    .B(_08640_),
    .Y(_00289_));
 XOR2x2_ASAP7_75t_R _16689_ (.A(_00422_),
    .B(net6529),
    .Y(_08641_));
 AND2x2_ASAP7_75t_R _16690_ (.A(net6684),
    .B(net125),
    .Y(_08642_));
 AO21x1_ASAP7_75t_R _16691_ (.A1(_08641_),
    .A2(net6675),
    .B(_08642_),
    .Y(_00300_));
 XOR2x2_ASAP7_75t_R _16692_ (.A(_00423_),
    .B(net6522),
    .Y(_08643_));
 AND2x2_ASAP7_75t_R _16693_ (.A(net6684),
    .B(net126),
    .Y(_08644_));
 AO21x1_ASAP7_75t_R _16694_ (.A1(_08643_),
    .A2(net6674),
    .B(_08644_),
    .Y(_00311_));
 XOR2x2_ASAP7_75t_R _16695_ (.A(_00424_),
    .B(net6519),
    .Y(_08645_));
 AND2x2_ASAP7_75t_R _16696_ (.A(net6684),
    .B(net127),
    .Y(_08646_));
 AO21x1_ASAP7_75t_R _16697_ (.A1(_08645_),
    .A2(net6675),
    .B(_08646_),
    .Y(_00314_));
 XOR2x2_ASAP7_75t_R _16698_ (.A(_00425_),
    .B(_00864_),
    .Y(_08647_));
 AND2x2_ASAP7_75t_R _16699_ (.A(net6684),
    .B(net2),
    .Y(_08648_));
 AO21x1_ASAP7_75t_R _16700_ (.A1(_08647_),
    .A2(net6675),
    .B(_08648_),
    .Y(_00315_));
 XOR2x2_ASAP7_75t_R _16701_ (.A(_00426_),
    .B(_00865_),
    .Y(_08649_));
 AND2x2_ASAP7_75t_R _16702_ (.A(net6686),
    .B(net3),
    .Y(_08650_));
 AO21x1_ASAP7_75t_R _16703_ (.A1(_08649_),
    .A2(net6675),
    .B(_08650_),
    .Y(_00316_));
 XOR2x2_ASAP7_75t_R _16704_ (.A(_00427_),
    .B(_00866_),
    .Y(_08651_));
 AND2x2_ASAP7_75t_R _16706_ (.A(net6684),
    .B(net4),
    .Y(_08653_));
 AO21x1_ASAP7_75t_R _16707_ (.A1(_08651_),
    .A2(net6675),
    .B(_08653_),
    .Y(_00317_));
 XOR2x2_ASAP7_75t_R _16708_ (.A(_00428_),
    .B(_00867_),
    .Y(_08654_));
 AND2x2_ASAP7_75t_R _16710_ (.A(net6684),
    .B(net5),
    .Y(_08656_));
 AO21x1_ASAP7_75t_R _16711_ (.A1(_08654_),
    .A2(net6675),
    .B(_08656_),
    .Y(_00318_));
 XOR2x2_ASAP7_75t_R _16712_ (.A(net6541),
    .B(net6514),
    .Y(_08657_));
 AND2x2_ASAP7_75t_R _16713_ (.A(net6680),
    .B(net6),
    .Y(_08658_));
 AO21x1_ASAP7_75t_R _16714_ (.A1(_08657_),
    .A2(net6674),
    .B(_08658_),
    .Y(_00319_));
 XOR2x2_ASAP7_75t_R _16715_ (.A(_00430_),
    .B(net6513),
    .Y(_08659_));
 AND2x2_ASAP7_75t_R _16716_ (.A(net6680),
    .B(net7),
    .Y(_08660_));
 AO21x1_ASAP7_75t_R _16717_ (.A1(_08659_),
    .A2(net6674),
    .B(_08660_),
    .Y(_00320_));
 XOR2x2_ASAP7_75t_R _16718_ (.A(_00431_),
    .B(net6538),
    .Y(_08661_));
 AND2x2_ASAP7_75t_R _16719_ (.A(net6680),
    .B(net8),
    .Y(_08662_));
 AO21x1_ASAP7_75t_R _16720_ (.A1(_08661_),
    .A2(net6674),
    .B(_08662_),
    .Y(_00290_));
 XOR2x2_ASAP7_75t_R _16721_ (.A(_00432_),
    .B(net6537),
    .Y(_08663_));
 AND2x2_ASAP7_75t_R _16722_ (.A(net6680),
    .B(net9),
    .Y(_08664_));
 AO21x1_ASAP7_75t_R _16723_ (.A1(_08663_),
    .A2(net6674),
    .B(_08664_),
    .Y(_00291_));
 XOR2x2_ASAP7_75t_R _16724_ (.A(_00433_),
    .B(_00841_),
    .Y(_08665_));
 AND2x2_ASAP7_75t_R _16725_ (.A(net6680),
    .B(net10),
    .Y(_08666_));
 AO21x1_ASAP7_75t_R _16726_ (.A1(_08665_),
    .A2(net6674),
    .B(_08666_),
    .Y(_00292_));
 XOR2x2_ASAP7_75t_R _16727_ (.A(_00434_),
    .B(_00842_),
    .Y(_08667_));
 AND2x2_ASAP7_75t_R _16728_ (.A(net6680),
    .B(net11),
    .Y(_08668_));
 AO21x1_ASAP7_75t_R _16729_ (.A1(_08667_),
    .A2(net6674),
    .B(_08668_),
    .Y(_00293_));
 XOR2x2_ASAP7_75t_R _16730_ (.A(_00435_),
    .B(_00843_),
    .Y(_08669_));
 AND2x2_ASAP7_75t_R _16731_ (.A(net6680),
    .B(net13),
    .Y(_08670_));
 AO21x1_ASAP7_75t_R _16732_ (.A1(_08669_),
    .A2(net6674),
    .B(_08670_),
    .Y(_00294_));
 XOR2x2_ASAP7_75t_R _16733_ (.A(_00436_),
    .B(_00844_),
    .Y(_08671_));
 AND2x2_ASAP7_75t_R _16734_ (.A(net6683),
    .B(net14),
    .Y(_08672_));
 AO21x1_ASAP7_75t_R _16735_ (.A1(_08671_),
    .A2(net6674),
    .B(_08672_),
    .Y(_00295_));
 XNOR2x2_ASAP7_75t_R _16739_ (.A(_00437_),
    .B(net6533),
    .Y(_08676_));
 NOR2x1_ASAP7_75t_R _16740_ (.A(net6688),
    .B(_08676_),
    .Y(_08677_));
 AO21x1_ASAP7_75t_R _16741_ (.A1(net6688),
    .A2(net15),
    .B(_08677_),
    .Y(_00296_));
 XNOR2x2_ASAP7_75t_R _16743_ (.A(_00438_),
    .B(net6532),
    .Y(_08679_));
 NOR2x1_ASAP7_75t_R _16744_ (.A(net6688),
    .B(_08679_),
    .Y(_08680_));
 AO21x1_ASAP7_75t_R _16745_ (.A1(net6688),
    .A2(net16),
    .B(_08680_),
    .Y(_00297_));
 AND2x2_ASAP7_75t_R _16747_ (.A(net6684),
    .B(net17),
    .Y(_08682_));
 AO21x1_ASAP7_75t_R _16748_ (.A1(_08052_),
    .A2(net6677),
    .B(_08682_),
    .Y(_00298_));
 XNOR2x2_ASAP7_75t_R _16749_ (.A(_00439_),
    .B(net6530),
    .Y(_08683_));
 NOR2x1_ASAP7_75t_R _16750_ (.A(net6688),
    .B(_08683_),
    .Y(_08684_));
 AO21x1_ASAP7_75t_R _16751_ (.A1(net6688),
    .A2(net18),
    .B(_08684_),
    .Y(_00299_));
 XNOR2x2_ASAP7_75t_R _16752_ (.A(_00440_),
    .B(_00850_),
    .Y(_08685_));
 NOR2x1_ASAP7_75t_R _16753_ (.A(net6682),
    .B(_08685_),
    .Y(_08686_));
 AO21x1_ASAP7_75t_R _16754_ (.A1(net6682),
    .A2(net19),
    .B(_08686_),
    .Y(_00301_));
 XNOR2x2_ASAP7_75t_R _16755_ (.A(_00441_),
    .B(_00851_),
    .Y(_08687_));
 NOR2x1_ASAP7_75t_R _16756_ (.A(net6688),
    .B(_08687_),
    .Y(_08688_));
 AO21x1_ASAP7_75t_R _16757_ (.A1(net6688),
    .A2(net20),
    .B(_08688_),
    .Y(_00302_));
 XNOR2x2_ASAP7_75t_R _16758_ (.A(_00442_),
    .B(_00852_),
    .Y(_08689_));
 NOR2x1_ASAP7_75t_R _16759_ (.A(net6682),
    .B(_08689_),
    .Y(_08690_));
 AO21x1_ASAP7_75t_R _16760_ (.A1(net6682),
    .A2(net21),
    .B(_08690_),
    .Y(_00303_));
 XNOR2x2_ASAP7_75t_R _16761_ (.A(_00443_),
    .B(_00853_),
    .Y(_08691_));
 NOR2x1_ASAP7_75t_R _16762_ (.A(net6689),
    .B(_08691_),
    .Y(_08692_));
 AO21x1_ASAP7_75t_R _16763_ (.A1(net6689),
    .A2(net22),
    .B(_08692_),
    .Y(_00304_));
 XOR2x2_ASAP7_75t_R _16766_ (.A(_00830_),
    .B(_00854_),
    .Y(_08695_));
 XOR2x2_ASAP7_75t_R _16767_ (.A(_08695_),
    .B(_00413_),
    .Y(_08696_));
 NOR2x1_ASAP7_75t_R _16768_ (.A(net6688),
    .B(_08696_),
    .Y(_08697_));
 AO21x1_ASAP7_75t_R _16769_ (.A1(net6688),
    .A2(net24),
    .B(_08697_),
    .Y(_00305_));
 XOR2x2_ASAP7_75t_R _16770_ (.A(_00831_),
    .B(net6527),
    .Y(_08698_));
 XOR2x2_ASAP7_75t_R _16771_ (.A(_08698_),
    .B(_00414_),
    .Y(_08699_));
 NOR2x1_ASAP7_75t_R _16772_ (.A(net6688),
    .B(_08699_),
    .Y(_08700_));
 AO21x1_ASAP7_75t_R _16773_ (.A1(net6688),
    .A2(net25),
    .B(_08700_),
    .Y(_00306_));
 XOR2x2_ASAP7_75t_R _16774_ (.A(_00832_),
    .B(_00856_),
    .Y(_08701_));
 XOR2x2_ASAP7_75t_R _16775_ (.A(_08701_),
    .B(_00415_),
    .Y(_08702_));
 NOR2x1_ASAP7_75t_R _16776_ (.A(net6688),
    .B(_08702_),
    .Y(_08703_));
 AO21x1_ASAP7_75t_R _16777_ (.A1(net6688),
    .A2(net26),
    .B(_08703_),
    .Y(_00307_));
 XOR2x2_ASAP7_75t_R _16778_ (.A(_00833_),
    .B(net6525),
    .Y(_08704_));
 XOR2x2_ASAP7_75t_R _16779_ (.A(_08704_),
    .B(_00416_),
    .Y(_08705_));
 NOR2x1_ASAP7_75t_R _16780_ (.A(net6688),
    .B(_08705_),
    .Y(_08706_));
 AO21x1_ASAP7_75t_R _16781_ (.A1(net6688),
    .A2(net27),
    .B(_08706_),
    .Y(_00308_));
 XOR2x2_ASAP7_75t_R _16783_ (.A(_00834_),
    .B(_00858_),
    .Y(_08708_));
 XOR2x2_ASAP7_75t_R _16784_ (.A(_08708_),
    .B(_00417_),
    .Y(_08709_));
 NOR2x1_ASAP7_75t_R _16785_ (.A(net6688),
    .B(_08709_),
    .Y(_08710_));
 AO21x1_ASAP7_75t_R _16786_ (.A1(net6688),
    .A2(net28),
    .B(_08710_),
    .Y(_00309_));
 XOR2x2_ASAP7_75t_R _16787_ (.A(_00835_),
    .B(_00859_),
    .Y(_08711_));
 XOR2x2_ASAP7_75t_R _16788_ (.A(_08711_),
    .B(_00418_),
    .Y(_08712_));
 NOR2x1_ASAP7_75t_R _16789_ (.A(net6688),
    .B(_08712_),
    .Y(_08713_));
 AO21x1_ASAP7_75t_R _16790_ (.A1(net6688),
    .A2(net29),
    .B(_08713_),
    .Y(_00310_));
 XOR2x2_ASAP7_75t_R _16791_ (.A(_00836_),
    .B(_00861_),
    .Y(_08714_));
 XOR2x2_ASAP7_75t_R _16792_ (.A(_08714_),
    .B(_00419_),
    .Y(_08715_));
 NOR2x1_ASAP7_75t_R _16793_ (.A(net6688),
    .B(_08715_),
    .Y(_08716_));
 AO21x1_ASAP7_75t_R _16794_ (.A1(net6688),
    .A2(net30),
    .B(_08716_),
    .Y(_00312_));
 XOR2x2_ASAP7_75t_R _16795_ (.A(_00837_),
    .B(_00862_),
    .Y(_08717_));
 XOR2x2_ASAP7_75t_R _16796_ (.A(_08717_),
    .B(_00420_),
    .Y(_08718_));
 NOR2x1_ASAP7_75t_R _16797_ (.A(net6688),
    .B(_08718_),
    .Y(_08719_));
 AO21x1_ASAP7_75t_R _16798_ (.A1(net6688),
    .A2(net31),
    .B(_08719_),
    .Y(_00313_));
 XOR2x2_ASAP7_75t_R _16799_ (.A(_00838_),
    .B(_00870_),
    .Y(_08720_));
 XOR2x2_ASAP7_75t_R _16800_ (.A(net6471),
    .B(net6540),
    .Y(_08721_));
 NOR2x1_ASAP7_75t_R _16801_ (.A(net6686),
    .B(_08721_),
    .Y(_08722_));
 AO21x1_ASAP7_75t_R _16802_ (.A1(net6686),
    .A2(net89),
    .B(_08722_),
    .Y(_00321_));
 XOR2x2_ASAP7_75t_R _16803_ (.A(_00881_),
    .B(_00849_),
    .Y(_08723_));
 XOR2x2_ASAP7_75t_R _16804_ (.A(net6470),
    .B(_00422_),
    .Y(_08724_));
 NOR2x1_ASAP7_75t_R _16805_ (.A(net6684),
    .B(_08724_),
    .Y(_08725_));
 AO21x1_ASAP7_75t_R _16806_ (.A1(net6684),
    .A2(net90),
    .B(_08725_),
    .Y(_00332_));
 XOR2x2_ASAP7_75t_R _16808_ (.A(_00860_),
    .B(_00892_),
    .Y(_08727_));
 XOR2x2_ASAP7_75t_R _16809_ (.A(_08727_),
    .B(_00423_),
    .Y(_08728_));
 NOR2x1_ASAP7_75t_R _16810_ (.A(net6683),
    .B(_08728_),
    .Y(_08729_));
 AO21x1_ASAP7_75t_R _16811_ (.A1(net6683),
    .A2(net91),
    .B(_08729_),
    .Y(_00343_));
 XOR2x2_ASAP7_75t_R _16812_ (.A(_00863_),
    .B(_00895_),
    .Y(_08730_));
 XOR2x2_ASAP7_75t_R _16813_ (.A(_08730_),
    .B(_00424_),
    .Y(_08731_));
 NOR2x1_ASAP7_75t_R _16814_ (.A(net6684),
    .B(_08731_),
    .Y(_08732_));
 AO21x1_ASAP7_75t_R _16815_ (.A1(net6684),
    .A2(net92),
    .B(_08732_),
    .Y(_00346_));
 XOR2x2_ASAP7_75t_R _16816_ (.A(_08647_),
    .B(net6497),
    .Y(_08733_));
 NOR2x1_ASAP7_75t_R _16817_ (.A(net6684),
    .B(_08733_),
    .Y(_08734_));
 AO21x1_ASAP7_75t_R _16818_ (.A1(net6684),
    .A2(net93),
    .B(_08734_),
    .Y(_00347_));
 XOR2x2_ASAP7_75t_R _16819_ (.A(_08649_),
    .B(net6496),
    .Y(_08735_));
 NOR2x1_ASAP7_75t_R _16820_ (.A(net6686),
    .B(_08735_),
    .Y(_08736_));
 AO21x1_ASAP7_75t_R _16821_ (.A1(net6686),
    .A2(net94),
    .B(_08736_),
    .Y(_00348_));
 XOR2x2_ASAP7_75t_R _16823_ (.A(_08651_),
    .B(_00898_),
    .Y(_08738_));
 NOR2x1_ASAP7_75t_R _16824_ (.A(net6686),
    .B(_08738_),
    .Y(_08739_));
 AO21x1_ASAP7_75t_R _16825_ (.A1(net6686),
    .A2(net96),
    .B(_08739_),
    .Y(_00349_));
 XOR2x2_ASAP7_75t_R _16826_ (.A(_08654_),
    .B(_00899_),
    .Y(_08740_));
 NOR2x1_ASAP7_75t_R _16827_ (.A(net6684),
    .B(_08740_),
    .Y(_08741_));
 AO21x1_ASAP7_75t_R _16828_ (.A1(net6684),
    .A2(net97),
    .B(_08741_),
    .Y(_00350_));
 XOR2x2_ASAP7_75t_R _16829_ (.A(_00868_),
    .B(_00900_),
    .Y(_08742_));
 XOR2x2_ASAP7_75t_R _16830_ (.A(net6469),
    .B(net6541),
    .Y(_08743_));
 NOR2x1_ASAP7_75t_R _16831_ (.A(net6683),
    .B(_08743_),
    .Y(_08744_));
 AO21x1_ASAP7_75t_R _16832_ (.A1(net6683),
    .A2(net98),
    .B(_08744_),
    .Y(_00351_));
 INVx1_ASAP7_75t_R _16834_ (.A(net6493),
    .Y(_08746_));
 OA21x2_ASAP7_75t_R _16835_ (.A1(_08659_),
    .A2(_08746_),
    .B(net6677),
    .Y(_08747_));
 NAND2x1_ASAP7_75t_R _16836_ (.A(_08746_),
    .B(_08659_),
    .Y(_08748_));
 AO22x1_ASAP7_75t_R _16837_ (.A1(net6683),
    .A2(net99),
    .B1(_08747_),
    .B2(_08748_),
    .Y(_00352_));
 XOR2x2_ASAP7_75t_R _16838_ (.A(_00839_),
    .B(_00871_),
    .Y(_08749_));
 XOR2x2_ASAP7_75t_R _16839_ (.A(_08749_),
    .B(_00431_),
    .Y(_08750_));
 NOR2x1_ASAP7_75t_R _16840_ (.A(net6683),
    .B(_08750_),
    .Y(_08751_));
 AO21x1_ASAP7_75t_R _16841_ (.A1(net6683),
    .A2(net100),
    .B(_08751_),
    .Y(_00322_));
 XOR2x2_ASAP7_75t_R _16842_ (.A(_00840_),
    .B(_00872_),
    .Y(_08752_));
 XOR2x2_ASAP7_75t_R _16843_ (.A(_08752_),
    .B(_00432_),
    .Y(_08753_));
 NOR2x1_ASAP7_75t_R _16844_ (.A(net6683),
    .B(_08753_),
    .Y(_08754_));
 AO21x1_ASAP7_75t_R _16845_ (.A1(net6683),
    .A2(net101),
    .B(_08754_),
    .Y(_00323_));
 XOR2x2_ASAP7_75t_R _16846_ (.A(_08665_),
    .B(_00873_),
    .Y(_08755_));
 NOR2x1_ASAP7_75t_R _16847_ (.A(net6683),
    .B(_08755_),
    .Y(_08756_));
 AO21x1_ASAP7_75t_R _16848_ (.A1(net6683),
    .A2(net102),
    .B(_08756_),
    .Y(_00324_));
 XOR2x2_ASAP7_75t_R _16850_ (.A(_08667_),
    .B(_00874_),
    .Y(_08758_));
 NOR2x1_ASAP7_75t_R _16851_ (.A(net6683),
    .B(_08758_),
    .Y(_08759_));
 AO21x1_ASAP7_75t_R _16852_ (.A1(net6683),
    .A2(net103),
    .B(_08759_),
    .Y(_00325_));
 XOR2x2_ASAP7_75t_R _16853_ (.A(_08669_),
    .B(_00875_),
    .Y(_08760_));
 NOR2x1_ASAP7_75t_R _16854_ (.A(net6683),
    .B(_08760_),
    .Y(_08761_));
 AO21x1_ASAP7_75t_R _16855_ (.A1(net6683),
    .A2(net104),
    .B(_08761_),
    .Y(_00326_));
 XOR2x2_ASAP7_75t_R _16856_ (.A(_08671_),
    .B(_00876_),
    .Y(_08762_));
 NOR2x1_ASAP7_75t_R _16857_ (.A(net6683),
    .B(_08762_),
    .Y(_08763_));
 AO21x1_ASAP7_75t_R _16858_ (.A1(net6683),
    .A2(net105),
    .B(_08763_),
    .Y(_00327_));
 INVx1_ASAP7_75t_R _16859_ (.A(net6508),
    .Y(_08764_));
 XOR2x2_ASAP7_75t_R _16860_ (.A(_08676_),
    .B(_08764_),
    .Y(_08765_));
 NOR2x1_ASAP7_75t_R _16861_ (.A(net6688),
    .B(_08765_),
    .Y(_08766_));
 AO21x1_ASAP7_75t_R _16862_ (.A1(net6688),
    .A2(net107),
    .B(_08766_),
    .Y(_00328_));
 INVx1_ASAP7_75t_R _16864_ (.A(net6507),
    .Y(_08768_));
 XOR2x2_ASAP7_75t_R _16865_ (.A(_08679_),
    .B(_08768_),
    .Y(_08769_));
 NOR2x1_ASAP7_75t_R _16866_ (.A(net6688),
    .B(_08769_),
    .Y(_08770_));
 AO21x1_ASAP7_75t_R _16867_ (.A1(net6688),
    .A2(net108),
    .B(_08770_),
    .Y(_00329_));
 INVx1_ASAP7_75t_R _16868_ (.A(net6506),
    .Y(_08771_));
 XOR2x2_ASAP7_75t_R _16869_ (.A(_08052_),
    .B(_08771_),
    .Y(_08772_));
 AND2x2_ASAP7_75t_R _16871_ (.A(net6689),
    .B(net109),
    .Y(_08774_));
 AO21x1_ASAP7_75t_R _16872_ (.A1(_08772_),
    .A2(net6678),
    .B(_08774_),
    .Y(_00330_));
 INVx1_ASAP7_75t_R _16873_ (.A(_00880_),
    .Y(_08775_));
 XOR2x2_ASAP7_75t_R _16874_ (.A(_08683_),
    .B(_08775_),
    .Y(_08776_));
 NOR2x1_ASAP7_75t_R _16875_ (.A(net6688),
    .B(_08776_),
    .Y(_08777_));
 AO21x1_ASAP7_75t_R _16876_ (.A1(net6688),
    .A2(net110),
    .B(_08777_),
    .Y(_00331_));
 INVx1_ASAP7_75t_R _16877_ (.A(_00882_),
    .Y(_08778_));
 XOR2x2_ASAP7_75t_R _16878_ (.A(_08685_),
    .B(_08778_),
    .Y(_08779_));
 NOR2x1_ASAP7_75t_R _16879_ (.A(net6682),
    .B(_08779_),
    .Y(_08780_));
 AO21x1_ASAP7_75t_R _16880_ (.A1(net6682),
    .A2(net111),
    .B(_08780_),
    .Y(_00333_));
 XNOR2x2_ASAP7_75t_R _16881_ (.A(_00883_),
    .B(_08687_),
    .Y(_08781_));
 NOR2x1_ASAP7_75t_R _16882_ (.A(net6688),
    .B(_08781_),
    .Y(_08782_));
 AO21x1_ASAP7_75t_R _16883_ (.A1(net6688),
    .A2(net112),
    .B(_08782_),
    .Y(_00334_));
 XNOR2x2_ASAP7_75t_R _16884_ (.A(_00884_),
    .B(_08689_),
    .Y(_08783_));
 NOR2x1_ASAP7_75t_R _16885_ (.A(net6682),
    .B(_08783_),
    .Y(_08784_));
 AO21x1_ASAP7_75t_R _16886_ (.A1(net6682),
    .A2(net113),
    .B(_08784_),
    .Y(_00335_));
 XNOR2x2_ASAP7_75t_R _16887_ (.A(net6504),
    .B(_08691_),
    .Y(_08785_));
 NOR2x1_ASAP7_75t_R _16888_ (.A(net6689),
    .B(_08785_),
    .Y(_08786_));
 AO21x1_ASAP7_75t_R _16889_ (.A1(net6689),
    .A2(net114),
    .B(_08786_),
    .Y(_00336_));
 XOR2x2_ASAP7_75t_R _16890_ (.A(net6503),
    .B(_08696_),
    .Y(_08787_));
 AND2x2_ASAP7_75t_R _16891_ (.A(net6688),
    .B(net115),
    .Y(_08788_));
 AO21x1_ASAP7_75t_R _16892_ (.A1(net6383),
    .A2(net6678),
    .B(_08788_),
    .Y(_00337_));
 INVx1_ASAP7_75t_R _16893_ (.A(_00414_),
    .Y(_08789_));
 XOR2x2_ASAP7_75t_R _16894_ (.A(_00887_),
    .B(_00855_),
    .Y(_08790_));
 XNOR2x2_ASAP7_75t_R _16895_ (.A(_08790_),
    .B(_00831_),
    .Y(_08791_));
 NAND2x1p5_ASAP7_75t_R _16896_ (.A(_08791_),
    .B(_08789_),
    .Y(_08792_));
 XOR2x2_ASAP7_75t_R _16897_ (.A(_08790_),
    .B(_00831_),
    .Y(_08793_));
 NAND2x1_ASAP7_75t_R _16898_ (.A(_00414_),
    .B(_08793_),
    .Y(_08794_));
 AND3x1_ASAP7_75t_R _16899_ (.A(_08792_),
    .B(_08794_),
    .C(net6678),
    .Y(_08795_));
 AO21x1_ASAP7_75t_R _16900_ (.A1(net6688),
    .A2(net116),
    .B(_08795_),
    .Y(_00338_));
 INVx1_ASAP7_75t_R _16902_ (.A(_00888_),
    .Y(_08797_));
 XOR2x2_ASAP7_75t_R _16903_ (.A(_08702_),
    .B(_08797_),
    .Y(_08798_));
 NOR2x1_ASAP7_75t_R _16904_ (.A(net6688),
    .B(_08798_),
    .Y(_08799_));
 AO21x1_ASAP7_75t_R _16905_ (.A1(net6688),
    .A2(net118),
    .B(_08799_),
    .Y(_00339_));
 XOR2x2_ASAP7_75t_R _16906_ (.A(_00857_),
    .B(_00889_),
    .Y(_08800_));
 XOR2x2_ASAP7_75t_R _16907_ (.A(_08800_),
    .B(_00833_),
    .Y(_08801_));
 NOR2x1_ASAP7_75t_R _16908_ (.A(_00416_),
    .B(_08801_),
    .Y(_08802_));
 INVx1_ASAP7_75t_R _16909_ (.A(_00416_),
    .Y(_08803_));
 XNOR2x2_ASAP7_75t_R _16910_ (.A(_00833_),
    .B(_08800_),
    .Y(_08804_));
 NOR2x1_ASAP7_75t_R _16911_ (.A(_08803_),
    .B(_08804_),
    .Y(_08805_));
 NOR2x1_ASAP7_75t_R _16912_ (.A(_08802_),
    .B(_08805_),
    .Y(_08806_));
 AND2x2_ASAP7_75t_R _16913_ (.A(net6689),
    .B(net119),
    .Y(_08807_));
 AO21x1_ASAP7_75t_R _16914_ (.A1(_08806_),
    .A2(net6678),
    .B(_08807_),
    .Y(_00340_));
 XOR2x2_ASAP7_75t_R _16915_ (.A(_08709_),
    .B(_00890_),
    .Y(_08808_));
 AND2x2_ASAP7_75t_R _16916_ (.A(net6688),
    .B(net120),
    .Y(_08809_));
 AO21x1_ASAP7_75t_R _16917_ (.A1(_08808_),
    .A2(net6678),
    .B(_08809_),
    .Y(_00341_));
 XOR2x2_ASAP7_75t_R _16918_ (.A(_08712_),
    .B(_00891_),
    .Y(_08810_));
 AND2x2_ASAP7_75t_R _16919_ (.A(net6688),
    .B(net121),
    .Y(_08811_));
 AO21x1_ASAP7_75t_R _16920_ (.A1(_08810_),
    .A2(net6678),
    .B(_08811_),
    .Y(_00342_));
 XOR2x2_ASAP7_75t_R _16921_ (.A(_08715_),
    .B(_00893_),
    .Y(_08812_));
 AND2x2_ASAP7_75t_R _16922_ (.A(net6688),
    .B(net122),
    .Y(_08813_));
 AO21x1_ASAP7_75t_R _16923_ (.A1(_08812_),
    .A2(net6678),
    .B(_08813_),
    .Y(_00344_));
 XOR2x2_ASAP7_75t_R _16924_ (.A(_08718_),
    .B(_00894_),
    .Y(_08814_));
 AND2x2_ASAP7_75t_R _16925_ (.A(net6688),
    .B(net123),
    .Y(_08815_));
 AO21x1_ASAP7_75t_R _16926_ (.A1(_08814_),
    .A2(net6678),
    .B(_08815_),
    .Y(_00345_));
 XOR2x2_ASAP7_75t_R _16927_ (.A(_00421_),
    .B(_00902_),
    .Y(_08816_));
 XOR2x2_ASAP7_75t_R _16928_ (.A(_08720_),
    .B(_08816_),
    .Y(_08817_));
 AND2x2_ASAP7_75t_R _16929_ (.A(net6684),
    .B(net54),
    .Y(_08818_));
 AO21x1_ASAP7_75t_R _16930_ (.A1(net6389),
    .A2(net6675),
    .B(_08818_),
    .Y(_00353_));
 XOR2x2_ASAP7_75t_R _16931_ (.A(_00422_),
    .B(_00913_),
    .Y(_08819_));
 XOR2x2_ASAP7_75t_R _16932_ (.A(_08723_),
    .B(_08819_),
    .Y(_08820_));
 AND2x2_ASAP7_75t_R _16933_ (.A(net6684),
    .B(net55),
    .Y(_08821_));
 AO21x1_ASAP7_75t_R _16934_ (.A1(_08820_),
    .A2(net6675),
    .B(_08821_),
    .Y(_00364_));
 INVx1_ASAP7_75t_R _16935_ (.A(net6480),
    .Y(_08822_));
 AO21x1_ASAP7_75t_R _16936_ (.A1(_08728_),
    .A2(_08822_),
    .B(net6683),
    .Y(_08823_));
 NOR2x1_ASAP7_75t_R _16937_ (.A(_08822_),
    .B(_08728_),
    .Y(_08824_));
 OA22x2_ASAP7_75t_R _16938_ (.A1(net6674),
    .A2(net56),
    .B1(_08823_),
    .B2(_08824_),
    .Y(_00375_));
 XOR2x2_ASAP7_75t_R _16939_ (.A(_00424_),
    .B(_00927_),
    .Y(_08825_));
 XOR2x2_ASAP7_75t_R _16940_ (.A(_08730_),
    .B(_08825_),
    .Y(_08826_));
 AND2x2_ASAP7_75t_R _16942_ (.A(net6684),
    .B(net57),
    .Y(_08828_));
 AO21x1_ASAP7_75t_R _16943_ (.A1(_08826_),
    .A2(net6675),
    .B(_08828_),
    .Y(_00378_));
 XOR2x2_ASAP7_75t_R _16944_ (.A(_08733_),
    .B(_00928_),
    .Y(_08829_));
 AND2x2_ASAP7_75t_R _16946_ (.A(net6684),
    .B(net58),
    .Y(_08831_));
 AO21x1_ASAP7_75t_R _16947_ (.A1(_08829_),
    .A2(_08030_),
    .B(_08831_),
    .Y(_00379_));
 XOR2x2_ASAP7_75t_R _16948_ (.A(_08735_),
    .B(_00929_),
    .Y(_08832_));
 AND2x2_ASAP7_75t_R _16949_ (.A(net6684),
    .B(net59),
    .Y(_08833_));
 AO21x1_ASAP7_75t_R _16950_ (.A1(_08832_),
    .A2(net6675),
    .B(_08833_),
    .Y(_00380_));
 XOR2x2_ASAP7_75t_R _16951_ (.A(_08738_),
    .B(_00930_),
    .Y(_08834_));
 AND2x2_ASAP7_75t_R _16952_ (.A(net6684),
    .B(net60),
    .Y(_08835_));
 AO21x1_ASAP7_75t_R _16953_ (.A1(_08834_),
    .A2(_08030_),
    .B(_08835_),
    .Y(_00381_));
 XOR2x2_ASAP7_75t_R _16954_ (.A(_08740_),
    .B(_00931_),
    .Y(_08836_));
 AND2x2_ASAP7_75t_R _16955_ (.A(net6684),
    .B(net61),
    .Y(_08837_));
 AO21x1_ASAP7_75t_R _16956_ (.A1(_08836_),
    .A2(net6675),
    .B(_08837_),
    .Y(_00382_));
 XOR2x2_ASAP7_75t_R _16957_ (.A(_00429_),
    .B(_00932_),
    .Y(_08838_));
 XOR2x2_ASAP7_75t_R _16958_ (.A(_08742_),
    .B(_08838_),
    .Y(_08839_));
 AND2x2_ASAP7_75t_R _16959_ (.A(net6683),
    .B(net63),
    .Y(_08840_));
 AO21x1_ASAP7_75t_R _16960_ (.A1(_08839_),
    .A2(net6674),
    .B(_08840_),
    .Y(_00383_));
 XOR2x2_ASAP7_75t_R _16961_ (.A(_00901_),
    .B(_00933_),
    .Y(_08841_));
 XOR2x2_ASAP7_75t_R _16962_ (.A(_08659_),
    .B(net6468),
    .Y(_08842_));
 AND2x2_ASAP7_75t_R _16963_ (.A(net6680),
    .B(net64),
    .Y(_08843_));
 AO21x1_ASAP7_75t_R _16964_ (.A1(_08842_),
    .A2(net6674),
    .B(_08843_),
    .Y(_00384_));
 INVx1_ASAP7_75t_R _16965_ (.A(net6491),
    .Y(_08844_));
 AO21x1_ASAP7_75t_R _16966_ (.A1(_08750_),
    .A2(_08844_),
    .B(net6683),
    .Y(_08845_));
 NOR2x1_ASAP7_75t_R _16967_ (.A(_08844_),
    .B(_08750_),
    .Y(_08846_));
 OA22x2_ASAP7_75t_R _16968_ (.A1(net6674),
    .A2(net65),
    .B1(_08845_),
    .B2(_08846_),
    .Y(_00354_));
 XOR2x2_ASAP7_75t_R _16969_ (.A(_00432_),
    .B(_00904_),
    .Y(_08847_));
 XOR2x2_ASAP7_75t_R _16970_ (.A(_08752_),
    .B(_08847_),
    .Y(_08848_));
 AND2x2_ASAP7_75t_R _16971_ (.A(net6680),
    .B(net66),
    .Y(_08849_));
 AO21x1_ASAP7_75t_R _16972_ (.A1(_08848_),
    .A2(net6674),
    .B(_08849_),
    .Y(_00355_));
 XOR2x2_ASAP7_75t_R _16973_ (.A(_08755_),
    .B(_00905_),
    .Y(_08850_));
 AND2x2_ASAP7_75t_R _16974_ (.A(net6683),
    .B(net67),
    .Y(_08851_));
 AO21x1_ASAP7_75t_R _16975_ (.A1(_08850_),
    .A2(net6674),
    .B(_08851_),
    .Y(_00356_));
 XOR2x2_ASAP7_75t_R _16976_ (.A(_08758_),
    .B(_00906_),
    .Y(_08852_));
 AND2x2_ASAP7_75t_R _16977_ (.A(net6684),
    .B(net68),
    .Y(_08853_));
 AO21x1_ASAP7_75t_R _16978_ (.A1(_08852_),
    .A2(_08030_),
    .B(_08853_),
    .Y(_00357_));
 XOR2x2_ASAP7_75t_R _16979_ (.A(_08760_),
    .B(_00907_),
    .Y(_08854_));
 AND2x2_ASAP7_75t_R _16981_ (.A(net6684),
    .B(net69),
    .Y(_08856_));
 AO21x1_ASAP7_75t_R _16982_ (.A1(_08854_),
    .A2(_08030_),
    .B(_08856_),
    .Y(_00358_));
 XOR2x2_ASAP7_75t_R _16983_ (.A(_08762_),
    .B(_00908_),
    .Y(_08857_));
 AND2x2_ASAP7_75t_R _16985_ (.A(net6681),
    .B(net70),
    .Y(_08859_));
 AO21x1_ASAP7_75t_R _16986_ (.A1(_08857_),
    .A2(net6677),
    .B(_08859_),
    .Y(_00359_));
 XOR2x2_ASAP7_75t_R _16987_ (.A(_08765_),
    .B(net6489),
    .Y(_08860_));
 AND2x2_ASAP7_75t_R _16988_ (.A(net6689),
    .B(net71),
    .Y(_08861_));
 AO21x1_ASAP7_75t_R _16989_ (.A1(_08860_),
    .A2(net6678),
    .B(_08861_),
    .Y(_00360_));
 XOR2x2_ASAP7_75t_R _16990_ (.A(_08769_),
    .B(net6488),
    .Y(_08862_));
 AND2x2_ASAP7_75t_R _16991_ (.A(net6688),
    .B(net72),
    .Y(_08863_));
 AO21x1_ASAP7_75t_R _16992_ (.A1(_08862_),
    .A2(net6678),
    .B(_08863_),
    .Y(_00361_));
 AND2x2_ASAP7_75t_R _16993_ (.A(net6689),
    .B(net74),
    .Y(_08864_));
 AO21x1_ASAP7_75t_R _16994_ (.A1(_08054_),
    .A2(net6678),
    .B(_08864_),
    .Y(_00362_));
 XOR2x2_ASAP7_75t_R _16995_ (.A(_08776_),
    .B(_00912_),
    .Y(_08865_));
 AND2x2_ASAP7_75t_R _16996_ (.A(net6688),
    .B(net75),
    .Y(_08866_));
 AO21x1_ASAP7_75t_R _16997_ (.A1(_08865_),
    .A2(net6678),
    .B(_08866_),
    .Y(_00363_));
 XOR2x2_ASAP7_75t_R _16998_ (.A(_08779_),
    .B(net6486),
    .Y(_08867_));
 AND2x2_ASAP7_75t_R _16999_ (.A(net6682),
    .B(net76),
    .Y(_08868_));
 AO21x1_ASAP7_75t_R _17000_ (.A1(_08867_),
    .A2(net6677),
    .B(_08868_),
    .Y(_00365_));
 XOR2x2_ASAP7_75t_R _17001_ (.A(_08781_),
    .B(_00915_),
    .Y(_08869_));
 AND2x2_ASAP7_75t_R _17002_ (.A(net6689),
    .B(net77),
    .Y(_08870_));
 AO21x1_ASAP7_75t_R _17003_ (.A1(_08869_),
    .A2(net6678),
    .B(_08870_),
    .Y(_00366_));
 XOR2x2_ASAP7_75t_R _17004_ (.A(_08783_),
    .B(_00916_),
    .Y(_08871_));
 AND2x2_ASAP7_75t_R _17005_ (.A(net6682),
    .B(net78),
    .Y(_08872_));
 AO21x1_ASAP7_75t_R _17006_ (.A1(_08871_),
    .A2(net6677),
    .B(_08872_),
    .Y(_00367_));
 XOR2x2_ASAP7_75t_R _17007_ (.A(_08785_),
    .B(net6485),
    .Y(_08873_));
 AND2x2_ASAP7_75t_R _17008_ (.A(net6689),
    .B(net79),
    .Y(_08874_));
 AO21x1_ASAP7_75t_R _17009_ (.A1(_08873_),
    .A2(net6678),
    .B(_08874_),
    .Y(_00368_));
 INVx1_ASAP7_75t_R _17010_ (.A(net6484),
    .Y(_08875_));
 OA21x2_ASAP7_75t_R _17011_ (.A1(net6383),
    .A2(_08875_),
    .B(net6677),
    .Y(_08876_));
 NAND2x1_ASAP7_75t_R _17012_ (.A(_08875_),
    .B(net6383),
    .Y(_08877_));
 AO22x1_ASAP7_75t_R _17013_ (.A1(net6689),
    .A2(net80),
    .B1(_08876_),
    .B2(_08877_),
    .Y(_00369_));
 NAND2x1_ASAP7_75t_R _17014_ (.A(_00414_),
    .B(_08791_),
    .Y(_08878_));
 NAND2x1_ASAP7_75t_R _17015_ (.A(_08789_),
    .B(net6390),
    .Y(_08879_));
 AO21x1_ASAP7_75t_R _17016_ (.A1(_08878_),
    .A2(_08879_),
    .B(net6483),
    .Y(_08880_));
 INVx1_ASAP7_75t_R _17017_ (.A(_00919_),
    .Y(_08881_));
 AO21x1_ASAP7_75t_R _17018_ (.A1(_08792_),
    .A2(_08794_),
    .B(net6467),
    .Y(_08882_));
 AND3x1_ASAP7_75t_R _17019_ (.A(_08880_),
    .B(_08882_),
    .C(net6678),
    .Y(_08883_));
 AO21x1_ASAP7_75t_R _17020_ (.A1(net6688),
    .A2(net81),
    .B(_08883_),
    .Y(_00370_));
 AOI21x1_ASAP7_75t_R _17021_ (.A1(net6482),
    .A2(_08798_),
    .B(net6688),
    .Y(_08884_));
 XOR2x2_ASAP7_75t_R _17022_ (.A(_00856_),
    .B(_00888_),
    .Y(_08885_));
 XNOR2x2_ASAP7_75t_R _17023_ (.A(_00832_),
    .B(_08885_),
    .Y(_08886_));
 NAND2x1_ASAP7_75t_R _17024_ (.A(_00415_),
    .B(_08886_),
    .Y(_08887_));
 INVx1_ASAP7_75t_R _17025_ (.A(_00415_),
    .Y(_08888_));
 XOR2x2_ASAP7_75t_R _17026_ (.A(_08885_),
    .B(_00832_),
    .Y(_08889_));
 NAND2x1_ASAP7_75t_R _17027_ (.A(_08888_),
    .B(_08889_),
    .Y(_08890_));
 AO21x1_ASAP7_75t_R _17028_ (.A1(_08887_),
    .A2(_08890_),
    .B(net6482),
    .Y(_08891_));
 AO22x1_ASAP7_75t_R _17029_ (.A1(net6688),
    .A2(net82),
    .B1(_08884_),
    .B2(_08891_),
    .Y(_00371_));
 INVx1_ASAP7_75t_R _17030_ (.A(net6481),
    .Y(_08892_));
 XOR2x2_ASAP7_75t_R _17031_ (.A(_08806_),
    .B(_08892_),
    .Y(_08893_));
 AND2x2_ASAP7_75t_R _17032_ (.A(net6688),
    .B(net83),
    .Y(_08894_));
 AO21x1_ASAP7_75t_R _17033_ (.A1(_08893_),
    .A2(net6678),
    .B(_08894_),
    .Y(_00372_));
 INVx1_ASAP7_75t_R _17034_ (.A(_00922_),
    .Y(_08895_));
 XOR2x2_ASAP7_75t_R _17035_ (.A(_08808_),
    .B(_08895_),
    .Y(_08896_));
 AND2x2_ASAP7_75t_R _17036_ (.A(net6688),
    .B(net85),
    .Y(_08897_));
 AO21x1_ASAP7_75t_R _17037_ (.A1(_08896_),
    .A2(net6677),
    .B(_08897_),
    .Y(_00373_));
 INVx1_ASAP7_75t_R _17038_ (.A(_00923_),
    .Y(_08898_));
 XOR2x2_ASAP7_75t_R _17039_ (.A(_08810_),
    .B(_08898_),
    .Y(_08899_));
 AND2x2_ASAP7_75t_R _17040_ (.A(net6688),
    .B(net86),
    .Y(_08900_));
 AO21x1_ASAP7_75t_R _17041_ (.A1(_08899_),
    .A2(net6677),
    .B(_08900_),
    .Y(_00374_));
 XOR2x2_ASAP7_75t_R _17042_ (.A(_08812_),
    .B(_00925_),
    .Y(_08901_));
 NOR2x1_ASAP7_75t_R _17043_ (.A(net6688),
    .B(_08901_),
    .Y(_08902_));
 AO21x1_ASAP7_75t_R _17044_ (.A1(net6688),
    .A2(net87),
    .B(_08902_),
    .Y(_00376_));
 XOR2x2_ASAP7_75t_R _17046_ (.A(_08814_),
    .B(_00926_),
    .Y(_08904_));
 NOR2x1_ASAP7_75t_R _17047_ (.A(net6686),
    .B(_08904_),
    .Y(_08905_));
 AO21x1_ASAP7_75t_R _17048_ (.A1(net6686),
    .A2(net88),
    .B(_08905_),
    .Y(_00377_));
 INVx1_ASAP7_75t_R _17050_ (.A(net1),
    .Y(_08907_));
 INVx1_ASAP7_75t_R _17051_ (.A(_00934_),
    .Y(_08908_));
 XOR2x2_ASAP7_75t_R _17052_ (.A(_08817_),
    .B(_08908_),
    .Y(_08909_));
 NOR2x1_ASAP7_75t_R _17053_ (.A(net129),
    .B(_08909_),
    .Y(_08910_));
 AO21x1_ASAP7_75t_R _17054_ (.A1(net6685),
    .A2(_08907_),
    .B(_08910_),
    .Y(_08911_));
 INVx1_ASAP7_75t_R _17056_ (.A(net40),
    .Y(_08912_));
 INVx1_ASAP7_75t_R _17057_ (.A(_00945_),
    .Y(_08913_));
 XOR2x2_ASAP7_75t_R _17058_ (.A(_08820_),
    .B(_08913_),
    .Y(_08914_));
 NOR2x1p5_ASAP7_75t_R _17059_ (.A(net129),
    .B(_08914_),
    .Y(_08915_));
 AOI21x1_ASAP7_75t_R _17060_ (.A1(net129),
    .A2(_08912_),
    .B(_08915_),
    .Y(_08916_));
 INVx1_ASAP7_75t_R _17061_ (.A(net6323),
    .Y(_01025_));
 OR2x2_ASAP7_75t_R _17062_ (.A(net51),
    .B(_08030_),
    .Y(_08917_));
 XOR2x2_ASAP7_75t_R _17063_ (.A(_00924_),
    .B(_00956_),
    .Y(_08918_));
 XOR2x2_ASAP7_75t_R _17064_ (.A(_08918_),
    .B(_00423_),
    .Y(_08919_));
 XOR2x2_ASAP7_75t_R _17065_ (.A(_08919_),
    .B(_08727_),
    .Y(_08920_));
 NAND2x1_ASAP7_75t_R _17066_ (.A(net6674),
    .B(_08920_),
    .Y(_08921_));
 NAND2x1_ASAP7_75t_R _17067_ (.A(_08917_),
    .B(_08921_),
    .Y(_08922_));
 INVx1_ASAP7_75t_R _17068_ (.A(_08922_),
    .Y(_08923_));
 INVx1_ASAP7_75t_R _17070_ (.A(_00959_),
    .Y(_08924_));
 NOR2x1_ASAP7_75t_R _17071_ (.A(_08924_),
    .B(_08826_),
    .Y(_08925_));
 AND2x2_ASAP7_75t_R _17072_ (.A(_08826_),
    .B(_08924_),
    .Y(_08926_));
 OAI21x1_ASAP7_75t_R _17073_ (.A1(_08925_),
    .A2(_08926_),
    .B(net6675),
    .Y(_08927_));
 OAI21x1_ASAP7_75t_R _17074_ (.A1(net6675),
    .A2(net62),
    .B(_08927_),
    .Y(_08928_));
 INVx2_ASAP7_75t_R _17075_ (.A(_08928_),
    .Y(_08929_));
 XOR2x2_ASAP7_75t_R _17078_ (.A(_08829_),
    .B(_00960_),
    .Y(_08931_));
 NOR2x1_ASAP7_75t_R _17079_ (.A(net73),
    .B(_08030_),
    .Y(_08932_));
 AOI21x1_ASAP7_75t_R _17080_ (.A1(_08030_),
    .A2(_08931_),
    .B(_08932_),
    .Y(_08933_));
 XOR2x2_ASAP7_75t_R _17082_ (.A(_08832_),
    .B(_00961_),
    .Y(_08934_));
 NOR2x1_ASAP7_75t_R _17083_ (.A(net84),
    .B(_08030_),
    .Y(_08935_));
 AOI21x1_ASAP7_75t_R _17084_ (.A1(_08030_),
    .A2(_08934_),
    .B(_08935_),
    .Y(_08936_));
 XOR2x2_ASAP7_75t_R _17087_ (.A(_08834_),
    .B(_00962_),
    .Y(_08938_));
 NAND2x1_ASAP7_75t_R _17088_ (.A(_08030_),
    .B(_08938_),
    .Y(_08939_));
 OA21x2_ASAP7_75t_R _17089_ (.A1(_08030_),
    .A2(net95),
    .B(_08939_),
    .Y(_08940_));
 XOR2x2_ASAP7_75t_R _17092_ (.A(_08836_),
    .B(_00963_),
    .Y(_08942_));
 NAND2x1_ASAP7_75t_R _17093_ (.A(net6675),
    .B(_08942_),
    .Y(_08943_));
 OA21x2_ASAP7_75t_R _17094_ (.A1(net6675),
    .A2(net106),
    .B(_08943_),
    .Y(_08944_));
 INVx1_ASAP7_75t_R _17097_ (.A(net117),
    .Y(_08946_));
 INVx1_ASAP7_75t_R _17098_ (.A(_00964_),
    .Y(_08947_));
 XOR2x2_ASAP7_75t_R _17099_ (.A(_08839_),
    .B(_08947_),
    .Y(_08948_));
 NOR2x1_ASAP7_75t_R _17100_ (.A(net6690),
    .B(_08948_),
    .Y(_08949_));
 AOI21x1_ASAP7_75t_R _17101_ (.A1(net6690),
    .A2(_08946_),
    .B(_08949_),
    .Y(_08950_));
 INVx1_ASAP7_75t_R _17103_ (.A(net6311),
    .Y(_01000_));
 XOR2x2_ASAP7_75t_R _17104_ (.A(_08841_),
    .B(_00430_),
    .Y(_08951_));
 XOR2x2_ASAP7_75t_R _17105_ (.A(_00486_),
    .B(_00869_),
    .Y(_08952_));
 XOR2x2_ASAP7_75t_R _17106_ (.A(_08951_),
    .B(_08952_),
    .Y(_08953_));
 NAND2x1_ASAP7_75t_R _17107_ (.A(_08030_),
    .B(_08953_),
    .Y(_08954_));
 OAI21x1_ASAP7_75t_R _17108_ (.A1(_08030_),
    .A2(net128),
    .B(_08954_),
    .Y(_08955_));
 OR2x2_ASAP7_75t_R _17110_ (.A(net12),
    .B(_08030_),
    .Y(_08956_));
 XOR2x2_ASAP7_75t_R _17111_ (.A(_00903_),
    .B(_00935_),
    .Y(_08957_));
 XOR2x2_ASAP7_75t_R _17112_ (.A(_08957_),
    .B(_00431_),
    .Y(_08958_));
 XOR2x2_ASAP7_75t_R _17113_ (.A(_08958_),
    .B(_08749_),
    .Y(_08959_));
 NAND2x1_ASAP7_75t_R _17114_ (.A(_08030_),
    .B(_08959_),
    .Y(_08960_));
 NAND2x2_ASAP7_75t_R _17115_ (.A(_08956_),
    .B(_08960_),
    .Y(_08961_));
 INVx2_ASAP7_75t_R _17116_ (.A(_08961_),
    .Y(_08962_));
 INVx1_ASAP7_75t_R _17118_ (.A(_00936_),
    .Y(_08963_));
 NOR2x1_ASAP7_75t_R _17119_ (.A(_08963_),
    .B(_08848_),
    .Y(_08964_));
 AND2x2_ASAP7_75t_R _17120_ (.A(_08848_),
    .B(_08963_),
    .Y(_08965_));
 OAI21x1_ASAP7_75t_R _17121_ (.A1(_08964_),
    .A2(_08965_),
    .B(net6674),
    .Y(_08966_));
 OAI21x1_ASAP7_75t_R _17122_ (.A1(net6674),
    .A2(net23),
    .B(_08966_),
    .Y(_08967_));
 INVx2_ASAP7_75t_R _17123_ (.A(_08967_),
    .Y(_08968_));
 XOR2x2_ASAP7_75t_R _17126_ (.A(_08850_),
    .B(_00937_),
    .Y(_08970_));
 NOR2x1_ASAP7_75t_R _17127_ (.A(net32),
    .B(net6675),
    .Y(_08971_));
 AOI21x1_ASAP7_75t_R _17128_ (.A1(_08030_),
    .A2(_08970_),
    .B(_08971_),
    .Y(_08972_));
 XOR2x2_ASAP7_75t_R _17131_ (.A(_08852_),
    .B(_00938_),
    .Y(_08974_));
 NOR2x1_ASAP7_75t_R _17132_ (.A(net33),
    .B(net6675),
    .Y(_08975_));
 AOI21x1_ASAP7_75t_R _17133_ (.A1(_08030_),
    .A2(_08974_),
    .B(_08975_),
    .Y(_08976_));
 XOR2x2_ASAP7_75t_R _17136_ (.A(_08854_),
    .B(_00939_),
    .Y(_08978_));
 NAND2x1_ASAP7_75t_R _17137_ (.A(net6675),
    .B(_08978_),
    .Y(_08979_));
 OA21x2_ASAP7_75t_R _17138_ (.A1(net6675),
    .A2(net34),
    .B(_08979_),
    .Y(_08980_));
 XOR2x2_ASAP7_75t_R _17141_ (.A(_08857_),
    .B(_00940_),
    .Y(_08982_));
 NAND2x1_ASAP7_75t_R _17142_ (.A(net6675),
    .B(_08982_),
    .Y(_08983_));
 OA21x2_ASAP7_75t_R _17143_ (.A1(net6676),
    .A2(net35),
    .B(_08983_),
    .Y(_08984_));
 XOR2x2_ASAP7_75t_R _17145_ (.A(_00918_),
    .B(_00950_),
    .Y(_08985_));
 INVx1_ASAP7_75t_R _17146_ (.A(_08985_),
    .Y(_08986_));
 INVx1_ASAP7_75t_R _17147_ (.A(_00886_),
    .Y(_08987_));
 XOR2x2_ASAP7_75t_R _17148_ (.A(_08696_),
    .B(_08987_),
    .Y(_08988_));
 NAND2x1_ASAP7_75t_R _17149_ (.A(_08986_),
    .B(_08988_),
    .Y(_08989_));
 AOI21x1_ASAP7_75t_R _17150_ (.A1(_08985_),
    .A2(net6383),
    .B(net6687),
    .Y(_08990_));
 AND2x2_ASAP7_75t_R _17151_ (.A(net6690),
    .B(net45),
    .Y(_08991_));
 AOI21x1_ASAP7_75t_R _17152_ (.A1(_08989_),
    .A2(_08990_),
    .B(_08991_),
    .Y(_08992_));
 XOR2x2_ASAP7_75t_R _17154_ (.A(_00919_),
    .B(_00951_),
    .Y(_08993_));
 AOI21x1_ASAP7_75t_R _17155_ (.A1(_08794_),
    .A2(_08792_),
    .B(_08993_),
    .Y(_08994_));
 AO31x2_ASAP7_75t_R _17156_ (.A1(_08993_),
    .A2(_08794_),
    .A3(_08792_),
    .B(net6690),
    .Y(_08995_));
 NAND2x1_ASAP7_75t_R _17157_ (.A(net6690),
    .B(net46),
    .Y(_08996_));
 OAI21x1_ASAP7_75t_R _17158_ (.A1(_08995_),
    .A2(_08994_),
    .B(_08996_),
    .Y(_08997_));
 INVx2_ASAP7_75t_R _17159_ (.A(net6300),
    .Y(_01047_));
 NOR2x1_ASAP7_75t_R _17160_ (.A(net47),
    .B(net6676),
    .Y(_08998_));
 INVx1_ASAP7_75t_R _17161_ (.A(_08998_),
    .Y(_08999_));
 NAND2x1_ASAP7_75t_R _17162_ (.A(_00415_),
    .B(_08889_),
    .Y(_09000_));
 NAND2x1_ASAP7_75t_R _17163_ (.A(_08888_),
    .B(_08886_),
    .Y(_09001_));
 XOR2x2_ASAP7_75t_R _17164_ (.A(_00920_),
    .B(_00952_),
    .Y(_09002_));
 AOI21x1_ASAP7_75t_R _17165_ (.A1(_09000_),
    .A2(_09001_),
    .B(_09002_),
    .Y(_09003_));
 INVx1_ASAP7_75t_R _17166_ (.A(_09002_),
    .Y(_09004_));
 AOI21x1_ASAP7_75t_R _17167_ (.A1(_08890_),
    .A2(_08887_),
    .B(_09004_),
    .Y(_09005_));
 OAI21x1_ASAP7_75t_R _17168_ (.A1(_09003_),
    .A2(_09005_),
    .B(net6679),
    .Y(_09006_));
 NAND2x1_ASAP7_75t_R _17169_ (.A(_08999_),
    .B(_09006_),
    .Y(_09007_));
 NOR2x1_ASAP7_75t_R _17171_ (.A(_08803_),
    .B(_08801_),
    .Y(_09008_));
 NOR2x1_ASAP7_75t_R _17172_ (.A(_00416_),
    .B(_08804_),
    .Y(_09009_));
 XNOR2x2_ASAP7_75t_R _17173_ (.A(_00921_),
    .B(_00953_),
    .Y(_09010_));
 INVx1_ASAP7_75t_R _17174_ (.A(_09010_),
    .Y(_09011_));
 OAI21x1_ASAP7_75t_R _17175_ (.A1(_09008_),
    .A2(_09009_),
    .B(_09011_),
    .Y(_09012_));
 OAI21x1_ASAP7_75t_R _17176_ (.A1(_08802_),
    .A2(_08805_),
    .B(_09010_),
    .Y(_09013_));
 NAND2x1_ASAP7_75t_R _17177_ (.A(_09012_),
    .B(_09013_),
    .Y(_09014_));
 NOR2x1_ASAP7_75t_R _17178_ (.A(net48),
    .B(net6676),
    .Y(_09015_));
 AOI21x1_ASAP7_75t_R _17179_ (.A1(net6676),
    .A2(_09014_),
    .B(_09015_),
    .Y(_09016_));
 XNOR2x2_ASAP7_75t_R _17182_ (.A(_00922_),
    .B(_00954_),
    .Y(_09018_));
 XOR2x2_ASAP7_75t_R _17183_ (.A(_08808_),
    .B(_09018_),
    .Y(_09019_));
 NOR2x1_ASAP7_75t_R _17184_ (.A(net49),
    .B(net6677),
    .Y(_09020_));
 AOI21x1_ASAP7_75t_R _17185_ (.A1(net6676),
    .A2(_09019_),
    .B(_09020_),
    .Y(_09021_));
 XNOR2x2_ASAP7_75t_R _17188_ (.A(_00923_),
    .B(_00955_),
    .Y(_09023_));
 XOR2x2_ASAP7_75t_R _17189_ (.A(_08810_),
    .B(_09023_),
    .Y(_09024_));
 NAND2x1_ASAP7_75t_R _17190_ (.A(net6675),
    .B(_09024_),
    .Y(_09025_));
 OAI21x1_ASAP7_75t_R _17191_ (.A1(net6675),
    .A2(net50),
    .B(_09025_),
    .Y(_09026_));
 INVx1_ASAP7_75t_R _17192_ (.A(_09026_),
    .Y(_09027_));
 XNOR2x2_ASAP7_75t_R _17194_ (.A(_00957_),
    .B(_08901_),
    .Y(_09028_));
 NOR2x1_ASAP7_75t_R _17195_ (.A(net52),
    .B(net6676),
    .Y(_09029_));
 AOI21x1_ASAP7_75t_R _17196_ (.A1(net6676),
    .A2(_09028_),
    .B(_09029_),
    .Y(_09030_));
 XNOR2x2_ASAP7_75t_R _17199_ (.A(_00958_),
    .B(_08904_),
    .Y(_09032_));
 NAND2x1_ASAP7_75t_R _17200_ (.A(net6675),
    .B(_09032_),
    .Y(_09033_));
 OA21x2_ASAP7_75t_R _17201_ (.A1(net6675),
    .A2(net53),
    .B(_09033_),
    .Y(_09034_));
 INVx6_ASAP7_75t_R _17203_ (.A(_08955_),
    .Y(_00995_));
 NOR2x1_ASAP7_75t_R _17205_ (.A(net5260),
    .B(net6308),
    .Y(_09035_));
 INVx1_ASAP7_75t_R _17206_ (.A(_09035_),
    .Y(_09036_));
 INVx1_ASAP7_75t_R _17209_ (.A(_00997_),
    .Y(_09039_));
 AO21x1_ASAP7_75t_R _17210_ (.A1(net6367),
    .A2(net6465),
    .B(net5241),
    .Y(_09040_));
 AO21x1_ASAP7_75t_R _17212_ (.A1(_09036_),
    .A2(_09040_),
    .B(net5948),
    .Y(_09042_));
 INVx2_ASAP7_75t_R _17213_ (.A(_08972_),
    .Y(_09043_));
 INVx1_ASAP7_75t_R _17215_ (.A(_01004_),
    .Y(_09045_));
 NOR2x1_ASAP7_75t_R _17216_ (.A(_09045_),
    .B(net6308),
    .Y(_09046_));
 INVx1_ASAP7_75t_R _17217_ (.A(_01006_),
    .Y(_09047_));
 AO21x1_ASAP7_75t_R _17218_ (.A1(net6367),
    .A2(net6465),
    .B(_09047_),
    .Y(_09048_));
 INVx1_ASAP7_75t_R _17219_ (.A(_09048_),
    .Y(_09049_));
 OAI21x1_ASAP7_75t_R _17221_ (.A1(_09046_),
    .A2(_09049_),
    .B(net5948),
    .Y(_09051_));
 AND3x1_ASAP7_75t_R _17222_ (.A(_09042_),
    .B(net5927),
    .C(_09051_),
    .Y(_09052_));
 NAND2x1_ASAP7_75t_R _17223_ (.A(net6309),
    .B(net5952),
    .Y(_09053_));
 NAND2x1_ASAP7_75t_R _17224_ (.A(_08962_),
    .B(net6310),
    .Y(_09054_));
 AO21x1_ASAP7_75t_R _17227_ (.A1(_09053_),
    .A2(net5556),
    .B(net6305),
    .Y(_09057_));
 AOI21x1_ASAP7_75t_R _17230_ (.A1(net5951),
    .A2(net6311),
    .B(net5946),
    .Y(_09060_));
 NAND2x1_ASAP7_75t_R _17231_ (.A(_09060_),
    .B(_09053_),
    .Y(_09061_));
 AO31x2_ASAP7_75t_R _17232_ (.A1(_09057_),
    .A2(net6304),
    .A3(_09061_),
    .B(net5943),
    .Y(_09062_));
 NOR2x1_ASAP7_75t_R _17233_ (.A(net5317),
    .B(net6308),
    .Y(_09063_));
 INVx1_ASAP7_75t_R _17234_ (.A(_01001_),
    .Y(_09064_));
 AO21x1_ASAP7_75t_R _17235_ (.A1(net6367),
    .A2(net6465),
    .B(_09064_),
    .Y(_09065_));
 INVx1_ASAP7_75t_R _17236_ (.A(_09065_),
    .Y(_09066_));
 OAI21x1_ASAP7_75t_R _17238_ (.A1(_09063_),
    .A2(_09066_),
    .B(net5945),
    .Y(_09068_));
 OAI21x1_ASAP7_75t_R _17241_ (.A1(net5950),
    .A2(net6310),
    .B(net6307),
    .Y(_09071_));
 AND2x2_ASAP7_75t_R _17242_ (.A(_09071_),
    .B(net5926),
    .Y(_09072_));
 INVx1_ASAP7_75t_R _17243_ (.A(_08980_),
    .Y(_09073_));
 AOI21x1_ASAP7_75t_R _17245_ (.A1(_09068_),
    .A2(_09072_),
    .B(net5554),
    .Y(_09075_));
 INVx1_ASAP7_75t_R _17246_ (.A(net5260),
    .Y(_09076_));
 NOR2x2_ASAP7_75t_R _17247_ (.A(_09076_),
    .B(net6308),
    .Y(_09077_));
 NOR2x1p5_ASAP7_75t_R _17248_ (.A(net6307),
    .B(_09077_),
    .Y(_09078_));
 INVx1_ASAP7_75t_R _17249_ (.A(_09078_),
    .Y(_09079_));
 INVx1_ASAP7_75t_R _17250_ (.A(net5320),
    .Y(_09080_));
 NOR2x1_ASAP7_75t_R _17251_ (.A(_09080_),
    .B(net5950),
    .Y(_09081_));
 NAND2x1_ASAP7_75t_R _17252_ (.A(net5950),
    .B(net5952),
    .Y(_09082_));
 OA21x2_ASAP7_75t_R _17253_ (.A1(net5950),
    .A2(net5319),
    .B(net6307),
    .Y(_09083_));
 AOI21x1_ASAP7_75t_R _17255_ (.A1(_09082_),
    .A2(_09083_),
    .B(net5926),
    .Y(_09085_));
 OAI21x1_ASAP7_75t_R _17256_ (.A1(_09079_),
    .A2(_09081_),
    .B(_09085_),
    .Y(_09086_));
 AOI21x1_ASAP7_75t_R _17257_ (.A1(_09075_),
    .A2(_09086_),
    .B(net5942),
    .Y(_09087_));
 OAI21x1_ASAP7_75t_R _17258_ (.A1(_09052_),
    .A2(_09062_),
    .B(_09087_),
    .Y(_09088_));
 NAND2x1_ASAP7_75t_R _17259_ (.A(_09064_),
    .B(_08962_),
    .Y(_09089_));
 AND2x2_ASAP7_75t_R _17260_ (.A(_09089_),
    .B(net5948),
    .Y(_09090_));
 INVx1_ASAP7_75t_R _17261_ (.A(_01005_),
    .Y(_09091_));
 AO21x1_ASAP7_75t_R _17262_ (.A1(net6367),
    .A2(net6465),
    .B(_09091_),
    .Y(_09092_));
 NOR2x1_ASAP7_75t_R _17264_ (.A(_01007_),
    .B(net6308),
    .Y(_09094_));
 INVx1_ASAP7_75t_R _17265_ (.A(_09094_),
    .Y(_09095_));
 NOR2x1_ASAP7_75t_R _17266_ (.A(net5948),
    .B(_09095_),
    .Y(_09096_));
 AO21x1_ASAP7_75t_R _17267_ (.A1(_09090_),
    .A2(net5240),
    .B(_09096_),
    .Y(_09097_));
 NOR2x1_ASAP7_75t_R _17268_ (.A(net6304),
    .B(_09097_),
    .Y(_09098_));
 NOR2x1_ASAP7_75t_R _17270_ (.A(_09064_),
    .B(net6308),
    .Y(_09100_));
 NOR2x1_ASAP7_75t_R _17272_ (.A(net6305),
    .B(_09095_),
    .Y(_09102_));
 AOI21x1_ASAP7_75t_R _17273_ (.A1(net6305),
    .A2(net4975),
    .B(_09102_),
    .Y(_09103_));
 NOR2x2_ASAP7_75t_R _17275_ (.A(_09045_),
    .B(net5949),
    .Y(_09105_));
 AOI21x1_ASAP7_75t_R _17277_ (.A1(net6305),
    .A2(_09105_),
    .B(_09043_),
    .Y(_09107_));
 AO21x1_ASAP7_75t_R _17279_ (.A1(_09103_),
    .A2(_09107_),
    .B(net5943),
    .Y(_09109_));
 AO21x1_ASAP7_75t_R _17280_ (.A1(_09095_),
    .A2(_09048_),
    .B(net5948),
    .Y(_09110_));
 AO21x1_ASAP7_75t_R _17281_ (.A1(net5951),
    .A2(net5317),
    .B(net6306),
    .Y(_09111_));
 AND2x2_ASAP7_75t_R _17282_ (.A(_09111_),
    .B(net6304),
    .Y(_09112_));
 AOI21x1_ASAP7_75t_R _17283_ (.A1(_09110_),
    .A2(_09112_),
    .B(net5554),
    .Y(_09113_));
 NAND2x1_ASAP7_75t_R _17284_ (.A(net6309),
    .B(_08962_),
    .Y(_09114_));
 AO21x2_ASAP7_75t_R _17285_ (.A1(net6367),
    .A2(net6465),
    .B(_09076_),
    .Y(_09115_));
 AND3x1_ASAP7_75t_R _17286_ (.A(net5553),
    .B(net6305),
    .C(net4787),
    .Y(_09116_));
 AO21x1_ASAP7_75t_R _17287_ (.A1(net6311),
    .A2(_08962_),
    .B(net6307),
    .Y(_09117_));
 NOR2x1_ASAP7_75t_R _17288_ (.A(_09105_),
    .B(_09117_),
    .Y(_09118_));
 OAI21x1_ASAP7_75t_R _17290_ (.A1(_09116_),
    .A2(_09118_),
    .B(net5928),
    .Y(_09120_));
 INVx1_ASAP7_75t_R _17291_ (.A(_08984_),
    .Y(_09121_));
 AOI21x1_ASAP7_75t_R _17292_ (.A1(_09113_),
    .A2(_09120_),
    .B(_09121_),
    .Y(_09122_));
 OAI21x1_ASAP7_75t_R _17293_ (.A1(_09098_),
    .A2(_09109_),
    .B(_09122_),
    .Y(_09123_));
 INVx1_ASAP7_75t_R _17294_ (.A(_08976_),
    .Y(_09124_));
 AOI21x1_ASAP7_75t_R _17296_ (.A1(_09088_),
    .A2(_09123_),
    .B(net5924),
    .Y(_09126_));
 AO21x1_ASAP7_75t_R _17297_ (.A1(net6367),
    .A2(net6465),
    .B(net5260),
    .Y(_09127_));
 NAND2x1_ASAP7_75t_R _17298_ (.A(net6306),
    .B(net5025),
    .Y(_09128_));
 NAND2x1_ASAP7_75t_R _17299_ (.A(_01014_),
    .B(net5948),
    .Y(_09129_));
 AO21x1_ASAP7_75t_R _17300_ (.A1(_09128_),
    .A2(_09129_),
    .B(net5929),
    .Y(_09130_));
 NOR2x1_ASAP7_75t_R _17301_ (.A(_08962_),
    .B(net6310),
    .Y(_09131_));
 INVx1_ASAP7_75t_R _17302_ (.A(_09131_),
    .Y(_09132_));
 INVx1_ASAP7_75t_R _17303_ (.A(_09100_),
    .Y(_09133_));
 AO21x1_ASAP7_75t_R _17304_ (.A1(_09132_),
    .A2(_09133_),
    .B(net5948),
    .Y(_09134_));
 NAND2x1_ASAP7_75t_R _17305_ (.A(_09047_),
    .B(net5951),
    .Y(_09135_));
 NOR2x1_ASAP7_75t_R _17306_ (.A(net6307),
    .B(_09131_),
    .Y(_09136_));
 AOI21x1_ASAP7_75t_R _17307_ (.A1(_09135_),
    .A2(_09136_),
    .B(net6304),
    .Y(_09137_));
 NAND2x1_ASAP7_75t_R _17308_ (.A(_09134_),
    .B(_09137_),
    .Y(_09138_));
 AOI21x1_ASAP7_75t_R _17309_ (.A1(_09130_),
    .A2(_09138_),
    .B(net5943),
    .Y(_09139_));
 NOR2x1_ASAP7_75t_R _17310_ (.A(_00997_),
    .B(net6308),
    .Y(_09140_));
 INVx1_ASAP7_75t_R _17311_ (.A(_09140_),
    .Y(_09141_));
 AOI21x1_ASAP7_75t_R _17312_ (.A1(_09141_),
    .A2(_09136_),
    .B(net6304),
    .Y(_09142_));
 NOR2x1_ASAP7_75t_R _17313_ (.A(net5570),
    .B(net6308),
    .Y(_09143_));
 AOI211x1_ASAP7_75t_R _17314_ (.A1(net6305),
    .A2(net5549),
    .B(_09078_),
    .C(_09043_),
    .Y(_09144_));
 AO21x1_ASAP7_75t_R _17315_ (.A1(net6367),
    .A2(net6465),
    .B(net5318),
    .Y(_09145_));
 NOR2x1_ASAP7_75t_R _17316_ (.A(net5948),
    .B(_09145_),
    .Y(_09146_));
 NOR2x1_ASAP7_75t_R _17317_ (.A(_09146_),
    .B(net5554),
    .Y(_09147_));
 OAI21x1_ASAP7_75t_R _17318_ (.A1(_09142_),
    .A2(_09144_),
    .B(_09147_),
    .Y(_09148_));
 NAND2x1_ASAP7_75t_R _17319_ (.A(net5942),
    .B(_09148_),
    .Y(_09149_));
 OAI21x1_ASAP7_75t_R _17320_ (.A1(_09139_),
    .A2(_09149_),
    .B(net5924),
    .Y(_09150_));
 NAND2x1_ASAP7_75t_R _17321_ (.A(net6308),
    .B(net6309),
    .Y(_09151_));
 AO21x1_ASAP7_75t_R _17322_ (.A1(_09095_),
    .A2(net5923),
    .B(net5945),
    .Y(_09152_));
 AO21x1_ASAP7_75t_R _17323_ (.A1(net6308),
    .A2(_09064_),
    .B(net5945),
    .Y(_09153_));
 INVx1_ASAP7_75t_R _17324_ (.A(_09114_),
    .Y(_09154_));
 OA21x2_ASAP7_75t_R _17325_ (.A1(_09153_),
    .A2(_09154_),
    .B(net6304),
    .Y(_09155_));
 NAND2x1_ASAP7_75t_R _17326_ (.A(net5320),
    .B(net5949),
    .Y(_09156_));
 NAND2x1_ASAP7_75t_R _17327_ (.A(net5236),
    .B(_09136_),
    .Y(_09157_));
 AO22x1_ASAP7_75t_R _17328_ (.A1(_09152_),
    .A2(_09142_),
    .B1(_09155_),
    .B2(_09157_),
    .Y(_09158_));
 NOR2x1_ASAP7_75t_R _17329_ (.A(_09047_),
    .B(net6308),
    .Y(_09159_));
 OAI21x1_ASAP7_75t_R _17331_ (.A1(net4973),
    .A2(net5238),
    .B(net6305),
    .Y(_09161_));
 AO21x1_ASAP7_75t_R _17332_ (.A1(net6367),
    .A2(net6465),
    .B(_01006_),
    .Y(_09162_));
 NAND2x1_ASAP7_75t_R _17333_ (.A(_09162_),
    .B(_09078_),
    .Y(_09163_));
 AOI21x1_ASAP7_75t_R _17335_ (.A1(_09161_),
    .A2(_09163_),
    .B(net6304),
    .Y(_09165_));
 AND2x2_ASAP7_75t_R _17336_ (.A(_09115_),
    .B(net5945),
    .Y(_09166_));
 NOR2x1_ASAP7_75t_R _17337_ (.A(net5926),
    .B(_09166_),
    .Y(_09167_));
 INVx2_ASAP7_75t_R _17338_ (.A(_09077_),
    .Y(_09168_));
 AO21x1_ASAP7_75t_R _17339_ (.A1(_09168_),
    .A2(net5923),
    .B(net5944),
    .Y(_09169_));
 AO21x1_ASAP7_75t_R _17340_ (.A1(_09167_),
    .A2(_09169_),
    .B(net5943),
    .Y(_09170_));
 OAI21x1_ASAP7_75t_R _17341_ (.A1(_09165_),
    .A2(_09170_),
    .B(_09121_),
    .Y(_09171_));
 AOI21x1_ASAP7_75t_R _17342_ (.A1(net5943),
    .A2(_09158_),
    .B(_09171_),
    .Y(_09172_));
 NOR2x1_ASAP7_75t_R _17343_ (.A(_09150_),
    .B(_09172_),
    .Y(_09173_));
 NOR2x1_ASAP7_75t_R _17344_ (.A(_09126_),
    .B(_09173_),
    .Y(_00008_));
 AO21x1_ASAP7_75t_R _17345_ (.A1(net6367),
    .A2(net6465),
    .B(_00997_),
    .Y(_09174_));
 NAND2x1_ASAP7_75t_R _17346_ (.A(net5946),
    .B(_09174_),
    .Y(_09175_));
 NOR2x1_ASAP7_75t_R _17347_ (.A(net5027),
    .B(_09175_),
    .Y(_09176_));
 AO21x1_ASAP7_75t_R _17348_ (.A1(_09063_),
    .A2(net6305),
    .B(net6304),
    .Y(_09177_));
 OAI21x1_ASAP7_75t_R _17350_ (.A1(_09176_),
    .A2(_09177_),
    .B(net6303),
    .Y(_09179_));
 NOR2x1_ASAP7_75t_R _17351_ (.A(_09039_),
    .B(net6308),
    .Y(_09180_));
 INVx1_ASAP7_75t_R _17352_ (.A(_09180_),
    .Y(_09181_));
 OA21x2_ASAP7_75t_R _17354_ (.A1(net5950),
    .A2(_09080_),
    .B(net5945),
    .Y(_09183_));
 AOI21x1_ASAP7_75t_R _17355_ (.A1(net5551),
    .A2(_09183_),
    .B(net5926),
    .Y(_09184_));
 OA21x2_ASAP7_75t_R _17356_ (.A1(net5944),
    .A2(_09181_),
    .B(_09184_),
    .Y(_09185_));
 OAI21x1_ASAP7_75t_R _17357_ (.A1(_09179_),
    .A2(_09185_),
    .B(net5943),
    .Y(_09186_));
 NAND2x1_ASAP7_75t_R _17358_ (.A(net6308),
    .B(net6310),
    .Y(_09187_));
 INVx1_ASAP7_75t_R _17359_ (.A(_09159_),
    .Y(_09188_));
 AO21x1_ASAP7_75t_R _17360_ (.A1(net5922),
    .A2(_09188_),
    .B(net5947),
    .Y(_09189_));
 AO21x1_ASAP7_75t_R _17362_ (.A1(net4598),
    .A2(net5237),
    .B(net6305),
    .Y(_09191_));
 AO21x1_ASAP7_75t_R _17364_ (.A1(_09189_),
    .A2(_09191_),
    .B(net5927),
    .Y(_09193_));
 NAND2x1_ASAP7_75t_R _17365_ (.A(net6309),
    .B(net6311),
    .Y(_09194_));
 NAND2x1_ASAP7_75t_R _17366_ (.A(_09194_),
    .B(_09136_),
    .Y(_09195_));
 AO21x1_ASAP7_75t_R _17367_ (.A1(net5556),
    .A2(net4787),
    .B(net5947),
    .Y(_09196_));
 AO21x1_ASAP7_75t_R _17368_ (.A1(_09195_),
    .A2(_09196_),
    .B(net6304),
    .Y(_09197_));
 AOI21x1_ASAP7_75t_R _17369_ (.A1(_09193_),
    .A2(_09197_),
    .B(net6303),
    .Y(_09198_));
 OAI21x1_ASAP7_75t_R _17370_ (.A1(_09186_),
    .A2(_09198_),
    .B(net5942),
    .Y(_09199_));
 NAND2x1_ASAP7_75t_R _17371_ (.A(net5317),
    .B(_08962_),
    .Y(_09200_));
 INVx1_ASAP7_75t_R _17372_ (.A(_09187_),
    .Y(_09201_));
 NOR2x1_ASAP7_75t_R _17373_ (.A(net5947),
    .B(_09201_),
    .Y(_09202_));
 AO221x1_ASAP7_75t_R _17374_ (.A1(net4598),
    .A2(_09136_),
    .B1(_09200_),
    .B2(_09202_),
    .C(net5927),
    .Y(_09203_));
 OA21x2_ASAP7_75t_R _17375_ (.A1(net4977),
    .A2(net6305),
    .B(net5927),
    .Y(_09204_));
 NOR2x1_ASAP7_75t_R _17376_ (.A(net6309),
    .B(_08962_),
    .Y(_09205_));
 INVx1_ASAP7_75t_R _17377_ (.A(_09205_),
    .Y(_09206_));
 AO21x1_ASAP7_75t_R _17378_ (.A1(_09206_),
    .A2(_09194_),
    .B(net5948),
    .Y(_09207_));
 AOI21x1_ASAP7_75t_R _17379_ (.A1(_09204_),
    .A2(_09207_),
    .B(net5924),
    .Y(_09208_));
 AO21x1_ASAP7_75t_R _17380_ (.A1(net5552),
    .A2(net5237),
    .B(net5947),
    .Y(_09209_));
 AOI21x1_ASAP7_75t_R _17381_ (.A1(_01009_),
    .A2(net5947),
    .B(net5927),
    .Y(_09210_));
 AO21x1_ASAP7_75t_R _17383_ (.A1(_09209_),
    .A2(_09210_),
    .B(net6303),
    .Y(_09212_));
 AND3x1_ASAP7_75t_R _17385_ (.A(net5236),
    .B(net5947),
    .C(net4787),
    .Y(_09214_));
 AO21x1_ASAP7_75t_R _17386_ (.A1(_09133_),
    .A2(net5237),
    .B(net5948),
    .Y(_09215_));
 NAND2x1_ASAP7_75t_R _17387_ (.A(net5929),
    .B(_09215_),
    .Y(_09216_));
 NOR2x1_ASAP7_75t_R _17388_ (.A(_09214_),
    .B(_09216_),
    .Y(_09217_));
 OAI21x1_ASAP7_75t_R _17390_ (.A1(_09212_),
    .A2(_09217_),
    .B(net5554),
    .Y(_09219_));
 AOI21x1_ASAP7_75t_R _17391_ (.A1(_09203_),
    .A2(_09208_),
    .B(_09219_),
    .Y(_09220_));
 AO21x1_ASAP7_75t_R _17392_ (.A1(net5555),
    .A2(_09206_),
    .B(net6303),
    .Y(_09221_));
 INVx1_ASAP7_75t_R _17393_ (.A(_09151_),
    .Y(_09222_));
 NOR2x1_ASAP7_75t_R _17394_ (.A(_09222_),
    .B(_09111_),
    .Y(_09223_));
 OR3x1_ASAP7_75t_R _17395_ (.A(_09221_),
    .B(net5930),
    .C(_09223_),
    .Y(_09224_));
 AO21x1_ASAP7_75t_R _17396_ (.A1(net5556),
    .A2(_09048_),
    .B(net5948),
    .Y(_09225_));
 AO21x1_ASAP7_75t_R _17397_ (.A1(_09181_),
    .A2(_09065_),
    .B(net6306),
    .Y(_09226_));
 AO21x1_ASAP7_75t_R _17398_ (.A1(_09225_),
    .A2(_09226_),
    .B(net5928),
    .Y(_09227_));
 AOI21x1_ASAP7_75t_R _17399_ (.A1(_01015_),
    .A2(net5946),
    .B(net6304),
    .Y(_09228_));
 OAI21x1_ASAP7_75t_R _17400_ (.A1(net4972),
    .A2(_09105_),
    .B(net6306),
    .Y(_09229_));
 OA22x2_ASAP7_75t_R _17401_ (.A1(_09228_),
    .A2(net6303),
    .B1(_09229_),
    .B2(net6304),
    .Y(_09230_));
 NAND2x1_ASAP7_75t_R _17402_ (.A(_09227_),
    .B(_09230_),
    .Y(_09231_));
 AOI21x1_ASAP7_75t_R _17403_ (.A1(_09224_),
    .A2(_09231_),
    .B(net5943),
    .Y(_09232_));
 AND2x2_ASAP7_75t_R _17404_ (.A(net5555),
    .B(_09162_),
    .Y(_09233_));
 OAI21x1_ASAP7_75t_R _17406_ (.A1(_09233_),
    .A2(_09223_),
    .B(net5930),
    .Y(_09235_));
 AO21x1_ASAP7_75t_R _17407_ (.A1(net5922),
    .A2(_09095_),
    .B(net5948),
    .Y(_09236_));
 AO21x1_ASAP7_75t_R _17409_ (.A1(_09188_),
    .A2(net5025),
    .B(net6305),
    .Y(_09238_));
 AO21x1_ASAP7_75t_R _17410_ (.A1(_09236_),
    .A2(_09238_),
    .B(net5927),
    .Y(_09239_));
 AOI21x1_ASAP7_75t_R _17411_ (.A1(_09235_),
    .A2(_09239_),
    .B(net5924),
    .Y(_09240_));
 INVx1_ASAP7_75t_R _17412_ (.A(_01007_),
    .Y(_09241_));
 OAI21x1_ASAP7_75t_R _17413_ (.A1(_09241_),
    .A2(net5951),
    .B(net6307),
    .Y(_09242_));
 INVx1_ASAP7_75t_R _17414_ (.A(_09242_),
    .Y(_09243_));
 AOI211x1_ASAP7_75t_R _17415_ (.A1(_09243_),
    .A2(net5236),
    .B(_09176_),
    .C(net5927),
    .Y(_09244_));
 AO21x1_ASAP7_75t_R _17416_ (.A1(net5922),
    .A2(_09181_),
    .B(net5944),
    .Y(_09245_));
 NOR2x1_ASAP7_75t_R _17417_ (.A(net6304),
    .B(net4599),
    .Y(_09246_));
 AO21x1_ASAP7_75t_R _17418_ (.A1(_09245_),
    .A2(_09246_),
    .B(net6303),
    .Y(_09247_));
 OAI21x1_ASAP7_75t_R _17419_ (.A1(_09244_),
    .A2(_09247_),
    .B(net5943),
    .Y(_09248_));
 OAI21x1_ASAP7_75t_R _17421_ (.A1(_09240_),
    .A2(_09248_),
    .B(net5550),
    .Y(_09250_));
 OAI22x1_ASAP7_75t_R _17422_ (.A1(_09199_),
    .A2(_09220_),
    .B1(_09232_),
    .B2(_09250_),
    .Y(_00009_));
 INVx1_ASAP7_75t_R _17423_ (.A(_09092_),
    .Y(_09251_));
 NOR2x1_ASAP7_75t_R _17424_ (.A(_08968_),
    .B(_09251_),
    .Y(_09252_));
 NAND2x1_ASAP7_75t_R _17425_ (.A(_09082_),
    .B(net4713),
    .Y(_09253_));
 NAND2x1_ASAP7_75t_R _17426_ (.A(net5025),
    .B(_09078_),
    .Y(_09254_));
 AO21x1_ASAP7_75t_R _17427_ (.A1(_09253_),
    .A2(_09254_),
    .B(net6304),
    .Y(_09255_));
 INVx1_ASAP7_75t_R _17428_ (.A(_09143_),
    .Y(_09256_));
 NOR2x1_ASAP7_75t_R _17430_ (.A(net6306),
    .B(_09222_),
    .Y(_09258_));
 AO21x1_ASAP7_75t_R _17431_ (.A1(net6367),
    .A2(net6465),
    .B(_00999_),
    .Y(_09259_));
 AO21x1_ASAP7_75t_R _17432_ (.A1(_09060_),
    .A2(_09259_),
    .B(_09043_),
    .Y(_09260_));
 AO21x1_ASAP7_75t_R _17433_ (.A1(net5235),
    .A2(_09258_),
    .B(_09260_),
    .Y(_09261_));
 AOI21x1_ASAP7_75t_R _17434_ (.A1(_09255_),
    .A2(_09261_),
    .B(net5924),
    .Y(_09262_));
 INVx1_ASAP7_75t_R _17435_ (.A(_01002_),
    .Y(_09263_));
 AO21x1_ASAP7_75t_R _17436_ (.A1(net6367),
    .A2(net6465),
    .B(_09263_),
    .Y(_09264_));
 AND2x2_ASAP7_75t_R _17437_ (.A(_09264_),
    .B(net5948),
    .Y(_09265_));
 NAND2x1_ASAP7_75t_R _17438_ (.A(net5552),
    .B(_09265_),
    .Y(_09266_));
 AO21x1_ASAP7_75t_R _17439_ (.A1(_09256_),
    .A2(net5237),
    .B(net5947),
    .Y(_09267_));
 AO21x1_ASAP7_75t_R _17440_ (.A1(_09266_),
    .A2(_09267_),
    .B(net6304),
    .Y(_09268_));
 AO21x1_ASAP7_75t_R _17441_ (.A1(net5556),
    .A2(net5237),
    .B(net6306),
    .Y(_09269_));
 AO21x1_ASAP7_75t_R _17442_ (.A1(_09256_),
    .A2(_09259_),
    .B(net5947),
    .Y(_09270_));
 AO21x1_ASAP7_75t_R _17443_ (.A1(_09269_),
    .A2(_09270_),
    .B(net5929),
    .Y(_09271_));
 AOI21x1_ASAP7_75t_R _17444_ (.A1(_09268_),
    .A2(_09271_),
    .B(net6303),
    .Y(_09272_));
 NOR3x1_ASAP7_75t_R _17445_ (.A(_09262_),
    .B(_09272_),
    .C(net5554),
    .Y(_09273_));
 INVx1_ASAP7_75t_R _17446_ (.A(_09259_),
    .Y(_09274_));
 OAI21x1_ASAP7_75t_R _17447_ (.A1(_09063_),
    .A2(_09274_),
    .B(net6305),
    .Y(_09275_));
 AO21x1_ASAP7_75t_R _17448_ (.A1(net5553),
    .A2(_09065_),
    .B(net6305),
    .Y(_09276_));
 AOI21x1_ASAP7_75t_R _17449_ (.A1(_09275_),
    .A2(_09276_),
    .B(net5929),
    .Y(_09277_));
 AO21x1_ASAP7_75t_R _17450_ (.A1(_09133_),
    .A2(net5237),
    .B(net6306),
    .Y(_09278_));
 NAND2x1_ASAP7_75t_R _17451_ (.A(_08962_),
    .B(net5931),
    .Y(_09279_));
 AO21x1_ASAP7_75t_R _17452_ (.A1(_09279_),
    .A2(net5025),
    .B(net5948),
    .Y(_09280_));
 AOI21x1_ASAP7_75t_R _17453_ (.A1(_09278_),
    .A2(_09280_),
    .B(net6304),
    .Y(_09281_));
 OAI21x1_ASAP7_75t_R _17454_ (.A1(_09277_),
    .A2(_09281_),
    .B(net5924),
    .Y(_09282_));
 NOR2x1_ASAP7_75t_R _17455_ (.A(net5316),
    .B(net5951),
    .Y(_09283_));
 OAI21x1_ASAP7_75t_R _17456_ (.A1(net4788),
    .A2(_09205_),
    .B(net6306),
    .Y(_09284_));
 OA21x2_ASAP7_75t_R _17457_ (.A1(_09117_),
    .A2(_09283_),
    .B(_09284_),
    .Y(_09285_));
 INVx1_ASAP7_75t_R _17458_ (.A(_09175_),
    .Y(_09286_));
 AOI21x1_ASAP7_75t_R _17459_ (.A1(net5236),
    .A2(_09286_),
    .B(_09083_),
    .Y(_09287_));
 AOI21x1_ASAP7_75t_R _17460_ (.A1(net5928),
    .A2(_09287_),
    .B(_09124_),
    .Y(_09288_));
 OAI21x1_ASAP7_75t_R _17461_ (.A1(net5928),
    .A2(_09285_),
    .B(_09288_),
    .Y(_09289_));
 NAND2x1_ASAP7_75t_R _17462_ (.A(_09282_),
    .B(_09289_),
    .Y(_09290_));
 OAI21x1_ASAP7_75t_R _17463_ (.A1(net5943),
    .A2(_09290_),
    .B(net5550),
    .Y(_09291_));
 NAND2x1_ASAP7_75t_R _17464_ (.A(net5946),
    .B(net5026),
    .Y(_09292_));
 AO21x1_ASAP7_75t_R _17465_ (.A1(net5553),
    .A2(_09162_),
    .B(net5946),
    .Y(_09293_));
 OA21x2_ASAP7_75t_R _17466_ (.A1(_09046_),
    .A2(_09292_),
    .B(_09293_),
    .Y(_09294_));
 NAND2x1_ASAP7_75t_R _17467_ (.A(_01015_),
    .B(net6307),
    .Y(_09295_));
 NAND2x1_ASAP7_75t_R _17468_ (.A(_09194_),
    .B(_09206_),
    .Y(_09296_));
 AOI21x1_ASAP7_75t_R _17469_ (.A1(net5946),
    .A2(_09296_),
    .B(net6304),
    .Y(_09297_));
 AOI21x1_ASAP7_75t_R _17470_ (.A1(_09295_),
    .A2(_09297_),
    .B(net6303),
    .Y(_09298_));
 OA21x2_ASAP7_75t_R _17471_ (.A1(net5925),
    .A2(_09294_),
    .B(_09298_),
    .Y(_09299_));
 AO21x1_ASAP7_75t_R _17472_ (.A1(_09133_),
    .A2(net5025),
    .B(net6306),
    .Y(_09300_));
 INVx1_ASAP7_75t_R _17473_ (.A(_01014_),
    .Y(_09301_));
 NAND2x1_ASAP7_75t_R _17474_ (.A(_09301_),
    .B(net6306),
    .Y(_09302_));
 AND3x1_ASAP7_75t_R _17475_ (.A(_09300_),
    .B(net5929),
    .C(_09302_),
    .Y(_09303_));
 AO21x1_ASAP7_75t_R _17476_ (.A1(net5552),
    .A2(net4787),
    .B(net5947),
    .Y(_09304_));
 AO21x1_ASAP7_75t_R _17477_ (.A1(net5556),
    .A2(_01011_),
    .B(net6305),
    .Y(_09305_));
 NAND2x1_ASAP7_75t_R _17478_ (.A(_09304_),
    .B(_09305_),
    .Y(_09306_));
 OAI21x1_ASAP7_75t_R _17479_ (.A1(net5929),
    .A2(_09306_),
    .B(net6303),
    .Y(_09307_));
 OAI21x1_ASAP7_75t_R _17480_ (.A1(_09303_),
    .A2(_09307_),
    .B(net5943),
    .Y(_09308_));
 NAND2x1_ASAP7_75t_R _17481_ (.A(net6305),
    .B(net4973),
    .Y(_09309_));
 NAND2x1_ASAP7_75t_R _17482_ (.A(net4970),
    .B(_09078_),
    .Y(_09310_));
 AOI21x1_ASAP7_75t_R _17483_ (.A1(_09309_),
    .A2(_09310_),
    .B(net6304),
    .Y(_09311_));
 NAND2x1_ASAP7_75t_R _17484_ (.A(net5556),
    .B(_09286_),
    .Y(_09312_));
 AOI21x1_ASAP7_75t_R _17485_ (.A1(_09229_),
    .A2(_09312_),
    .B(net5928),
    .Y(_09313_));
 OAI21x1_ASAP7_75t_R _17486_ (.A1(_09311_),
    .A2(_09313_),
    .B(net6303),
    .Y(_09314_));
 OA21x2_ASAP7_75t_R _17487_ (.A1(_01011_),
    .A2(net5947),
    .B(net6304),
    .Y(_09315_));
 AOI21x1_ASAP7_75t_R _17488_ (.A1(_09315_),
    .A2(_09276_),
    .B(net6303),
    .Y(_09316_));
 NAND2x1_ASAP7_75t_R _17489_ (.A(_01013_),
    .B(net5945),
    .Y(_09317_));
 NAND2x1_ASAP7_75t_R _17490_ (.A(_09317_),
    .B(_09153_),
    .Y(_09318_));
 OR2x2_ASAP7_75t_R _17491_ (.A(net6304),
    .B(_09318_),
    .Y(_09319_));
 AOI21x1_ASAP7_75t_R _17492_ (.A1(_09316_),
    .A2(_09319_),
    .B(net5943),
    .Y(_09320_));
 AOI21x1_ASAP7_75t_R _17493_ (.A1(_09314_),
    .A2(_09320_),
    .B(_09121_),
    .Y(_09321_));
 OAI21x1_ASAP7_75t_R _17494_ (.A1(_09299_),
    .A2(_09308_),
    .B(_09321_),
    .Y(_09322_));
 OAI21x1_ASAP7_75t_R _17495_ (.A1(_09273_),
    .A2(_09291_),
    .B(_09322_),
    .Y(_00010_));
 NOR2x1_ASAP7_75t_R _17496_ (.A(net5944),
    .B(_09168_),
    .Y(_09323_));
 AO21x1_ASAP7_75t_R _17497_ (.A1(_09323_),
    .A2(net6303),
    .B(_09102_),
    .Y(_09324_));
 OR3x1_ASAP7_75t_R _17498_ (.A(net5950),
    .B(_09076_),
    .C(net6307),
    .Y(_09325_));
 OAI21x1_ASAP7_75t_R _17499_ (.A1(net5238),
    .A2(_09154_),
    .B(net6307),
    .Y(_09326_));
 AOI21x1_ASAP7_75t_R _17500_ (.A1(_09325_),
    .A2(_09326_),
    .B(net6303),
    .Y(_09327_));
 OAI21x1_ASAP7_75t_R _17501_ (.A1(_09324_),
    .A2(_09327_),
    .B(net6304),
    .Y(_09328_));
 NOR2x1_ASAP7_75t_R _17502_ (.A(net4788),
    .B(_09071_),
    .Y(_09329_));
 AO21x1_ASAP7_75t_R _17503_ (.A1(net5556),
    .A2(_09183_),
    .B(_09329_),
    .Y(_09330_));
 OA21x2_ASAP7_75t_R _17504_ (.A1(_09256_),
    .A2(net6305),
    .B(net6303),
    .Y(_09331_));
 AOI21x1_ASAP7_75t_R _17505_ (.A1(_09253_),
    .A2(_09331_),
    .B(net6304),
    .Y(_09332_));
 OAI21x1_ASAP7_75t_R _17506_ (.A1(net6303),
    .A2(_09330_),
    .B(_09332_),
    .Y(_09333_));
 AOI21x1_ASAP7_75t_R _17507_ (.A1(_09328_),
    .A2(_09333_),
    .B(net5943),
    .Y(_09334_));
 NAND2x1_ASAP7_75t_R _17508_ (.A(_09124_),
    .B(_09260_),
    .Y(_09335_));
 NOR2x1_ASAP7_75t_R _17509_ (.A(net4971),
    .B(_09117_),
    .Y(_09336_));
 INVx1_ASAP7_75t_R _17510_ (.A(_09336_),
    .Y(_09337_));
 AOI21x1_ASAP7_75t_R _17511_ (.A1(_09229_),
    .A2(_09337_),
    .B(net6304),
    .Y(_09338_));
 OAI21x1_ASAP7_75t_R _17512_ (.A1(_09335_),
    .A2(_09338_),
    .B(net5943),
    .Y(_09339_));
 NAND2x1_ASAP7_75t_R _17513_ (.A(_09207_),
    .B(_09137_),
    .Y(_09340_));
 AO21x1_ASAP7_75t_R _17514_ (.A1(_09036_),
    .A2(_09259_),
    .B(net5948),
    .Y(_09341_));
 AO21x1_ASAP7_75t_R _17515_ (.A1(net5951),
    .A2(net5570),
    .B(net6307),
    .Y(_09342_));
 OA21x2_ASAP7_75t_R _17516_ (.A1(_09342_),
    .A2(_09201_),
    .B(net6304),
    .Y(_09343_));
 NAND2x1_ASAP7_75t_R _17517_ (.A(_09341_),
    .B(_09343_),
    .Y(_09344_));
 AOI21x1_ASAP7_75t_R _17518_ (.A1(_09340_),
    .A2(_09344_),
    .B(net5924),
    .Y(_09345_));
 NOR2x1_ASAP7_75t_R _17519_ (.A(_09339_),
    .B(_09345_),
    .Y(_09346_));
 OAI21x1_ASAP7_75t_R _17520_ (.A1(_09334_),
    .A2(_09346_),
    .B(_09121_),
    .Y(_09347_));
 AND3x1_ASAP7_75t_R _17521_ (.A(_09168_),
    .B(net5944),
    .C(net5923),
    .Y(_09348_));
 AO21x1_ASAP7_75t_R _17522_ (.A1(_09053_),
    .A2(net5922),
    .B(net5944),
    .Y(_09349_));
 NAND2x1_ASAP7_75t_R _17523_ (.A(net5926),
    .B(_09349_),
    .Y(_09350_));
 AO21x1_ASAP7_75t_R _17524_ (.A1(net5556),
    .A2(_01011_),
    .B(net5944),
    .Y(_09351_));
 AOI21x1_ASAP7_75t_R _17525_ (.A1(_09167_),
    .A2(_09351_),
    .B(net6303),
    .Y(_09352_));
 OAI21x1_ASAP7_75t_R _17526_ (.A1(_09348_),
    .A2(_09350_),
    .B(_09352_),
    .Y(_09353_));
 NAND2x1_ASAP7_75t_R _17527_ (.A(net5236),
    .B(_09265_),
    .Y(_09354_));
 AOI21x1_ASAP7_75t_R _17528_ (.A1(_09284_),
    .A2(_09354_),
    .B(net6304),
    .Y(_09355_));
 OAI21x1_ASAP7_75t_R _17529_ (.A1(_09046_),
    .A2(_09201_),
    .B(net6305),
    .Y(_09356_));
 AO21x1_ASAP7_75t_R _17530_ (.A1(_09188_),
    .A2(net4787),
    .B(net6305),
    .Y(_09357_));
 AOI21x1_ASAP7_75t_R _17531_ (.A1(_09356_),
    .A2(_09357_),
    .B(net5927),
    .Y(_09358_));
 OAI21x1_ASAP7_75t_R _17532_ (.A1(_09355_),
    .A2(_09358_),
    .B(net6303),
    .Y(_09359_));
 AOI21x1_ASAP7_75t_R _17533_ (.A1(_09353_),
    .A2(_09359_),
    .B(net5943),
    .Y(_09360_));
 OA21x2_ASAP7_75t_R _17534_ (.A1(net5950),
    .A2(net5319),
    .B(net5945),
    .Y(_09361_));
 NAND2x1_ASAP7_75t_R _17535_ (.A(_09036_),
    .B(net4713),
    .Y(_09362_));
 AOI21x1_ASAP7_75t_R _17536_ (.A1(_09362_),
    .A2(_09184_),
    .B(net6303),
    .Y(_09363_));
 OAI21x1_ASAP7_75t_R _17537_ (.A1(_09361_),
    .A2(_09350_),
    .B(_09363_),
    .Y(_09364_));
 OAI21x1_ASAP7_75t_R _17538_ (.A1(_09046_),
    .A2(_09066_),
    .B(net5944),
    .Y(_09365_));
 AO21x1_ASAP7_75t_R _17539_ (.A1(_09181_),
    .A2(net5024),
    .B(net5944),
    .Y(_09366_));
 AOI21x1_ASAP7_75t_R _17540_ (.A1(_09365_),
    .A2(_09366_),
    .B(net6304),
    .Y(_09367_));
 OAI21x1_ASAP7_75t_R _17541_ (.A1(net4788),
    .A2(net5238),
    .B(net6307),
    .Y(_09368_));
 NAND2x1_ASAP7_75t_R _17542_ (.A(net5931),
    .B(net5952),
    .Y(_09369_));
 AO21x1_ASAP7_75t_R _17543_ (.A1(_09369_),
    .A2(net5922),
    .B(net6307),
    .Y(_09370_));
 AOI21x1_ASAP7_75t_R _17544_ (.A1(_09368_),
    .A2(_09370_),
    .B(net5926),
    .Y(_09371_));
 OAI21x1_ASAP7_75t_R _17545_ (.A1(_09367_),
    .A2(_09371_),
    .B(net6303),
    .Y(_09372_));
 AOI21x1_ASAP7_75t_R _17546_ (.A1(_09364_),
    .A2(_09372_),
    .B(net5554),
    .Y(_09373_));
 OAI21x1_ASAP7_75t_R _17547_ (.A1(_09360_),
    .A2(_09373_),
    .B(net5942),
    .Y(_09374_));
 NAND2x1_ASAP7_75t_R _17548_ (.A(_09347_),
    .B(_09374_),
    .Y(_00011_));
 NOR2x1_ASAP7_75t_R _17549_ (.A(net6306),
    .B(net4971),
    .Y(_09375_));
 NOR2x1_ASAP7_75t_R _17550_ (.A(net5239),
    .B(net4711),
    .Y(_09376_));
 AO21x1_ASAP7_75t_R _17551_ (.A1(_09376_),
    .A2(net6304),
    .B(net5554),
    .Y(_09377_));
 AO21x1_ASAP7_75t_R _17552_ (.A1(net5556),
    .A2(_01016_),
    .B(net6306),
    .Y(_09378_));
 AND3x1_ASAP7_75t_R _17553_ (.A(_09225_),
    .B(_09378_),
    .C(net5930),
    .Y(_09379_));
 OAI21x1_ASAP7_75t_R _17554_ (.A1(_09377_),
    .A2(_09379_),
    .B(net6303),
    .Y(_09380_));
 AO21x1_ASAP7_75t_R _17555_ (.A1(net5949),
    .A2(net5320),
    .B(net5945),
    .Y(_09381_));
 INVx1_ASAP7_75t_R _17556_ (.A(_09381_),
    .Y(_09382_));
 AOI22x1_ASAP7_75t_R _17557_ (.A1(net4714),
    .A2(net5240),
    .B1(net4787),
    .B2(_09382_),
    .Y(_09383_));
 NOR2x1_ASAP7_75t_R _17558_ (.A(net6306),
    .B(_09127_),
    .Y(_09384_));
 OR3x1_ASAP7_75t_R _17559_ (.A(_09146_),
    .B(_09043_),
    .C(net5549),
    .Y(_09385_));
 OAI21x1_ASAP7_75t_R _17560_ (.A1(net4786),
    .A2(_09385_),
    .B(net5554),
    .Y(_09386_));
 AOI21x1_ASAP7_75t_R _17561_ (.A1(net5928),
    .A2(_09383_),
    .B(_09386_),
    .Y(_09387_));
 OAI21x1_ASAP7_75t_R _17562_ (.A1(_09380_),
    .A2(_09387_),
    .B(net5942),
    .Y(_09388_));
 NAND2x1_ASAP7_75t_R _17563_ (.A(net6304),
    .B(_09275_),
    .Y(_09389_));
 AO21x1_ASAP7_75t_R _17564_ (.A1(net4714),
    .A2(net5923),
    .B(_09389_),
    .Y(_09390_));
 AND3x1_ASAP7_75t_R _17565_ (.A(_09135_),
    .B(net5948),
    .C(net5923),
    .Y(_09391_));
 OA21x2_ASAP7_75t_R _17566_ (.A1(_09216_),
    .A2(_09391_),
    .B(net5554),
    .Y(_09392_));
 NAND2x1_ASAP7_75t_R _17567_ (.A(_09206_),
    .B(net5555),
    .Y(_09393_));
 AOI21x1_ASAP7_75t_R _17568_ (.A1(_09393_),
    .A2(_09297_),
    .B(net5554),
    .Y(_09394_));
 AND3x1_ASAP7_75t_R _17569_ (.A(_09279_),
    .B(net5946),
    .C(_09048_),
    .Y(_09395_));
 NAND2x1_ASAP7_75t_R _17570_ (.A(net6311),
    .B(net5931),
    .Y(_09396_));
 NAND2x1_ASAP7_75t_R _17571_ (.A(net5553),
    .B(_09396_),
    .Y(_09397_));
 AND2x2_ASAP7_75t_R _17572_ (.A(_09397_),
    .B(net6307),
    .Y(_09398_));
 OAI21x1_ASAP7_75t_R _17573_ (.A1(_09395_),
    .A2(_09398_),
    .B(net6304),
    .Y(_09399_));
 AO21x1_ASAP7_75t_R _17574_ (.A1(_09394_),
    .A2(_09399_),
    .B(net6303),
    .Y(_09400_));
 AOI21x1_ASAP7_75t_R _17575_ (.A1(_09390_),
    .A2(_09392_),
    .B(_09400_),
    .Y(_09401_));
 INVx1_ASAP7_75t_R _17576_ (.A(_09117_),
    .Y(_09402_));
 AO21x1_ASAP7_75t_R _17577_ (.A1(_09402_),
    .A2(net5240),
    .B(net5925),
    .Y(_09403_));
 OAI21x1_ASAP7_75t_R _17578_ (.A1(_09398_),
    .A2(_09403_),
    .B(net5554),
    .Y(_09404_));
 AND3x1_ASAP7_75t_R _17579_ (.A(_09057_),
    .B(net5928),
    .C(_09110_),
    .Y(_09405_));
 NOR2x1_ASAP7_75t_R _17580_ (.A(_09404_),
    .B(_09405_),
    .Y(_09406_));
 INVx1_ASAP7_75t_R _17581_ (.A(_09081_),
    .Y(_09407_));
 AOI22x1_ASAP7_75t_R _17582_ (.A1(net5555),
    .A2(_09407_),
    .B1(net6308),
    .B2(net5948),
    .Y(_09408_));
 AO21x1_ASAP7_75t_R _17583_ (.A1(_09408_),
    .A2(net5930),
    .B(net5554),
    .Y(_09409_));
 AND3x1_ASAP7_75t_R _17584_ (.A(_09206_),
    .B(net6306),
    .C(_09135_),
    .Y(_09410_));
 NOR3x1_ASAP7_75t_R _17585_ (.A(_09410_),
    .B(net5930),
    .C(_09223_),
    .Y(_09411_));
 OAI21x1_ASAP7_75t_R _17586_ (.A1(_09409_),
    .A2(_09411_),
    .B(net5924),
    .Y(_09412_));
 INVx1_ASAP7_75t_R _17587_ (.A(_09142_),
    .Y(_09413_));
 AND3x1_ASAP7_75t_R _17588_ (.A(_09200_),
    .B(net6305),
    .C(_09127_),
    .Y(_09414_));
 NAND2x1_ASAP7_75t_R _17589_ (.A(_09242_),
    .B(_09175_),
    .Y(_09415_));
 OA21x2_ASAP7_75t_R _17590_ (.A1(_09415_),
    .A2(net5925),
    .B(net5943),
    .Y(_09416_));
 OAI21x1_ASAP7_75t_R _17591_ (.A1(_09413_),
    .A2(_09414_),
    .B(_09416_),
    .Y(_09417_));
 NAND2x1_ASAP7_75t_R _17592_ (.A(net5553),
    .B(_09375_),
    .Y(_09418_));
 OA21x2_ASAP7_75t_R _17593_ (.A1(_09133_),
    .A2(net5948),
    .B(net6304),
    .Y(_09419_));
 NAND2x1_ASAP7_75t_R _17594_ (.A(_09418_),
    .B(_09419_),
    .Y(_09420_));
 OA21x2_ASAP7_75t_R _17595_ (.A1(net5241),
    .A2(net5946),
    .B(net5925),
    .Y(_09421_));
 AOI21x1_ASAP7_75t_R _17596_ (.A1(_09292_),
    .A2(_09421_),
    .B(net5943),
    .Y(_09422_));
 AOI21x1_ASAP7_75t_R _17597_ (.A1(_09420_),
    .A2(_09422_),
    .B(net5924),
    .Y(_09423_));
 AOI21x1_ASAP7_75t_R _17598_ (.A1(_09417_),
    .A2(_09423_),
    .B(net5942),
    .Y(_09424_));
 OAI21x1_ASAP7_75t_R _17599_ (.A1(_09406_),
    .A2(_09412_),
    .B(_09424_),
    .Y(_09425_));
 OAI21x1_ASAP7_75t_R _17600_ (.A1(_09388_),
    .A2(_09401_),
    .B(_09425_),
    .Y(_00012_));
 AO21x1_ASAP7_75t_R _17601_ (.A1(net5949),
    .A2(_09039_),
    .B(net5945),
    .Y(_09426_));
 NAND2x1_ASAP7_75t_R _17602_ (.A(net5571),
    .B(net5945),
    .Y(_09427_));
 AO21x1_ASAP7_75t_R _17603_ (.A1(_09426_),
    .A2(_09427_),
    .B(net6303),
    .Y(_09428_));
 AOI221x1_ASAP7_75t_R _17604_ (.A1(_09141_),
    .A2(_09083_),
    .B1(net6303),
    .B2(_09402_),
    .C(net6304),
    .Y(_09429_));
 OAI21x1_ASAP7_75t_R _17605_ (.A1(net5027),
    .A2(net5238),
    .B(net5945),
    .Y(_09430_));
 AO21x1_ASAP7_75t_R _17606_ (.A1(_09168_),
    .A2(_09259_),
    .B(net5945),
    .Y(_09431_));
 AOI21x1_ASAP7_75t_R _17607_ (.A1(_09430_),
    .A2(_09431_),
    .B(net6303),
    .Y(_09432_));
 OAI21x1_ASAP7_75t_R _17608_ (.A1(_09146_),
    .A2(_09183_),
    .B(net6303),
    .Y(_09433_));
 NAND2x1_ASAP7_75t_R _17609_ (.A(net6304),
    .B(_09433_),
    .Y(_09434_));
 OAI21x1_ASAP7_75t_R _17610_ (.A1(_09432_),
    .A2(_09434_),
    .B(net5554),
    .Y(_09435_));
 AOI21x1_ASAP7_75t_R _17611_ (.A1(_09428_),
    .A2(_09429_),
    .B(_09435_),
    .Y(_09436_));
 AND3x1_ASAP7_75t_R _17612_ (.A(_09082_),
    .B(net6305),
    .C(_09264_),
    .Y(_09437_));
 AO21x1_ASAP7_75t_R _17613_ (.A1(_09181_),
    .A2(_09259_),
    .B(net5945),
    .Y(_09438_));
 OA21x2_ASAP7_75t_R _17614_ (.A1(_09427_),
    .A2(_08962_),
    .B(net6304),
    .Y(_09439_));
 AOI21x1_ASAP7_75t_R _17615_ (.A1(_09438_),
    .A2(_09439_),
    .B(net6303),
    .Y(_09440_));
 OAI21x1_ASAP7_75t_R _17616_ (.A1(_09437_),
    .A2(_09413_),
    .B(_09440_),
    .Y(_09441_));
 AO22x1_ASAP7_75t_R _17617_ (.A1(net4713),
    .A2(net5551),
    .B1(_09361_),
    .B2(_09168_),
    .Y(_09442_));
 OA21x2_ASAP7_75t_R _17618_ (.A1(net5952),
    .A2(net6307),
    .B(net5926),
    .Y(_09443_));
 AOI21x1_ASAP7_75t_R _17619_ (.A1(_09061_),
    .A2(_09443_),
    .B(_09124_),
    .Y(_09444_));
 OAI21x1_ASAP7_75t_R _17620_ (.A1(net5926),
    .A2(_09442_),
    .B(_09444_),
    .Y(_09445_));
 AOI21x1_ASAP7_75t_R _17621_ (.A1(_09441_),
    .A2(_09445_),
    .B(net5554),
    .Y(_09446_));
 OAI21x1_ASAP7_75t_R _17622_ (.A1(_09436_),
    .A2(_09446_),
    .B(_09121_),
    .Y(_09447_));
 NAND2x1_ASAP7_75t_R _17623_ (.A(net4976),
    .B(net4713),
    .Y(_09448_));
 NAND2x1_ASAP7_75t_R _17624_ (.A(net5556),
    .B(_09265_),
    .Y(_09449_));
 AOI21x1_ASAP7_75t_R _17625_ (.A1(_09448_),
    .A2(_09449_),
    .B(net5927),
    .Y(_09450_));
 NAND2x1_ASAP7_75t_R _17626_ (.A(_09200_),
    .B(_09183_),
    .Y(_09451_));
 AOI21x1_ASAP7_75t_R _17627_ (.A1(_09152_),
    .A2(_09451_),
    .B(net6304),
    .Y(_09452_));
 OAI21x1_ASAP7_75t_R _17628_ (.A1(_09450_),
    .A2(_09452_),
    .B(net6303),
    .Y(_09453_));
 AO21x1_ASAP7_75t_R _17629_ (.A1(_09200_),
    .A2(net6305),
    .B(_09066_),
    .Y(_09454_));
 AOI21x1_ASAP7_75t_R _17630_ (.A1(net6305),
    .A2(_09168_),
    .B(net6304),
    .Y(_09455_));
 AO21x1_ASAP7_75t_R _17631_ (.A1(_09132_),
    .A2(_09256_),
    .B(net6305),
    .Y(_09456_));
 AOI21x1_ASAP7_75t_R _17632_ (.A1(_09455_),
    .A2(_09456_),
    .B(net6303),
    .Y(_09457_));
 OAI21x1_ASAP7_75t_R _17633_ (.A1(net5927),
    .A2(_09454_),
    .B(_09457_),
    .Y(_09458_));
 AOI21x1_ASAP7_75t_R _17634_ (.A1(_09453_),
    .A2(_09458_),
    .B(net5554),
    .Y(_09459_));
 INVx1_ASAP7_75t_R _17635_ (.A(_09384_),
    .Y(_09460_));
 NAND2x1_ASAP7_75t_R _17636_ (.A(_09279_),
    .B(_09243_),
    .Y(_09461_));
 AOI21x1_ASAP7_75t_R _17637_ (.A1(_09460_),
    .A2(_09461_),
    .B(net5925),
    .Y(_09462_));
 AO21x1_ASAP7_75t_R _17638_ (.A1(net6306),
    .A2(_09259_),
    .B(net6304),
    .Y(_09463_));
 AOI21x1_ASAP7_75t_R _17639_ (.A1(_09048_),
    .A2(net4600),
    .B(_09463_),
    .Y(_09464_));
 OAI21x1_ASAP7_75t_R _17640_ (.A1(_09462_),
    .A2(_09464_),
    .B(net5924),
    .Y(_09465_));
 AO21x1_ASAP7_75t_R _17641_ (.A1(net6309),
    .A2(net5946),
    .B(net6304),
    .Y(_09466_));
 AOI21x1_ASAP7_75t_R _17642_ (.A1(net6307),
    .A2(_09397_),
    .B(_09466_),
    .Y(_09467_));
 OAI21x1_ASAP7_75t_R _17643_ (.A1(net4972),
    .A2(_09105_),
    .B(net5946),
    .Y(_09468_));
 AO21x1_ASAP7_75t_R _17644_ (.A1(_09132_),
    .A2(_09396_),
    .B(net5946),
    .Y(_09469_));
 AOI21x1_ASAP7_75t_R _17645_ (.A1(_09468_),
    .A2(_09469_),
    .B(net5925),
    .Y(_09470_));
 OAI21x1_ASAP7_75t_R _17646_ (.A1(_09467_),
    .A2(_09470_),
    .B(net6303),
    .Y(_09471_));
 AOI21x1_ASAP7_75t_R _17647_ (.A1(_09465_),
    .A2(_09471_),
    .B(net5943),
    .Y(_09472_));
 OAI21x1_ASAP7_75t_R _17648_ (.A1(_09459_),
    .A2(_09472_),
    .B(net5942),
    .Y(_09473_));
 NAND2x1_ASAP7_75t_R _17649_ (.A(_09447_),
    .B(_09473_),
    .Y(_00013_));
 AO22x1_ASAP7_75t_R _17650_ (.A1(_09036_),
    .A2(_09243_),
    .B1(_09361_),
    .B2(net5551),
    .Y(_09474_));
 NOR2x1_ASAP7_75t_R _17651_ (.A(net5927),
    .B(_09323_),
    .Y(_09475_));
 AO21x1_ASAP7_75t_R _17652_ (.A1(_09475_),
    .A2(_09318_),
    .B(net5943),
    .Y(_09476_));
 AO21x1_ASAP7_75t_R _17653_ (.A1(net5927),
    .A2(_09474_),
    .B(_09476_),
    .Y(_09477_));
 AOI21x1_ASAP7_75t_R _17654_ (.A1(net5553),
    .A2(_09396_),
    .B(net6307),
    .Y(_09478_));
 AO21x1_ASAP7_75t_R _17655_ (.A1(net6309),
    .A2(net6307),
    .B(_09478_),
    .Y(_09479_));
 NOR2x1_ASAP7_75t_R _17656_ (.A(_09241_),
    .B(net5951),
    .Y(_09480_));
 OAI21x1_ASAP7_75t_R _17657_ (.A1(_09480_),
    .A2(_09342_),
    .B(_09309_),
    .Y(_09481_));
 AO21x1_ASAP7_75t_R _17658_ (.A1(_09481_),
    .A2(net6304),
    .B(net5554),
    .Y(_09482_));
 AO21x1_ASAP7_75t_R _17659_ (.A1(net5925),
    .A2(_09479_),
    .B(_09482_),
    .Y(_09483_));
 AOI21x1_ASAP7_75t_R _17660_ (.A1(_09477_),
    .A2(_09483_),
    .B(net5550),
    .Y(_09484_));
 AOI221x1_ASAP7_75t_R _17661_ (.A1(_01010_),
    .A2(net5947),
    .B1(net5552),
    .B2(net4713),
    .C(net6304),
    .Y(_09485_));
 OA21x2_ASAP7_75t_R _17662_ (.A1(net5922),
    .A2(net5948),
    .B(net6304),
    .Y(_09486_));
 AO21x1_ASAP7_75t_R _17663_ (.A1(net4598),
    .A2(_09259_),
    .B(net6306),
    .Y(_09487_));
 AO21x1_ASAP7_75t_R _17664_ (.A1(_09486_),
    .A2(_09487_),
    .B(net5943),
    .Y(_09488_));
 OAI21x1_ASAP7_75t_R _17665_ (.A1(_09485_),
    .A2(_09488_),
    .B(net5550),
    .Y(_09489_));
 AND3x1_ASAP7_75t_R _17666_ (.A(net5553),
    .B(net6306),
    .C(net4977),
    .Y(_09490_));
 AOI21x1_ASAP7_75t_R _17667_ (.A1(net5556),
    .A2(_09369_),
    .B(net6305),
    .Y(_09491_));
 OA21x2_ASAP7_75t_R _17668_ (.A1(_09490_),
    .A2(_09491_),
    .B(net5929),
    .Y(_09492_));
 AOI211x1_ASAP7_75t_R _17669_ (.A1(_09382_),
    .A2(net5922),
    .B(_09491_),
    .C(net5929),
    .Y(_09493_));
 NOR3x1_ASAP7_75t_R _17670_ (.A(_09492_),
    .B(net5554),
    .C(_09493_),
    .Y(_09494_));
 OAI21x1_ASAP7_75t_R _17671_ (.A1(_09489_),
    .A2(_09494_),
    .B(net6303),
    .Y(_09495_));
 NAND2x1_ASAP7_75t_R _17672_ (.A(_09082_),
    .B(_09083_),
    .Y(_09496_));
 NAND2x1_ASAP7_75t_R _17673_ (.A(_09210_),
    .B(_09496_),
    .Y(_09497_));
 OA21x2_ASAP7_75t_R _17674_ (.A1(net5947),
    .A2(_09036_),
    .B(net5927),
    .Y(_09498_));
 NAND2x1_ASAP7_75t_R _17675_ (.A(_09498_),
    .B(_09456_),
    .Y(_09499_));
 AOI21x1_ASAP7_75t_R _17676_ (.A1(_09497_),
    .A2(_09499_),
    .B(net5554),
    .Y(_09500_));
 AO21x1_ASAP7_75t_R _17677_ (.A1(net6308),
    .A2(_09045_),
    .B(net5946),
    .Y(_09501_));
 AOI21x1_ASAP7_75t_R _17678_ (.A1(_09501_),
    .A2(_09418_),
    .B(net5930),
    .Y(_09502_));
 AO21x1_ASAP7_75t_R _17679_ (.A1(_09089_),
    .A2(_09264_),
    .B(net6305),
    .Y(_09503_));
 AO21x1_ASAP7_75t_R _17680_ (.A1(_09503_),
    .A2(_09043_),
    .B(net5943),
    .Y(_09504_));
 NOR2x1_ASAP7_75t_R _17681_ (.A(_09502_),
    .B(_09504_),
    .Y(_09505_));
 OAI21x1_ASAP7_75t_R _17682_ (.A1(_09500_),
    .A2(_09505_),
    .B(net5550),
    .Y(_09506_));
 AO21x1_ASAP7_75t_R _17683_ (.A1(_09133_),
    .A2(net5923),
    .B(net6306),
    .Y(_09507_));
 AOI21x1_ASAP7_75t_R _17684_ (.A1(_09107_),
    .A2(_09507_),
    .B(net5943),
    .Y(_09508_));
 AOI21x1_ASAP7_75t_R _17685_ (.A1(net5025),
    .A2(net5555),
    .B(net6304),
    .Y(_09509_));
 AO21x1_ASAP7_75t_R _17686_ (.A1(_09132_),
    .A2(_09133_),
    .B(net6306),
    .Y(_09510_));
 NAND2x1_ASAP7_75t_R _17687_ (.A(_09509_),
    .B(_09510_),
    .Y(_09511_));
 AOI21x1_ASAP7_75t_R _17688_ (.A1(_09508_),
    .A2(_09511_),
    .B(net5550),
    .Y(_09512_));
 AO21x1_ASAP7_75t_R _17689_ (.A1(_09095_),
    .A2(_09040_),
    .B(net6305),
    .Y(_09513_));
 NAND2x1_ASAP7_75t_R _17690_ (.A(net5236),
    .B(net4713),
    .Y(_09514_));
 NAND3x1_ASAP7_75t_R _17691_ (.A(_09513_),
    .B(_09514_),
    .C(net5927),
    .Y(_09515_));
 NAND2x1_ASAP7_75t_R _17692_ (.A(net5025),
    .B(net5555),
    .Y(_09516_));
 AOI21x1_ASAP7_75t_R _17693_ (.A1(_09516_),
    .A2(_09343_),
    .B(net5554),
    .Y(_09517_));
 NAND2x1_ASAP7_75t_R _17694_ (.A(_09515_),
    .B(_09517_),
    .Y(_09518_));
 AOI21x1_ASAP7_75t_R _17695_ (.A1(_09512_),
    .A2(_09518_),
    .B(net6303),
    .Y(_09519_));
 NAND2x1_ASAP7_75t_R _17696_ (.A(_09506_),
    .B(_09519_),
    .Y(_09520_));
 OAI21x1_ASAP7_75t_R _17697_ (.A1(_09484_),
    .A2(_09495_),
    .B(_09520_),
    .Y(_00014_));
 AOI21x1_ASAP7_75t_R _17698_ (.A1(net6306),
    .A2(_09222_),
    .B(_09223_),
    .Y(_09521_));
 NOR2x1_ASAP7_75t_R _17699_ (.A(net5241),
    .B(net6306),
    .Y(_09522_));
 AOI21x1_ASAP7_75t_R _17700_ (.A1(net6306),
    .A2(_09283_),
    .B(_09522_),
    .Y(_09523_));
 AO21x1_ASAP7_75t_R _17701_ (.A1(_09523_),
    .A2(net5930),
    .B(net5924),
    .Y(_09524_));
 AOI21x1_ASAP7_75t_R _17702_ (.A1(net4530),
    .A2(_09521_),
    .B(_09524_),
    .Y(_09525_));
 OA21x2_ASAP7_75t_R _17703_ (.A1(_01016_),
    .A2(net6306),
    .B(net5930),
    .Y(_09526_));
 AO21x1_ASAP7_75t_R _17704_ (.A1(_09256_),
    .A2(net4787),
    .B(net5948),
    .Y(_09527_));
 AO21x1_ASAP7_75t_R _17705_ (.A1(_09526_),
    .A2(_09527_),
    .B(net6303),
    .Y(_09528_));
 AO21x1_ASAP7_75t_R _17706_ (.A1(net4598),
    .A2(net5025),
    .B(net6306),
    .Y(_09529_));
 AND3x1_ASAP7_75t_R _17707_ (.A(_09486_),
    .B(_09302_),
    .C(_09529_),
    .Y(_09530_));
 OAI21x1_ASAP7_75t_R _17708_ (.A1(_09528_),
    .A2(_09530_),
    .B(net5554),
    .Y(_09531_));
 NOR2x1_ASAP7_75t_R _17709_ (.A(_09525_),
    .B(_09531_),
    .Y(_09532_));
 AO21x1_ASAP7_75t_R _17710_ (.A1(_09188_),
    .A2(_09040_),
    .B(_08968_),
    .Y(_09533_));
 OAI21x1_ASAP7_75t_R _17711_ (.A1(net4788),
    .A2(net5238),
    .B(net5948),
    .Y(_09534_));
 AO21x1_ASAP7_75t_R _17712_ (.A1(_09533_),
    .A2(_09534_),
    .B(net6304),
    .Y(_09535_));
 AND3x1_ASAP7_75t_R _17713_ (.A(_09279_),
    .B(net6306),
    .C(_09174_),
    .Y(_09536_));
 OAI21x1_ASAP7_75t_R _17714_ (.A1(net4712),
    .A2(_09536_),
    .B(net6304),
    .Y(_09537_));
 AOI21x1_ASAP7_75t_R _17715_ (.A1(_09535_),
    .A2(_09537_),
    .B(net5924),
    .Y(_09538_));
 AO21x1_ASAP7_75t_R _17716_ (.A1(_09263_),
    .A2(net6305),
    .B(net5925),
    .Y(_09539_));
 OAI21x1_ASAP7_75t_R _17717_ (.A1(_09478_),
    .A2(_09539_),
    .B(net5924),
    .Y(_09540_));
 AO21x1_ASAP7_75t_R _17718_ (.A1(net5946),
    .A2(_09206_),
    .B(_09243_),
    .Y(_09541_));
 AOI21x1_ASAP7_75t_R _17719_ (.A1(net4974),
    .A2(_09541_),
    .B(net6304),
    .Y(_09542_));
 OAI21x1_ASAP7_75t_R _17720_ (.A1(_09540_),
    .A2(_09542_),
    .B(net5943),
    .Y(_09543_));
 OAI21x1_ASAP7_75t_R _17721_ (.A1(_09538_),
    .A2(_09543_),
    .B(net5942),
    .Y(_09544_));
 OAI21x1_ASAP7_75t_R _17722_ (.A1(net4596),
    .A2(_09214_),
    .B(net6304),
    .Y(_09545_));
 AO21x1_ASAP7_75t_R _17723_ (.A1(_09305_),
    .A2(_09514_),
    .B(net6304),
    .Y(_09546_));
 AOI21x1_ASAP7_75t_R _17724_ (.A1(_09545_),
    .A2(_09546_),
    .B(net6303),
    .Y(_09547_));
 NAND2x1_ASAP7_75t_R _17725_ (.A(net5930),
    .B(_09381_),
    .Y(_09548_));
 INVx1_ASAP7_75t_R _17726_ (.A(_09418_),
    .Y(_09549_));
 OAI21x1_ASAP7_75t_R _17727_ (.A1(_09548_),
    .A2(_09549_),
    .B(net6303),
    .Y(_09550_));
 AO21x1_ASAP7_75t_R _17728_ (.A1(_09286_),
    .A2(_09135_),
    .B(net5928),
    .Y(_09551_));
 AND3x1_ASAP7_75t_R _17729_ (.A(_09132_),
    .B(net6305),
    .C(_09089_),
    .Y(_09552_));
 NOR2x1_ASAP7_75t_R _17730_ (.A(_09551_),
    .B(_09552_),
    .Y(_09553_));
 OAI21x1_ASAP7_75t_R _17731_ (.A1(_09550_),
    .A2(_09553_),
    .B(net5943),
    .Y(_09554_));
 OAI21x1_ASAP7_75t_R _17732_ (.A1(_09547_),
    .A2(_09554_),
    .B(net5550),
    .Y(_09555_));
 AO21x1_ASAP7_75t_R _17733_ (.A1(net6311),
    .A2(net6307),
    .B(net5925),
    .Y(_09556_));
 NOR2x1_ASAP7_75t_R _17734_ (.A(_09222_),
    .B(_09117_),
    .Y(_09557_));
 OA21x2_ASAP7_75t_R _17735_ (.A1(_09556_),
    .A2(_09557_),
    .B(net6303),
    .Y(_09558_));
 AO21x1_ASAP7_75t_R _17736_ (.A1(_09279_),
    .A2(_09040_),
    .B(net5948),
    .Y(_09559_));
 NAND2x1_ASAP7_75t_R _17737_ (.A(_09559_),
    .B(_09297_),
    .Y(_09560_));
 OAI21x1_ASAP7_75t_R _17738_ (.A1(net6305),
    .A2(net4972),
    .B(_09455_),
    .Y(_09561_));
 AOI21x1_ASAP7_75t_R _17739_ (.A1(_09040_),
    .A2(net4597),
    .B(net5948),
    .Y(_09562_));
 OAI21x1_ASAP7_75t_R _17740_ (.A1(_09562_),
    .A2(net4714),
    .B(net6304),
    .Y(_09563_));
 AOI21x1_ASAP7_75t_R _17741_ (.A1(_09561_),
    .A2(_09563_),
    .B(net6303),
    .Y(_09564_));
 AOI211x1_ASAP7_75t_R _17742_ (.A1(_09558_),
    .A2(_09560_),
    .B(_09564_),
    .C(net5943),
    .Y(_09565_));
 OAI22x1_ASAP7_75t_R _17743_ (.A1(_09532_),
    .A2(_09544_),
    .B1(_09555_),
    .B2(_09565_),
    .Y(_00015_));
 AOI21x1_ASAP7_75t_R _17747_ (.A1(net129),
    .A2(_08907_),
    .B(_08910_),
    .Y(_09567_));
 NOR2x1_ASAP7_75t_R _17749_ (.A(net6321),
    .B(net6323),
    .Y(_09568_));
 INVx1_ASAP7_75t_R _17750_ (.A(_09568_),
    .Y(_09569_));
 NOR2x1_ASAP7_75t_R _17752_ (.A(net5569),
    .B(net5964),
    .Y(_09571_));
 NOR2x1_ASAP7_75t_R _17753_ (.A(net5960),
    .B(_09571_),
    .Y(_09572_));
 NOR2x1_ASAP7_75t_R _17754_ (.A(net5963),
    .B(net6296),
    .Y(_09573_));
 INVx1_ASAP7_75t_R _17755_ (.A(_09573_),
    .Y(_09574_));
 NAND2x1_ASAP7_75t_R _17758_ (.A(_01021_),
    .B(net5964),
    .Y(_09577_));
 AND3x1_ASAP7_75t_R _17759_ (.A(_09574_),
    .B(net5959),
    .C(net5548),
    .Y(_09578_));
 AOI21x1_ASAP7_75t_R _17760_ (.A1(_09569_),
    .A2(_09572_),
    .B(_09578_),
    .Y(_09579_));
 NAND2x1_ASAP7_75t_R _17761_ (.A(net6322),
    .B(net6323),
    .Y(_09580_));
 NAND2x1_ASAP7_75t_R _17764_ (.A(net5312),
    .B(net5963),
    .Y(_09583_));
 AND3x1_ASAP7_75t_R _17765_ (.A(net5921),
    .B(net6319),
    .C(_09583_),
    .Y(_09584_));
 NOR2x1_ASAP7_75t_R _17766_ (.A(_01019_),
    .B(net6321),
    .Y(_09585_));
 AO21x1_ASAP7_75t_R _17768_ (.A1(net6324),
    .A2(net6321),
    .B(net6320),
    .Y(_09587_));
 INVx1_ASAP7_75t_R _17769_ (.A(_00960_),
    .Y(_09588_));
 XOR2x2_ASAP7_75t_R _17770_ (.A(_08829_),
    .B(_09588_),
    .Y(_09589_));
 INVx1_ASAP7_75t_R _17771_ (.A(_08932_),
    .Y(_09590_));
 OAI21x1_ASAP7_75t_R _17772_ (.A1(net6683),
    .A2(_09589_),
    .B(_09590_),
    .Y(_09591_));
 OAI21x1_ASAP7_75t_R _17774_ (.A1(_09585_),
    .A2(_09587_),
    .B(net6293),
    .Y(_09593_));
 INVx1_ASAP7_75t_R _17775_ (.A(_08936_),
    .Y(_09594_));
 OAI21x1_ASAP7_75t_R _17777_ (.A1(_09584_),
    .A2(_09593_),
    .B(net5919),
    .Y(_09596_));
 AOI21x1_ASAP7_75t_R _17778_ (.A1(net6315),
    .A2(_09579_),
    .B(_09596_),
    .Y(_09597_));
 INVx1_ASAP7_75t_R _17779_ (.A(_08944_),
    .Y(_09598_));
 INVx1_ASAP7_75t_R _17782_ (.A(_01021_),
    .Y(_09601_));
 AO21x1_ASAP7_75t_R _17783_ (.A1(net6368),
    .A2(net6466),
    .B(_09601_),
    .Y(_09602_));
 INVx1_ASAP7_75t_R _17784_ (.A(net5563),
    .Y(_09603_));
 NOR2x2_ASAP7_75t_R _17785_ (.A(_09603_),
    .B(net6321),
    .Y(_09604_));
 NOR2x2_ASAP7_75t_R _17786_ (.A(_09604_),
    .B(net6320),
    .Y(_09605_));
 NAND2x1_ASAP7_75t_R _17787_ (.A(net5234),
    .B(_09605_),
    .Y(_09606_));
 NAND2x1_ASAP7_75t_R _17788_ (.A(_08923_),
    .B(net6296),
    .Y(_09607_));
 INVx1_ASAP7_75t_R _17789_ (.A(_01023_),
    .Y(_09608_));
 AO21x1_ASAP7_75t_R _17790_ (.A1(net6368),
    .A2(net6466),
    .B(_09608_),
    .Y(_09609_));
 AO21x1_ASAP7_75t_R _17792_ (.A1(net5547),
    .A2(net5233),
    .B(net5959),
    .Y(_09611_));
 AOI21x1_ASAP7_75t_R _17793_ (.A1(_09606_),
    .A2(_09611_),
    .B(net6295),
    .Y(_09612_));
 AO21x1_ASAP7_75t_R _17795_ (.A1(net5963),
    .A2(net5568),
    .B(net6320),
    .Y(_09614_));
 OAI21x1_ASAP7_75t_R _17796_ (.A1(net5963),
    .A2(net6296),
    .B(net6320),
    .Y(_09615_));
 OA21x2_ASAP7_75t_R _17797_ (.A1(_09614_),
    .A2(_09571_),
    .B(_09615_),
    .Y(_09616_));
 NOR2x1_ASAP7_75t_R _17798_ (.A(net6315),
    .B(_09616_),
    .Y(_09617_));
 OAI21x1_ASAP7_75t_R _17800_ (.A1(_09612_),
    .A2(_09617_),
    .B(net6313),
    .Y(_09619_));
 NAND2x1_ASAP7_75t_R _17801_ (.A(_09598_),
    .B(_09619_),
    .Y(_09620_));
 AO21x1_ASAP7_75t_R _17802_ (.A1(net6368),
    .A2(net6466),
    .B(_01024_),
    .Y(_09621_));
 NOR2x1_ASAP7_75t_R _17803_ (.A(net5956),
    .B(net5545),
    .Y(_09622_));
 NOR2x1_ASAP7_75t_R _17805_ (.A(net6295),
    .B(_09605_),
    .Y(_09624_));
 NOR2x1_ASAP7_75t_R _17806_ (.A(net5314),
    .B(net6321),
    .Y(_09625_));
 INVx1_ASAP7_75t_R _17807_ (.A(_09625_),
    .Y(_09626_));
 AO21x1_ASAP7_75t_R _17809_ (.A1(_09626_),
    .A2(_09621_),
    .B(net5957),
    .Y(_09628_));
 AOI21x1_ASAP7_75t_R _17810_ (.A1(_09624_),
    .A2(_09628_),
    .B(net6312),
    .Y(_09629_));
 OAI21x1_ASAP7_75t_R _17811_ (.A1(_09622_),
    .A2(_09593_),
    .B(_09629_),
    .Y(_09630_));
 AO21x1_ASAP7_75t_R _17812_ (.A1(net6368),
    .A2(net6466),
    .B(net5563),
    .Y(_09631_));
 NAND2x1_ASAP7_75t_R _17814_ (.A(net5963),
    .B(net6323),
    .Y(_09633_));
 AOI21x1_ASAP7_75t_R _17815_ (.A1(net5267),
    .A2(_09633_),
    .B(net5960),
    .Y(_09634_));
 INVx1_ASAP7_75t_R _17816_ (.A(_01026_),
    .Y(_09635_));
 AO21x1_ASAP7_75t_R _17817_ (.A1(net6368),
    .A2(net6466),
    .B(_09635_),
    .Y(_09636_));
 INVx1_ASAP7_75t_R _17818_ (.A(_09636_),
    .Y(_09637_));
 AO21x1_ASAP7_75t_R _17819_ (.A1(net6296),
    .A2(net5963),
    .B(net6320),
    .Y(_09638_));
 NOR2x1_ASAP7_75t_R _17820_ (.A(_09637_),
    .B(_09638_),
    .Y(_09639_));
 OAI21x1_ASAP7_75t_R _17823_ (.A1(_09634_),
    .A2(_09639_),
    .B(net6295),
    .Y(_09642_));
 NOR2x1_ASAP7_75t_R _17824_ (.A(_01029_),
    .B(net6321),
    .Y(_09643_));
 INVx1_ASAP7_75t_R _17825_ (.A(_09643_),
    .Y(_09644_));
 INVx1_ASAP7_75t_R _17826_ (.A(_01028_),
    .Y(_09645_));
 AO21x1_ASAP7_75t_R _17827_ (.A1(net6368),
    .A2(net6466),
    .B(_09645_),
    .Y(_09646_));
 AO21x1_ASAP7_75t_R _17829_ (.A1(_09644_),
    .A2(_09646_),
    .B(net5955),
    .Y(_09648_));
 AND2x2_ASAP7_75t_R _17831_ (.A(_09614_),
    .B(net6315),
    .Y(_09650_));
 AOI21x1_ASAP7_75t_R _17832_ (.A1(_09648_),
    .A2(_09650_),
    .B(net5920),
    .Y(_09651_));
 AOI21x1_ASAP7_75t_R _17833_ (.A1(_09642_),
    .A2(_09651_),
    .B(_09598_),
    .Y(_09652_));
 INVx1_ASAP7_75t_R _17834_ (.A(_08940_),
    .Y(_09653_));
 AOI21x1_ASAP7_75t_R _17836_ (.A1(_09630_),
    .A2(_09652_),
    .B(_09653_),
    .Y(_09655_));
 OAI21x1_ASAP7_75t_R _17837_ (.A1(_09597_),
    .A2(_09620_),
    .B(_09655_),
    .Y(_09656_));
 AOI21x1_ASAP7_75t_R _17838_ (.A1(net5964),
    .A2(net6296),
    .B(_08929_),
    .Y(_09657_));
 NAND2x1_ASAP7_75t_R _17839_ (.A(net6324),
    .B(net5965),
    .Y(_09658_));
 NAND2x1_ASAP7_75t_R _17840_ (.A(_09657_),
    .B(_09658_),
    .Y(_09659_));
 AO21x1_ASAP7_75t_R _17843_ (.A1(_09658_),
    .A2(net5547),
    .B(net6320),
    .Y(_09662_));
 AOI21x1_ASAP7_75t_R _17844_ (.A1(_09659_),
    .A2(_09662_),
    .B(net6295),
    .Y(_09663_));
 NAND2x1_ASAP7_75t_R _17845_ (.A(net5315),
    .B(net5964),
    .Y(_09664_));
 AO21x1_ASAP7_75t_R _17846_ (.A1(_09664_),
    .A2(_09646_),
    .B(net6320),
    .Y(_09665_));
 NOR2x1_ASAP7_75t_R _17847_ (.A(net5563),
    .B(net6321),
    .Y(_09666_));
 INVx1_ASAP7_75t_R _17848_ (.A(_09666_),
    .Y(_09667_));
 INVx1_ASAP7_75t_R _17849_ (.A(_01019_),
    .Y(_09668_));
 AO21x1_ASAP7_75t_R _17850_ (.A1(net6368),
    .A2(net6466),
    .B(_09668_),
    .Y(_09669_));
 AO21x1_ASAP7_75t_R _17852_ (.A1(_09667_),
    .A2(_09669_),
    .B(net5957),
    .Y(_09671_));
 AOI21x1_ASAP7_75t_R _17853_ (.A1(_09665_),
    .A2(_09671_),
    .B(net6318),
    .Y(_09672_));
 OA21x2_ASAP7_75t_R _17854_ (.A1(_09663_),
    .A2(_09672_),
    .B(net6312),
    .Y(_09673_));
 NAND2x1_ASAP7_75t_R _17855_ (.A(net5313),
    .B(net5964),
    .Y(_09674_));
 OA21x2_ASAP7_75t_R _17856_ (.A1(_09674_),
    .A2(net5955),
    .B(net6295),
    .Y(_09675_));
 AO21x1_ASAP7_75t_R _17857_ (.A1(net6368),
    .A2(net6466),
    .B(net5313),
    .Y(_09676_));
 AOI22x1_ASAP7_75t_R _17859_ (.A1(net4784),
    .A2(_09676_),
    .B1(net6320),
    .B2(_09637_),
    .Y(_09678_));
 NAND2x1_ASAP7_75t_R _17860_ (.A(_09675_),
    .B(_09678_),
    .Y(_09679_));
 AO21x1_ASAP7_75t_R _17861_ (.A1(net6368),
    .A2(net6466),
    .B(_09603_),
    .Y(_09680_));
 OA21x2_ASAP7_75t_R _17862_ (.A1(net6320),
    .A2(_09680_),
    .B(net6318),
    .Y(_09681_));
 AO21x1_ASAP7_75t_R _17863_ (.A1(_09580_),
    .A2(_09667_),
    .B(net5957),
    .Y(_09682_));
 AOI21x1_ASAP7_75t_R _17864_ (.A1(_09681_),
    .A2(_09682_),
    .B(net6312),
    .Y(_09683_));
 AO21x1_ASAP7_75t_R _17865_ (.A1(_09679_),
    .A2(_09683_),
    .B(net5953),
    .Y(_09684_));
 NOR2x1_ASAP7_75t_R _17866_ (.A(_09608_),
    .B(net6321),
    .Y(_09685_));
 INVx1_ASAP7_75t_R _17867_ (.A(_09685_),
    .Y(_09686_));
 AO21x1_ASAP7_75t_R _17868_ (.A1(_09574_),
    .A2(_09686_),
    .B(net5955),
    .Y(_09687_));
 NAND2x1_ASAP7_75t_R _17869_ (.A(_08922_),
    .B(net6296),
    .Y(_09688_));
 NAND2x1_ASAP7_75t_R _17870_ (.A(_09674_),
    .B(_09688_),
    .Y(_09689_));
 AOI21x1_ASAP7_75t_R _17871_ (.A1(net5956),
    .A2(_09689_),
    .B(net6317),
    .Y(_09690_));
 NAND2x1_ASAP7_75t_R _17872_ (.A(_09687_),
    .B(_09690_),
    .Y(_09691_));
 INVx2_ASAP7_75t_R _17873_ (.A(_09631_),
    .Y(_09692_));
 NOR2x1_ASAP7_75t_R _17874_ (.A(_01036_),
    .B(net6320),
    .Y(_09693_));
 AO21x1_ASAP7_75t_R _17875_ (.A1(_09692_),
    .A2(net6320),
    .B(_09693_),
    .Y(_09694_));
 OA21x2_ASAP7_75t_R _17877_ (.A1(_09694_),
    .A2(net6295),
    .B(net5920),
    .Y(_09696_));
 AOI21x1_ASAP7_75t_R _17878_ (.A1(_09691_),
    .A2(_09696_),
    .B(_09598_),
    .Y(_09697_));
 OA21x2_ASAP7_75t_R _17879_ (.A1(net5957),
    .A2(_09636_),
    .B(net6318),
    .Y(_09698_));
 NAND2x1_ASAP7_75t_R _17880_ (.A(net5958),
    .B(net5231),
    .Y(_09699_));
 OA21x2_ASAP7_75t_R _17881_ (.A1(net5958),
    .A2(net4968),
    .B(_09699_),
    .Y(_09700_));
 NAND2x1_ASAP7_75t_R _17882_ (.A(_09698_),
    .B(_09700_),
    .Y(_09701_));
 NAND2x1_ASAP7_75t_R _17883_ (.A(net6320),
    .B(net5231),
    .Y(_09702_));
 AO21x1_ASAP7_75t_R _17884_ (.A1(net5964),
    .A2(net5546),
    .B(net6320),
    .Y(_09703_));
 INVx1_ASAP7_75t_R _17885_ (.A(_01027_),
    .Y(_09704_));
 AO21x1_ASAP7_75t_R _17886_ (.A1(net6368),
    .A2(net6466),
    .B(_09704_),
    .Y(_09705_));
 INVx1_ASAP7_75t_R _17887_ (.A(_09705_),
    .Y(_09706_));
 OA21x2_ASAP7_75t_R _17888_ (.A1(_09703_),
    .A2(_09706_),
    .B(net6293),
    .Y(_09707_));
 AOI21x1_ASAP7_75t_R _17889_ (.A1(_09702_),
    .A2(_09707_),
    .B(net5920),
    .Y(_09708_));
 NAND2x1_ASAP7_75t_R _17890_ (.A(_09701_),
    .B(_09708_),
    .Y(_09709_));
 AOI21x1_ASAP7_75t_R _17891_ (.A1(_09697_),
    .A2(_09709_),
    .B(net5954),
    .Y(_09710_));
 OAI21x1_ASAP7_75t_R _17892_ (.A1(_09673_),
    .A2(_09684_),
    .B(_09710_),
    .Y(_09711_));
 NAND2x1_ASAP7_75t_R _17893_ (.A(_09656_),
    .B(_09711_),
    .Y(_00016_));
 INVx1_ASAP7_75t_R _17894_ (.A(net5544),
    .Y(_09712_));
 OA21x2_ASAP7_75t_R _17895_ (.A1(_09712_),
    .A2(net5023),
    .B(net5955),
    .Y(_09713_));
 AOI211x1_ASAP7_75t_R _17897_ (.A1(net6319),
    .A2(_09689_),
    .B(_09713_),
    .C(net6295),
    .Y(_09715_));
 NOR2x1_ASAP7_75t_R _17898_ (.A(net5958),
    .B(_09692_),
    .Y(_09716_));
 NAND2x1_ASAP7_75t_R _17899_ (.A(net5964),
    .B(net6324),
    .Y(_09717_));
 AND2x2_ASAP7_75t_R _17900_ (.A(_09716_),
    .B(_09717_),
    .Y(_09718_));
 NOR2x1_ASAP7_75t_R _17901_ (.A(net6323),
    .B(net6325),
    .Y(_09719_));
 OAI21x1_ASAP7_75t_R _17902_ (.A1(_09719_),
    .A2(_09587_),
    .B(net6293),
    .Y(_09720_));
 OAI21x1_ASAP7_75t_R _17903_ (.A1(_09718_),
    .A2(_09720_),
    .B(net5920),
    .Y(_09721_));
 NOR2x1_ASAP7_75t_R _17904_ (.A(_09715_),
    .B(_09721_),
    .Y(_09722_));
 AO21x1_ASAP7_75t_R _17905_ (.A1(net6321),
    .A2(_09668_),
    .B(net6320),
    .Y(_09723_));
 NOR2x1_ASAP7_75t_R _17906_ (.A(net5266),
    .B(net5229),
    .Y(_09724_));
 NOR2x1_ASAP7_75t_R _17907_ (.A(net5568),
    .B(net5961),
    .Y(_09725_));
 AO21x1_ASAP7_75t_R _17909_ (.A1(_09725_),
    .A2(net5963),
    .B(net6314),
    .Y(_09727_));
 OAI21x1_ASAP7_75t_R _17910_ (.A1(_09724_),
    .A2(_09727_),
    .B(net6313),
    .Y(_09728_));
 NAND2x1_ASAP7_75t_R _17911_ (.A(_01019_),
    .B(net5963),
    .Y(_09729_));
 INVx1_ASAP7_75t_R _17912_ (.A(_09602_),
    .Y(_09730_));
 NOR2x1_ASAP7_75t_R _17913_ (.A(net6320),
    .B(_09730_),
    .Y(_09731_));
 AOI21x1_ASAP7_75t_R _17914_ (.A1(_09569_),
    .A2(_09731_),
    .B(net6295),
    .Y(_09732_));
 OA21x2_ASAP7_75t_R _17915_ (.A1(net5960),
    .A2(_09729_),
    .B(_09732_),
    .Y(_09733_));
 OAI21x1_ASAP7_75t_R _17916_ (.A1(_09728_),
    .A2(_09733_),
    .B(net5953),
    .Y(_09734_));
 OAI21x1_ASAP7_75t_R _17917_ (.A1(_09722_),
    .A2(_09734_),
    .B(net5954),
    .Y(_09735_));
 AND2x2_ASAP7_75t_R _17918_ (.A(_09657_),
    .B(_09676_),
    .Y(_09736_));
 NAND2x1_ASAP7_75t_R _17919_ (.A(net6322),
    .B(net5965),
    .Y(_09737_));
 INVx1_ASAP7_75t_R _17920_ (.A(_09737_),
    .Y(_09738_));
 NOR2x1_ASAP7_75t_R _17921_ (.A(_09614_),
    .B(_09738_),
    .Y(_09739_));
 OAI21x1_ASAP7_75t_R _17922_ (.A1(_09736_),
    .A2(_09739_),
    .B(net6295),
    .Y(_09740_));
 AO21x1_ASAP7_75t_R _17923_ (.A1(net5918),
    .A2(_09644_),
    .B(net5955),
    .Y(_09741_));
 AO21x1_ASAP7_75t_R _17924_ (.A1(_09674_),
    .A2(net5267),
    .B(net6319),
    .Y(_09742_));
 AO21x1_ASAP7_75t_R _17925_ (.A1(_09741_),
    .A2(_09742_),
    .B(net6295),
    .Y(_09743_));
 AOI21x1_ASAP7_75t_R _17927_ (.A1(_09740_),
    .A2(_09743_),
    .B(net5919),
    .Y(_09745_));
 AOI21x1_ASAP7_75t_R _17928_ (.A1(net5312),
    .A2(net6322),
    .B(net5962),
    .Y(_09746_));
 AOI211x1_ASAP7_75t_R _17929_ (.A1(_09746_),
    .A2(net5548),
    .B(_09724_),
    .C(net6295),
    .Y(_09747_));
 AO21x1_ASAP7_75t_R _17930_ (.A1(_09688_),
    .A2(_09729_),
    .B(net5959),
    .Y(_09748_));
 NOR2x1_ASAP7_75t_R _17931_ (.A(net6317),
    .B(_09605_),
    .Y(_09749_));
 AO21x1_ASAP7_75t_R _17932_ (.A1(_09748_),
    .A2(_09749_),
    .B(net6313),
    .Y(_09750_));
 OAI21x1_ASAP7_75t_R _17933_ (.A1(_09747_),
    .A2(_09750_),
    .B(_09598_),
    .Y(_09751_));
 NOR2x1_ASAP7_75t_R _17934_ (.A(_09745_),
    .B(_09751_),
    .Y(_09752_));
 INVx1_ASAP7_75t_R _17935_ (.A(_09688_),
    .Y(_09753_));
 AO21x1_ASAP7_75t_R _17936_ (.A1(net5963),
    .A2(net5568),
    .B(net5960),
    .Y(_09754_));
 NOR2x1_ASAP7_75t_R _17937_ (.A(_09753_),
    .B(_09754_),
    .Y(_09755_));
 AO21x1_ASAP7_75t_R _17938_ (.A1(net4785),
    .A2(_09574_),
    .B(net6295),
    .Y(_09756_));
 OA21x2_ASAP7_75t_R _17939_ (.A1(net6319),
    .A2(net5233),
    .B(net6295),
    .Y(_09757_));
 INVx1_ASAP7_75t_R _17940_ (.A(_09580_),
    .Y(_09758_));
 OAI21x1_ASAP7_75t_R _17941_ (.A1(_09758_),
    .A2(_09719_),
    .B(net6319),
    .Y(_09759_));
 AOI21x1_ASAP7_75t_R _17942_ (.A1(_09757_),
    .A2(_09759_),
    .B(net5919),
    .Y(_09760_));
 OA21x2_ASAP7_75t_R _17943_ (.A1(_09755_),
    .A2(_09756_),
    .B(_09760_),
    .Y(_09761_));
 AO21x1_ASAP7_75t_R _17944_ (.A1(_01031_),
    .A2(net5959),
    .B(net6295),
    .Y(_09762_));
 OA21x2_ASAP7_75t_R _17945_ (.A1(_09568_),
    .A2(_09712_),
    .B(net6320),
    .Y(_09763_));
 OAI21x1_ASAP7_75t_R _17946_ (.A1(_09762_),
    .A2(_09763_),
    .B(net5919),
    .Y(_09764_));
 AND3x1_ASAP7_75t_R _17947_ (.A(net5548),
    .B(net5959),
    .C(net5021),
    .Y(_09765_));
 NAND2x1_ASAP7_75t_R _17948_ (.A(_09621_),
    .B(_09686_),
    .Y(_09766_));
 AO21x1_ASAP7_75t_R _17949_ (.A1(_09766_),
    .A2(net6320),
    .B(net6317),
    .Y(_09767_));
 NOR2x1_ASAP7_75t_R _17950_ (.A(_09765_),
    .B(_09767_),
    .Y(_09768_));
 OAI21x1_ASAP7_75t_R _17951_ (.A1(_09764_),
    .A2(_09768_),
    .B(net5953),
    .Y(_09769_));
 OAI21x1_ASAP7_75t_R _17952_ (.A1(_09761_),
    .A2(_09769_),
    .B(net5542),
    .Y(_09770_));
 AO21x1_ASAP7_75t_R _17953_ (.A1(net5547),
    .A2(_09646_),
    .B(net5955),
    .Y(_09771_));
 AO21x1_ASAP7_75t_R _17954_ (.A1(net6321),
    .A2(net5546),
    .B(net6320),
    .Y(_09772_));
 NAND2x1_ASAP7_75t_R _17955_ (.A(net6318),
    .B(_08936_),
    .Y(_09773_));
 INVx1_ASAP7_75t_R _17956_ (.A(_09773_),
    .Y(_09774_));
 OA21x2_ASAP7_75t_R _17957_ (.A1(_09585_),
    .A2(_09772_),
    .B(_09774_),
    .Y(_09775_));
 NAND2x1_ASAP7_75t_R _17958_ (.A(_09771_),
    .B(_09775_),
    .Y(_09776_));
 NOR2x1_ASAP7_75t_R _17959_ (.A(net6295),
    .B(_09739_),
    .Y(_09777_));
 NAND2x1_ASAP7_75t_R _17960_ (.A(net5921),
    .B(_09657_),
    .Y(_09778_));
 AND2x2_ASAP7_75t_R _17961_ (.A(_09778_),
    .B(net5920),
    .Y(_09779_));
 AO21x1_ASAP7_75t_R _17962_ (.A1(_09729_),
    .A2(_09636_),
    .B(net5960),
    .Y(_09780_));
 NAND2x1_ASAP7_75t_R _17963_ (.A(_01037_),
    .B(net5961),
    .Y(_09781_));
 OA21x2_ASAP7_75t_R _17964_ (.A1(_09781_),
    .A2(net6313),
    .B(net6295),
    .Y(_09782_));
 AOI22x1_ASAP7_75t_R _17965_ (.A1(_09777_),
    .A2(_09779_),
    .B1(_09780_),
    .B2(_09782_),
    .Y(_09783_));
 AOI21x1_ASAP7_75t_R _17966_ (.A1(_09776_),
    .A2(_09783_),
    .B(net5953),
    .Y(_09784_));
 OAI22x1_ASAP7_75t_R _17967_ (.A1(_09735_),
    .A2(_09752_),
    .B1(_09770_),
    .B2(_09784_),
    .Y(_00017_));
 OA21x2_ASAP7_75t_R _17968_ (.A1(_01033_),
    .A2(_08929_),
    .B(net6318),
    .Y(_09785_));
 OAI21x1_ASAP7_75t_R _17969_ (.A1(net6321),
    .A2(net6323),
    .B(_09609_),
    .Y(_09786_));
 NAND2x1_ASAP7_75t_R _17970_ (.A(net5961),
    .B(_09786_),
    .Y(_09787_));
 AOI21x1_ASAP7_75t_R _17971_ (.A1(_09785_),
    .A2(_09787_),
    .B(net6312),
    .Y(_09788_));
 AOI21x1_ASAP7_75t_R _17972_ (.A1(_01035_),
    .A2(net5960),
    .B(_09572_),
    .Y(_09789_));
 NAND2x1_ASAP7_75t_R _17973_ (.A(net6294),
    .B(_09789_),
    .Y(_09790_));
 NAND2x1_ASAP7_75t_R _17974_ (.A(_09788_),
    .B(_09790_),
    .Y(_09791_));
 INVx1_ASAP7_75t_R _17975_ (.A(net5547),
    .Y(_09792_));
 OAI21x1_ASAP7_75t_R _17976_ (.A1(_09792_),
    .A2(net5229),
    .B(_09780_),
    .Y(_09793_));
 AO21x1_ASAP7_75t_R _17977_ (.A1(_09667_),
    .A2(net5544),
    .B(net6320),
    .Y(_09794_));
 AOI21x1_ASAP7_75t_R _17978_ (.A1(_09794_),
    .A2(_09675_),
    .B(net5920),
    .Y(_09795_));
 OAI21x1_ASAP7_75t_R _17979_ (.A1(net6295),
    .A2(_09793_),
    .B(_09795_),
    .Y(_09796_));
 AOI21x1_ASAP7_75t_R _17980_ (.A1(_09791_),
    .A2(_09796_),
    .B(net5954),
    .Y(_09797_));
 AND3x1_ASAP7_75t_R _17981_ (.A(_09664_),
    .B(net5957),
    .C(net5268),
    .Y(_09798_));
 AND3x1_ASAP7_75t_R _17983_ (.A(_09633_),
    .B(net6320),
    .C(_09646_),
    .Y(_09800_));
 OAI21x1_ASAP7_75t_R _17984_ (.A1(_09798_),
    .A2(_09800_),
    .B(net6316),
    .Y(_09801_));
 INVx1_ASAP7_75t_R _17985_ (.A(_01037_),
    .Y(_09802_));
 OAI21x1_ASAP7_75t_R _17986_ (.A1(net6325),
    .A2(net6323),
    .B(net5921),
    .Y(_09803_));
 AOI21x1_ASAP7_75t_R _17987_ (.A1(net5961),
    .A2(_09803_),
    .B(net6314),
    .Y(_09804_));
 OAI21x1_ASAP7_75t_R _17988_ (.A1(_09802_),
    .A2(net5961),
    .B(_09804_),
    .Y(_09805_));
 NAND2x1_ASAP7_75t_R _17989_ (.A(_09801_),
    .B(_09805_),
    .Y(_09806_));
 AO21x1_ASAP7_75t_R _17990_ (.A1(net5547),
    .A2(_01033_),
    .B(net6320),
    .Y(_09807_));
 INVx1_ASAP7_75t_R _17991_ (.A(_09807_),
    .Y(_09808_));
 AO21x1_ASAP7_75t_R _17992_ (.A1(_09633_),
    .A2(_09716_),
    .B(_09773_),
    .Y(_09809_));
 AO21x1_ASAP7_75t_R _17993_ (.A1(net4968),
    .A2(net5267),
    .B(net6320),
    .Y(_09810_));
 OR2x2_ASAP7_75t_R _17994_ (.A(_01036_),
    .B(_08929_),
    .Y(_09811_));
 INVx1_ASAP7_75t_R _17995_ (.A(_09811_),
    .Y(_09812_));
 NAND2x1_ASAP7_75t_R _17996_ (.A(_08936_),
    .B(_09591_),
    .Y(_09813_));
 NOR2x1_ASAP7_75t_R _17997_ (.A(_09812_),
    .B(_09813_),
    .Y(_09814_));
 AOI21x1_ASAP7_75t_R _17998_ (.A1(_09810_),
    .A2(_09814_),
    .B(_09653_),
    .Y(_09815_));
 OAI21x1_ASAP7_75t_R _17999_ (.A1(_09808_),
    .A2(_09809_),
    .B(_09815_),
    .Y(_09816_));
 AOI21x1_ASAP7_75t_R _18000_ (.A1(net5920),
    .A2(_09806_),
    .B(_09816_),
    .Y(_09817_));
 OAI21x1_ASAP7_75t_R _18001_ (.A1(_09797_),
    .A2(_09817_),
    .B(net5953),
    .Y(_09818_));
 INVx1_ASAP7_75t_R _18002_ (.A(net5568),
    .Y(_09819_));
 NAND2x1_ASAP7_75t_R _18003_ (.A(_09819_),
    .B(net5963),
    .Y(_09820_));
 AO21x1_ASAP7_75t_R _18004_ (.A1(net6368),
    .A2(net6466),
    .B(_01021_),
    .Y(_09821_));
 AO21x1_ASAP7_75t_R _18005_ (.A1(_09820_),
    .A2(_09821_),
    .B(net5960),
    .Y(_09822_));
 AOI21x1_ASAP7_75t_R _18006_ (.A1(_09787_),
    .A2(_09822_),
    .B(net6295),
    .Y(_09823_));
 AND2x2_ASAP7_75t_R _18007_ (.A(_09716_),
    .B(_09633_),
    .Y(_09824_));
 OAI21x1_ASAP7_75t_R _18008_ (.A1(net6320),
    .A2(_09766_),
    .B(net6295),
    .Y(_09825_));
 NOR2x1_ASAP7_75t_R _18009_ (.A(_09824_),
    .B(_09825_),
    .Y(_09826_));
 OAI21x1_ASAP7_75t_R _18010_ (.A1(_09823_),
    .A2(_09826_),
    .B(net5920),
    .Y(_09827_));
 INVx3_ASAP7_75t_R _18011_ (.A(_09604_),
    .Y(_09828_));
 AOI21x1_ASAP7_75t_R _18012_ (.A1(_09828_),
    .A2(_09580_),
    .B(_08929_),
    .Y(_09829_));
 AO21x1_ASAP7_75t_R _18013_ (.A1(net6368),
    .A2(net6466),
    .B(net5312),
    .Y(_09830_));
 AND3x1_ASAP7_75t_R _18014_ (.A(net5547),
    .B(net5962),
    .C(_09830_),
    .Y(_09831_));
 OAI21x1_ASAP7_75t_R _18015_ (.A1(_09829_),
    .A2(_09831_),
    .B(net6314),
    .Y(_09832_));
 INVx1_ASAP7_75t_R _18016_ (.A(_09723_),
    .Y(_09833_));
 AOI21x1_ASAP7_75t_R _18017_ (.A1(net5548),
    .A2(_09833_),
    .B(_09572_),
    .Y(_09834_));
 AOI21x1_ASAP7_75t_R _18018_ (.A1(net6294),
    .A2(_09834_),
    .B(net5920),
    .Y(_09835_));
 NAND2x1_ASAP7_75t_R _18019_ (.A(_09832_),
    .B(_09835_),
    .Y(_09836_));
 AOI21x1_ASAP7_75t_R _18020_ (.A1(_09827_),
    .A2(_09836_),
    .B(net5954),
    .Y(_09837_));
 OA21x2_ASAP7_75t_R _18021_ (.A1(net5963),
    .A2(_09819_),
    .B(net5960),
    .Y(_09838_));
 NAND2x1_ASAP7_75t_R _18022_ (.A(_09569_),
    .B(_09838_),
    .Y(_09839_));
 AOI21x1_ASAP7_75t_R _18023_ (.A1(_09628_),
    .A2(_09839_),
    .B(net6318),
    .Y(_09840_));
 AO21x1_ASAP7_75t_R _18024_ (.A1(_09626_),
    .A2(_09821_),
    .B(net5956),
    .Y(_09841_));
 AO21x1_ASAP7_75t_R _18025_ (.A1(net5547),
    .A2(_09621_),
    .B(net6320),
    .Y(_09842_));
 AOI21x1_ASAP7_75t_R _18026_ (.A1(_09841_),
    .A2(_09842_),
    .B(net6295),
    .Y(_09843_));
 OAI21x1_ASAP7_75t_R _18027_ (.A1(_09840_),
    .A2(_09843_),
    .B(net5920),
    .Y(_09844_));
 NAND2x1p5_ASAP7_75t_R _18028_ (.A(net5267),
    .B(net4784),
    .Y(_09845_));
 NOR2x1_ASAP7_75t_R _18029_ (.A(_08929_),
    .B(_09706_),
    .Y(_09846_));
 NAND2x1_ASAP7_75t_R _18030_ (.A(_09717_),
    .B(_09846_),
    .Y(_09847_));
 AOI21x1_ASAP7_75t_R _18031_ (.A1(_09845_),
    .A2(_09847_),
    .B(net6317),
    .Y(_09848_));
 AO21x1_ASAP7_75t_R _18032_ (.A1(net5965),
    .A2(net6322),
    .B(net6320),
    .Y(_09849_));
 AOI21x1_ASAP7_75t_R _18033_ (.A1(_09821_),
    .A2(_09657_),
    .B(net6295),
    .Y(_09850_));
 OA21x2_ASAP7_75t_R _18034_ (.A1(_09625_),
    .A2(_09849_),
    .B(_09850_),
    .Y(_09851_));
 OAI21x1_ASAP7_75t_R _18035_ (.A1(_09848_),
    .A2(_09851_),
    .B(net6312),
    .Y(_09852_));
 AOI21x1_ASAP7_75t_R _18036_ (.A1(_09844_),
    .A2(_09852_),
    .B(net5543),
    .Y(_09853_));
 OAI21x1_ASAP7_75t_R _18037_ (.A1(_09837_),
    .A2(_09853_),
    .B(_09598_),
    .Y(_09854_));
 NAND2x1_ASAP7_75t_R _18038_ (.A(_09818_),
    .B(_09854_),
    .Y(_00018_));
 AO21x1_ASAP7_75t_R _18039_ (.A1(_09580_),
    .A2(_09667_),
    .B(net6320),
    .Y(_09855_));
 AO21x1_ASAP7_75t_R _18040_ (.A1(_09658_),
    .A2(_09688_),
    .B(net5957),
    .Y(_09856_));
 AOI21x1_ASAP7_75t_R _18041_ (.A1(_09855_),
    .A2(_09856_),
    .B(net6318),
    .Y(_09857_));
 NAND2x1_ASAP7_75t_R _18042_ (.A(_01033_),
    .B(net5547),
    .Y(_09858_));
 OAI21x1_ASAP7_75t_R _18043_ (.A1(net5957),
    .A2(_09858_),
    .B(_09681_),
    .Y(_09859_));
 NAND2x1_ASAP7_75t_R _18044_ (.A(net5920),
    .B(_09859_),
    .Y(_09860_));
 NOR2x1_ASAP7_75t_R _18045_ (.A(_09857_),
    .B(_09860_),
    .Y(_09861_));
 NAND2x1_ASAP7_75t_R _18046_ (.A(_09645_),
    .B(net5963),
    .Y(_09862_));
 INVx1_ASAP7_75t_R _18047_ (.A(_09862_),
    .Y(_09863_));
 NAND2x1_ASAP7_75t_R _18048_ (.A(net5957),
    .B(net5268),
    .Y(_09864_));
 NOR2x1_ASAP7_75t_R _18049_ (.A(_09863_),
    .B(_09864_),
    .Y(_09865_));
 INVx1_ASAP7_75t_R _18050_ (.A(_09615_),
    .Y(_09866_));
 NAND2x1_ASAP7_75t_R _18051_ (.A(net5232),
    .B(net5964),
    .Y(_09867_));
 AO21x1_ASAP7_75t_R _18052_ (.A1(_09866_),
    .A2(_09867_),
    .B(_09773_),
    .Y(_09868_));
 NAND2x1_ASAP7_75t_R _18053_ (.A(_09601_),
    .B(net5964),
    .Y(_09869_));
 AO21x1_ASAP7_75t_R _18054_ (.A1(_09869_),
    .A2(net5544),
    .B(net6320),
    .Y(_09870_));
 NOR2x1_ASAP7_75t_R _18055_ (.A(_09813_),
    .B(_09829_),
    .Y(_09871_));
 AOI21x1_ASAP7_75t_R _18056_ (.A1(_09871_),
    .A2(_09870_),
    .B(net5954),
    .Y(_09872_));
 OAI21x1_ASAP7_75t_R _18057_ (.A1(_09865_),
    .A2(_09868_),
    .B(_09872_),
    .Y(_09873_));
 NOR2x1_ASAP7_75t_R _18058_ (.A(_09861_),
    .B(_09873_),
    .Y(_09874_));
 INVx1_ASAP7_75t_R _18059_ (.A(net4529),
    .Y(_09875_));
 OAI21x1_ASAP7_75t_R _18060_ (.A1(net5266),
    .A2(_09875_),
    .B(_09732_),
    .Y(_09876_));
 AND2x2_ASAP7_75t_R _18061_ (.A(_09772_),
    .B(net6293),
    .Y(_09877_));
 AOI21x1_ASAP7_75t_R _18062_ (.A1(_09877_),
    .A2(_09856_),
    .B(net6312),
    .Y(_09878_));
 NAND2x1_ASAP7_75t_R _18063_ (.A(_09876_),
    .B(_09878_),
    .Y(_09879_));
 NOR2x1_ASAP7_75t_R _18064_ (.A(net5957),
    .B(_09585_),
    .Y(_09880_));
 NAND2x1_ASAP7_75t_R _18065_ (.A(_09680_),
    .B(_09880_),
    .Y(_09881_));
 AO21x1_ASAP7_75t_R _18066_ (.A1(_09664_),
    .A2(_09609_),
    .B(net6320),
    .Y(_09882_));
 AOI21x1_ASAP7_75t_R _18067_ (.A1(_09881_),
    .A2(_09882_),
    .B(net6318),
    .Y(_09883_));
 AO21x1_ASAP7_75t_R _18068_ (.A1(_09828_),
    .A2(_09636_),
    .B(_08929_),
    .Y(_09884_));
 NAND2x1_ASAP7_75t_R _18069_ (.A(net6323),
    .B(net6325),
    .Y(_09885_));
 AO21x1_ASAP7_75t_R _18070_ (.A1(_09885_),
    .A2(_09688_),
    .B(net6320),
    .Y(_09886_));
 AOI21x1_ASAP7_75t_R _18071_ (.A1(_09884_),
    .A2(_09886_),
    .B(net6293),
    .Y(_09887_));
 OAI21x1_ASAP7_75t_R _18072_ (.A1(_09883_),
    .A2(_09887_),
    .B(net6312),
    .Y(_09888_));
 AOI21x1_ASAP7_75t_R _18073_ (.A1(_09879_),
    .A2(_09888_),
    .B(net5543),
    .Y(_09889_));
 OAI21x1_ASAP7_75t_R _18074_ (.A1(_09874_),
    .A2(_09889_),
    .B(net5953),
    .Y(_09890_));
 NAND2x1_ASAP7_75t_R _18075_ (.A(net6320),
    .B(_09604_),
    .Y(_09891_));
 AOI21x1_ASAP7_75t_R _18076_ (.A1(net4782),
    .A2(_09699_),
    .B(net6295),
    .Y(_09892_));
 NAND2x1_ASAP7_75t_R _18077_ (.A(net5957),
    .B(_09625_),
    .Y(_09893_));
 AOI21x1_ASAP7_75t_R _18078_ (.A1(_09893_),
    .A2(_09847_),
    .B(net6318),
    .Y(_09894_));
 OAI21x1_ASAP7_75t_R _18079_ (.A1(_09892_),
    .A2(_09894_),
    .B(net6312),
    .Y(_09895_));
 NOR2x1_ASAP7_75t_R _18080_ (.A(net5023),
    .B(_09615_),
    .Y(_09896_));
 INVx1_ASAP7_75t_R _18081_ (.A(_09896_),
    .Y(_09897_));
 NAND2x1_ASAP7_75t_R _18082_ (.A(net5547),
    .B(_09731_),
    .Y(_09898_));
 AOI21x1_ASAP7_75t_R _18083_ (.A1(_09897_),
    .A2(_09898_),
    .B(net6318),
    .Y(_09899_));
 AO21x1_ASAP7_75t_R _18084_ (.A1(_09644_),
    .A2(net5021),
    .B(net6320),
    .Y(_09900_));
 OA21x2_ASAP7_75t_R _18085_ (.A1(net5964),
    .A2(net5315),
    .B(net6320),
    .Y(_09901_));
 NAND2x1_ASAP7_75t_R _18086_ (.A(_09633_),
    .B(_09901_),
    .Y(_09902_));
 AOI21x1_ASAP7_75t_R _18087_ (.A1(_09900_),
    .A2(_09902_),
    .B(net6295),
    .Y(_09903_));
 OAI21x1_ASAP7_75t_R _18088_ (.A1(_09899_),
    .A2(_09903_),
    .B(net5920),
    .Y(_09904_));
 AOI21x1_ASAP7_75t_R _18089_ (.A1(_09895_),
    .A2(_09904_),
    .B(net5954),
    .Y(_09905_));
 NAND3x1_ASAP7_75t_R _18090_ (.A(net5547),
    .B(net5958),
    .C(net4967),
    .Y(_09906_));
 AOI21x1_ASAP7_75t_R _18091_ (.A1(_09780_),
    .A2(_09906_),
    .B(net6317),
    .Y(_09907_));
 OAI21x1_ASAP7_75t_R _18092_ (.A1(_09850_),
    .A2(_09907_),
    .B(net5920),
    .Y(_09908_));
 AND3x1_ASAP7_75t_R _18093_ (.A(net4783),
    .B(net6320),
    .C(net5234),
    .Y(_09909_));
 AND2x2_ASAP7_75t_R _18094_ (.A(_09893_),
    .B(net6318),
    .Y(_09910_));
 OAI21x1_ASAP7_75t_R _18095_ (.A1(net6320),
    .A2(_09574_),
    .B(_09910_),
    .Y(_09911_));
 AOI21x1_ASAP7_75t_R _18096_ (.A1(_09759_),
    .A2(_09690_),
    .B(net5920),
    .Y(_09912_));
 OAI21x1_ASAP7_75t_R _18097_ (.A1(_09909_),
    .A2(_09911_),
    .B(_09912_),
    .Y(_09913_));
 AOI21x1_ASAP7_75t_R _18098_ (.A1(_09908_),
    .A2(_09913_),
    .B(net5543),
    .Y(_09914_));
 OAI21x1_ASAP7_75t_R _18099_ (.A1(_09905_),
    .A2(_09914_),
    .B(_09598_),
    .Y(_09915_));
 NAND2x1_ASAP7_75t_R _18100_ (.A(_09915_),
    .B(_09890_),
    .Y(_00019_));
 NOR2x1_ASAP7_75t_R _18101_ (.A(net5231),
    .B(net6295),
    .Y(_09916_));
 NAND2x1_ASAP7_75t_R _18102_ (.A(_08929_),
    .B(net4967),
    .Y(_09917_));
 AO21x1_ASAP7_75t_R _18103_ (.A1(_09916_),
    .A2(_09917_),
    .B(_09653_),
    .Y(_09918_));
 AO21x1_ASAP7_75t_R _18104_ (.A1(net5547),
    .A2(_01038_),
    .B(net6320),
    .Y(_09919_));
 AND3x1_ASAP7_75t_R _18105_ (.A(_09771_),
    .B(_09919_),
    .C(net6295),
    .Y(_09920_));
 OAI21x1_ASAP7_75t_R _18106_ (.A1(_09918_),
    .A2(_09920_),
    .B(net6312),
    .Y(_09921_));
 NAND2x1_ASAP7_75t_R _18107_ (.A(net5956),
    .B(net5020),
    .Y(_09922_));
 AND3x1_ASAP7_75t_R _18108_ (.A(_09910_),
    .B(_09628_),
    .C(_09922_),
    .Y(_09923_));
 AO21x1_ASAP7_75t_R _18109_ (.A1(_09869_),
    .A2(net5267),
    .B(net5958),
    .Y(_09924_));
 AO21x1_ASAP7_75t_R _18110_ (.A1(_09707_),
    .A2(_09924_),
    .B(net5954),
    .Y(_09925_));
 NOR2x1_ASAP7_75t_R _18111_ (.A(_09923_),
    .B(_09925_),
    .Y(_09926_));
 OAI21x1_ASAP7_75t_R _18112_ (.A1(_09921_),
    .A2(_09926_),
    .B(net5953),
    .Y(_09927_));
 OA211x2_ASAP7_75t_R _18113_ (.A1(_09738_),
    .A2(net5230),
    .B(_09822_),
    .C(net6317),
    .Y(_09928_));
 NOR2x1_ASAP7_75t_R _18114_ (.A(_09863_),
    .B(_09849_),
    .Y(_09929_));
 OAI21x1_ASAP7_75t_R _18115_ (.A1(_09929_),
    .A2(_09767_),
    .B(net5543),
    .Y(_09930_));
 AND3x1_ASAP7_75t_R _18116_ (.A(_09633_),
    .B(net5961),
    .C(_09646_),
    .Y(_09931_));
 NAND2x1_ASAP7_75t_R _18117_ (.A(_09885_),
    .B(_09737_),
    .Y(_09932_));
 NOR2x1_ASAP7_75t_R _18118_ (.A(net5961),
    .B(_09932_),
    .Y(_09933_));
 OAI21x1_ASAP7_75t_R _18119_ (.A1(_09931_),
    .A2(_09933_),
    .B(net6314),
    .Y(_09934_));
 AOI21x1_ASAP7_75t_R _18120_ (.A1(_09778_),
    .A2(_09804_),
    .B(_09653_),
    .Y(_09935_));
 AOI21x1_ASAP7_75t_R _18121_ (.A1(_09934_),
    .A2(_09935_),
    .B(net6313),
    .Y(_09936_));
 OA21x2_ASAP7_75t_R _18122_ (.A1(_09928_),
    .A2(_09930_),
    .B(_09936_),
    .Y(_09937_));
 NAND2x1_ASAP7_75t_R _18123_ (.A(net6318),
    .B(_09906_),
    .Y(_09938_));
 OAI21x1_ASAP7_75t_R _18124_ (.A1(_09933_),
    .A2(_09938_),
    .B(_09653_),
    .Y(_09939_));
 AND3x1_ASAP7_75t_R _18125_ (.A(_09662_),
    .B(net6295),
    .C(_09648_),
    .Y(_09940_));
 NOR2x1_ASAP7_75t_R _18126_ (.A(_09939_),
    .B(_09940_),
    .Y(_09941_));
 AOI22x1_ASAP7_75t_R _18127_ (.A1(_09657_),
    .A2(net5234),
    .B1(net6322),
    .B2(net5959),
    .Y(_09942_));
 AO21x1_ASAP7_75t_R _18128_ (.A1(_09942_),
    .A2(net6295),
    .B(_09653_),
    .Y(_09943_));
 NOR2x1_ASAP7_75t_R _18129_ (.A(net5960),
    .B(_09758_),
    .Y(_09944_));
 INVx1_ASAP7_75t_R _18130_ (.A(_09944_),
    .Y(_09945_));
 OA21x2_ASAP7_75t_R _18131_ (.A1(_09945_),
    .A2(_09863_),
    .B(_09777_),
    .Y(_09946_));
 OAI21x1_ASAP7_75t_R _18132_ (.A1(_09943_),
    .A2(_09946_),
    .B(net5919),
    .Y(_09947_));
 NOR2x1_ASAP7_75t_R _18133_ (.A(net5020),
    .B(_09754_),
    .Y(_09948_));
 NAND2x1_ASAP7_75t_R _18134_ (.A(net6316),
    .B(net5229),
    .Y(_09949_));
 OA21x2_ASAP7_75t_R _18135_ (.A1(_09949_),
    .A2(_09746_),
    .B(net5954),
    .Y(_09950_));
 OAI21x1_ASAP7_75t_R _18136_ (.A1(_09948_),
    .A2(_09593_),
    .B(_09950_),
    .Y(_09951_));
 OA21x2_ASAP7_75t_R _18137_ (.A1(_09668_),
    .A2(net5957),
    .B(net6293),
    .Y(_09952_));
 AOI21x1_ASAP7_75t_R _18138_ (.A1(_09864_),
    .A2(_09952_),
    .B(net5954),
    .Y(_09953_));
 NOR2x1_ASAP7_75t_R _18139_ (.A(_09568_),
    .B(_09917_),
    .Y(_09954_));
 AO21x1_ASAP7_75t_R _18140_ (.A1(net6320),
    .A2(_09685_),
    .B(net6293),
    .Y(_09955_));
 OR2x2_ASAP7_75t_R _18141_ (.A(_09954_),
    .B(_09955_),
    .Y(_09956_));
 AOI21x1_ASAP7_75t_R _18142_ (.A1(_09953_),
    .A2(_09956_),
    .B(net5920),
    .Y(_09957_));
 AOI21x1_ASAP7_75t_R _18143_ (.A1(_09951_),
    .A2(_09957_),
    .B(net5953),
    .Y(_09958_));
 OAI21x1_ASAP7_75t_R _18144_ (.A1(_09941_),
    .A2(_09947_),
    .B(_09958_),
    .Y(_09959_));
 OAI21x1_ASAP7_75t_R _18145_ (.A1(_09927_),
    .A2(_09937_),
    .B(_09959_),
    .Y(_00020_));
 OA21x2_ASAP7_75t_R _18146_ (.A1(_09731_),
    .A2(_09622_),
    .B(net6317),
    .Y(_09960_));
 AO21x1_ASAP7_75t_R _18147_ (.A1(_09729_),
    .A2(net5233),
    .B(net5960),
    .Y(_09961_));
 AOI21x1_ASAP7_75t_R _18148_ (.A1(_09638_),
    .A2(_09961_),
    .B(net6315),
    .Y(_09962_));
 OAI21x1_ASAP7_75t_R _18149_ (.A1(_09960_),
    .A2(_09962_),
    .B(net6312),
    .Y(_09963_));
 NOR2x1_ASAP7_75t_R _18150_ (.A(net5232),
    .B(net6320),
    .Y(_09964_));
 OA21x2_ASAP7_75t_R _18151_ (.A1(_09880_),
    .A2(_09964_),
    .B(net6293),
    .Y(_09965_));
 AO21x1_ASAP7_75t_R _18152_ (.A1(_09667_),
    .A2(_09636_),
    .B(net6320),
    .Y(_09966_));
 AO21x1_ASAP7_75t_R _18153_ (.A1(_09828_),
    .A2(_09821_),
    .B(net5957),
    .Y(_09967_));
 AOI21x1_ASAP7_75t_R _18154_ (.A1(_09966_),
    .A2(_09967_),
    .B(net6293),
    .Y(_09968_));
 OAI21x1_ASAP7_75t_R _18155_ (.A1(_09965_),
    .A2(_09968_),
    .B(net5920),
    .Y(_09969_));
 AOI21x1_ASAP7_75t_R _18156_ (.A1(_09963_),
    .A2(_09969_),
    .B(net5954),
    .Y(_09970_));
 OA21x2_ASAP7_75t_R _18157_ (.A1(_09792_),
    .A2(_09712_),
    .B(net6320),
    .Y(_09971_));
 AO21x1_ASAP7_75t_R _18158_ (.A1(net6321),
    .A2(_09964_),
    .B(net6293),
    .Y(_09972_));
 AO21x1_ASAP7_75t_R _18159_ (.A1(net5234),
    .A2(_09880_),
    .B(_09972_),
    .Y(_09973_));
 OAI21x1_ASAP7_75t_R _18160_ (.A1(_09971_),
    .A2(_09593_),
    .B(_09973_),
    .Y(_09974_));
 AOI21x1_ASAP7_75t_R _18161_ (.A1(_09569_),
    .A2(net4529),
    .B(_09773_),
    .Y(_09975_));
 OAI21x1_ASAP7_75t_R _18162_ (.A1(net5022),
    .A2(_09772_),
    .B(_09975_),
    .Y(_09976_));
 AOI21x1_ASAP7_75t_R _18163_ (.A1(net6296),
    .A2(_08929_),
    .B(_09813_),
    .Y(_09977_));
 AOI21x1_ASAP7_75t_R _18164_ (.A1(_09659_),
    .A2(_09977_),
    .B(_09653_),
    .Y(_09978_));
 NAND2x1_ASAP7_75t_R _18165_ (.A(_09976_),
    .B(_09978_),
    .Y(_09979_));
 AOI21x1_ASAP7_75t_R _18166_ (.A1(net5920),
    .A2(_09974_),
    .B(_09979_),
    .Y(_09980_));
 OAI21x1_ASAP7_75t_R _18167_ (.A1(_09970_),
    .A2(_09980_),
    .B(_09598_),
    .Y(_09981_));
 AO21x1_ASAP7_75t_R _18168_ (.A1(net4783),
    .A2(net6319),
    .B(net6315),
    .Y(_09982_));
 AO21x1_ASAP7_75t_R _18169_ (.A1(_09574_),
    .A2(net4969),
    .B(net6319),
    .Y(_09983_));
 INVx1_ASAP7_75t_R _18170_ (.A(_09983_),
    .Y(_09984_));
 AND2x2_ASAP7_75t_R _18171_ (.A(net6315),
    .B(net5233),
    .Y(_09985_));
 AOI21x1_ASAP7_75t_R _18172_ (.A1(_09754_),
    .A2(_09985_),
    .B(net6313),
    .Y(_09986_));
 OAI21x1_ASAP7_75t_R _18173_ (.A1(_09982_),
    .A2(_09984_),
    .B(_09986_),
    .Y(_09987_));
 NOR2x1_ASAP7_75t_R _18174_ (.A(_09730_),
    .B(_09614_),
    .Y(_09988_));
 AO21x1_ASAP7_75t_R _18175_ (.A1(_09944_),
    .A2(_09583_),
    .B(net6315),
    .Y(_09989_));
 NAND2x1_ASAP7_75t_R _18176_ (.A(net5547),
    .B(_09838_),
    .Y(_09990_));
 NAND2x1_ASAP7_75t_R _18177_ (.A(net5546),
    .B(net5964),
    .Y(_09991_));
 AOI21x1_ASAP7_75t_R _18178_ (.A1(_09991_),
    .A2(net4529),
    .B(net6294),
    .Y(_09992_));
 AOI21x1_ASAP7_75t_R _18179_ (.A1(_09990_),
    .A2(_09992_),
    .B(net5920),
    .Y(_09993_));
 OAI21x1_ASAP7_75t_R _18180_ (.A1(_09988_),
    .A2(_09989_),
    .B(_09993_),
    .Y(_09994_));
 AOI21x1_ASAP7_75t_R _18181_ (.A1(_09987_),
    .A2(_09994_),
    .B(_09653_),
    .Y(_09995_));
 NAND2x1_ASAP7_75t_R _18182_ (.A(_09633_),
    .B(_09746_),
    .Y(_09996_));
 AOI21x1_ASAP7_75t_R _18183_ (.A1(_09922_),
    .A2(_09996_),
    .B(net6295),
    .Y(_09997_));
 AO21x1_ASAP7_75t_R _18184_ (.A1(net6320),
    .A2(_09821_),
    .B(net6317),
    .Y(_09998_));
 AOI21x1_ASAP7_75t_R _18185_ (.A1(net4785),
    .A2(_09646_),
    .B(_09998_),
    .Y(_09999_));
 OAI21x1_ASAP7_75t_R _18186_ (.A1(_09997_),
    .A2(_09999_),
    .B(net5920),
    .Y(_10000_));
 AO21x1_ASAP7_75t_R _18187_ (.A1(net5965),
    .A2(net5962),
    .B(net6314),
    .Y(_10001_));
 NOR2x1_ASAP7_75t_R _18188_ (.A(_10001_),
    .B(_09933_),
    .Y(_10002_));
 AND3x1_ASAP7_75t_R _18189_ (.A(_09729_),
    .B(net5961),
    .C(_09636_),
    .Y(_10003_));
 NAND2x1_ASAP7_75t_R _18190_ (.A(net6296),
    .B(net6323),
    .Y(_10004_));
 AO21x1_ASAP7_75t_R _18191_ (.A1(_09866_),
    .A2(_10004_),
    .B(net6293),
    .Y(_10005_));
 NOR2x1_ASAP7_75t_R _18192_ (.A(_10003_),
    .B(_10005_),
    .Y(_10006_));
 OAI21x1_ASAP7_75t_R _18193_ (.A1(_10002_),
    .A2(_10006_),
    .B(net6313),
    .Y(_10007_));
 AOI21x1_ASAP7_75t_R _18194_ (.A1(_10000_),
    .A2(_10007_),
    .B(net5954),
    .Y(_10008_));
 OAI21x1_ASAP7_75t_R _18195_ (.A1(_09995_),
    .A2(_10008_),
    .B(net5953),
    .Y(_10009_));
 NAND2x1_ASAP7_75t_R _18196_ (.A(_09981_),
    .B(_10009_),
    .Y(_00021_));
 AND2x2_ASAP7_75t_R _18197_ (.A(_09657_),
    .B(net5267),
    .Y(_10010_));
 NAND2x1_ASAP7_75t_R _18198_ (.A(_09583_),
    .B(_09833_),
    .Y(_10011_));
 AOI21x1_ASAP7_75t_R _18199_ (.A1(net5548),
    .A2(net4529),
    .B(net6316),
    .Y(_10012_));
 NAND2x1_ASAP7_75t_R _18200_ (.A(_10011_),
    .B(_10012_),
    .Y(_10013_));
 OAI21x1_ASAP7_75t_R _18201_ (.A1(_10010_),
    .A2(_09911_),
    .B(_10013_),
    .Y(_10014_));
 INVx1_ASAP7_75t_R _18202_ (.A(_09910_),
    .Y(_10015_));
 OA21x2_ASAP7_75t_R _18203_ (.A1(_09674_),
    .A2(net5962),
    .B(net6313),
    .Y(_10016_));
 OAI21x1_ASAP7_75t_R _18204_ (.A1(net6319),
    .A2(_09830_),
    .B(_10016_),
    .Y(_10017_));
 NOR2x1_ASAP7_75t_R _18205_ (.A(net5962),
    .B(net6323),
    .Y(_10018_));
 NOR2x1_ASAP7_75t_R _18206_ (.A(_10018_),
    .B(_09813_),
    .Y(_10019_));
 OAI21x1_ASAP7_75t_R _18207_ (.A1(net6319),
    .A2(_09932_),
    .B(_10019_),
    .Y(_10020_));
 OAI21x1_ASAP7_75t_R _18208_ (.A1(_10015_),
    .A2(_10017_),
    .B(_10020_),
    .Y(_10021_));
 AOI21x1_ASAP7_75t_R _18209_ (.A1(net5919),
    .A2(_10014_),
    .B(_10021_),
    .Y(_10022_));
 AND3x1_ASAP7_75t_R _18210_ (.A(_09688_),
    .B(_09577_),
    .C(net6319),
    .Y(_10023_));
 AOI21x1_ASAP7_75t_R _18211_ (.A1(net5547),
    .A2(_09885_),
    .B(net6320),
    .Y(_10024_));
 NOR3x1_ASAP7_75t_R _18212_ (.A(_10023_),
    .B(net6295),
    .C(_10024_),
    .Y(_10025_));
 NOR2x1_ASAP7_75t_R _18213_ (.A(net5961),
    .B(_09786_),
    .Y(_10026_));
 OAI21x1_ASAP7_75t_R _18214_ (.A1(_10026_),
    .A2(_10024_),
    .B(net6295),
    .Y(_10027_));
 NAND2x1_ASAP7_75t_R _18215_ (.A(net6313),
    .B(_10027_),
    .Y(_10028_));
 OA21x2_ASAP7_75t_R _18216_ (.A1(_09667_),
    .A2(net5959),
    .B(net6295),
    .Y(_10029_));
 NAND2x1_ASAP7_75t_R _18217_ (.A(_10029_),
    .B(_09983_),
    .Y(_10030_));
 INVx1_ASAP7_75t_R _18218_ (.A(_09762_),
    .Y(_10031_));
 AOI21x1_ASAP7_75t_R _18219_ (.A1(_09611_),
    .A2(_10031_),
    .B(net6313),
    .Y(_10032_));
 AOI21x1_ASAP7_75t_R _18220_ (.A1(_10030_),
    .A2(_10032_),
    .B(net5953),
    .Y(_10033_));
 OAI21x1_ASAP7_75t_R _18221_ (.A1(_10025_),
    .A2(_10028_),
    .B(_10033_),
    .Y(_10034_));
 OAI21x1_ASAP7_75t_R _18222_ (.A1(_09598_),
    .A2(_10022_),
    .B(_10034_),
    .Y(_10035_));
 OAI21x1_ASAP7_75t_R _18223_ (.A1(_09758_),
    .A2(net5230),
    .B(_09698_),
    .Y(_10036_));
 AOI21x1_ASAP7_75t_R _18224_ (.A1(net5268),
    .A2(_09657_),
    .B(net6316),
    .Y(_10037_));
 OAI21x1_ASAP7_75t_R _18225_ (.A1(_09753_),
    .A2(net5230),
    .B(_10037_),
    .Y(_10038_));
 AOI21x1_ASAP7_75t_R _18226_ (.A1(_10036_),
    .A2(_10038_),
    .B(net6312),
    .Y(_10039_));
 NAND2x1_ASAP7_75t_R _18227_ (.A(_09667_),
    .B(_09746_),
    .Y(_10040_));
 AO21x1_ASAP7_75t_R _18228_ (.A1(_09633_),
    .A2(net5233),
    .B(net6320),
    .Y(_10041_));
 AOI21x1_ASAP7_75t_R _18229_ (.A1(_10040_),
    .A2(_10041_),
    .B(net6317),
    .Y(_10042_));
 NAND2x1_ASAP7_75t_R _18230_ (.A(net6318),
    .B(_09891_),
    .Y(_10043_));
 OAI21x1_ASAP7_75t_R _18231_ (.A1(_10043_),
    .A2(_09789_),
    .B(net6313),
    .Y(_10044_));
 OAI21x1_ASAP7_75t_R _18232_ (.A1(_10042_),
    .A2(_10044_),
    .B(net5953),
    .Y(_10045_));
 NOR2x1_ASAP7_75t_R _18233_ (.A(_10039_),
    .B(_10045_),
    .Y(_10046_));
 NAND2x1_ASAP7_75t_R _18234_ (.A(net5920),
    .B(_09825_),
    .Y(_10047_));
 OA21x2_ASAP7_75t_R _18235_ (.A1(_09954_),
    .A2(_09901_),
    .B(net6316),
    .Y(_10048_));
 NOR2x1_ASAP7_75t_R _18236_ (.A(_10047_),
    .B(_10048_),
    .Y(_10049_));
 NOR2x1_ASAP7_75t_R _18237_ (.A(net6320),
    .B(net5266),
    .Y(_10050_));
 AND2x2_ASAP7_75t_R _18238_ (.A(_10050_),
    .B(net5234),
    .Y(_10051_));
 NOR2x1_ASAP7_75t_R _18239_ (.A(net5955),
    .B(net5918),
    .Y(_10052_));
 OR3x1_ASAP7_75t_R _18240_ (.A(_10052_),
    .B(net6295),
    .C(net5920),
    .Y(_10053_));
 NAND2x1_ASAP7_75t_R _18241_ (.A(_09569_),
    .B(net4529),
    .Y(_10054_));
 AOI211x1_ASAP7_75t_R _18242_ (.A1(_01032_),
    .A2(net5959),
    .B(net5920),
    .C(net6317),
    .Y(_10055_));
 AOI21x1_ASAP7_75t_R _18243_ (.A1(_10054_),
    .A2(_10055_),
    .B(net5953),
    .Y(_10056_));
 OAI21x1_ASAP7_75t_R _18244_ (.A1(_10051_),
    .A2(_10053_),
    .B(_10056_),
    .Y(_10057_));
 OAI21x1_ASAP7_75t_R _18245_ (.A1(_10049_),
    .A2(_10057_),
    .B(net5542),
    .Y(_10058_));
 NOR2x1_ASAP7_75t_R _18246_ (.A(_10046_),
    .B(_10058_),
    .Y(_10059_));
 AOI21x1_ASAP7_75t_R _18247_ (.A1(net5954),
    .A2(_10035_),
    .B(_10059_),
    .Y(_00022_));
 NOR2x1_ASAP7_75t_R _18248_ (.A(net6315),
    .B(_09863_),
    .Y(_10060_));
 AO21x1_ASAP7_75t_R _18249_ (.A1(net5961),
    .A2(net5921),
    .B(_09746_),
    .Y(_10061_));
 AOI21x1_ASAP7_75t_R _18250_ (.A1(_10060_),
    .A2(_10061_),
    .B(net6313),
    .Y(_10062_));
 NOR2x1_ASAP7_75t_R _18251_ (.A(net6320),
    .B(_09932_),
    .Y(_10063_));
 OAI21x1_ASAP7_75t_R _18252_ (.A1(_09725_),
    .A2(_10063_),
    .B(net6318),
    .Y(_10064_));
 NAND2x1_ASAP7_75t_R _18253_ (.A(_10062_),
    .B(_10064_),
    .Y(_10065_));
 OA21x2_ASAP7_75t_R _18254_ (.A1(net5963),
    .A2(_01019_),
    .B(net6320),
    .Y(_10066_));
 OA21x2_ASAP7_75t_R _18255_ (.A1(_09637_),
    .A2(net5022),
    .B(net5961),
    .Y(_10067_));
 AOI211x1_ASAP7_75t_R _18256_ (.A1(net4966),
    .A2(_10066_),
    .B(_10067_),
    .C(_09813_),
    .Y(_10068_));
 AO21x1_ASAP7_75t_R _18257_ (.A1(_10066_),
    .A2(_09633_),
    .B(net5920),
    .Y(_10069_));
 OAI21x1_ASAP7_75t_R _18258_ (.A1(_10069_),
    .A2(_09938_),
    .B(net5954),
    .Y(_10070_));
 NOR2x1_ASAP7_75t_R _18259_ (.A(_10068_),
    .B(_10070_),
    .Y(_10071_));
 AOI21x1_ASAP7_75t_R _18260_ (.A1(_10065_),
    .A2(_10071_),
    .B(_09598_),
    .Y(_10072_));
 AOI211x1_ASAP7_75t_R _18261_ (.A1(_10050_),
    .A2(net5021),
    .B(_09812_),
    .C(_10052_),
    .Y(_10073_));
 AO21x1_ASAP7_75t_R _18262_ (.A1(net4969),
    .A2(net5021),
    .B(net5957),
    .Y(_10074_));
 OR2x2_ASAP7_75t_R _18263_ (.A(_01038_),
    .B(net6320),
    .Y(_10075_));
 AO21x1_ASAP7_75t_R _18264_ (.A1(_10074_),
    .A2(_10075_),
    .B(net6317),
    .Y(_10076_));
 OAI21x1_ASAP7_75t_R _18265_ (.A1(net6295),
    .A2(_10073_),
    .B(_10076_),
    .Y(_10077_));
 AOI21x1_ASAP7_75t_R _18266_ (.A1(_09991_),
    .A2(_09944_),
    .B(net5919),
    .Y(_10078_));
 NOR2x1_ASAP7_75t_R _18267_ (.A(_01019_),
    .B(net6320),
    .Y(_10079_));
 AO21x1_ASAP7_75t_R _18268_ (.A1(_09830_),
    .A2(net6320),
    .B(_10079_),
    .Y(_10080_));
 INVx1_ASAP7_75t_R _18269_ (.A(_09813_),
    .Y(_10081_));
 AO21x1_ASAP7_75t_R _18270_ (.A1(_10080_),
    .A2(_10081_),
    .B(net5954),
    .Y(_10082_));
 AOI21x1_ASAP7_75t_R _18271_ (.A1(_09777_),
    .A2(_10078_),
    .B(_10082_),
    .Y(_10083_));
 OAI21x1_ASAP7_75t_R _18272_ (.A1(net6313),
    .A2(_10077_),
    .B(_10083_),
    .Y(_10084_));
 AND2x2_ASAP7_75t_R _18273_ (.A(net5021),
    .B(net5955),
    .Y(_10085_));
 AOI211x1_ASAP7_75t_R _18274_ (.A1(net5548),
    .A2(_10085_),
    .B(_09896_),
    .C(net6294),
    .Y(_10086_));
 AND2x2_ASAP7_75t_R _18275_ (.A(_10012_),
    .B(_09807_),
    .Y(_10087_));
 OAI21x1_ASAP7_75t_R _18276_ (.A1(_10086_),
    .A2(_10087_),
    .B(net5920),
    .Y(_10088_));
 AOI221x1_ASAP7_75t_R _18277_ (.A1(_09991_),
    .A2(_09866_),
    .B1(net4966),
    .B2(_09833_),
    .C(_09773_),
    .Y(_10089_));
 AO21x1_ASAP7_75t_R _18278_ (.A1(net6320),
    .A2(_09577_),
    .B(_09813_),
    .Y(_10090_));
 OAI21x1_ASAP7_75t_R _18279_ (.A1(net4528),
    .A2(_10090_),
    .B(net5954),
    .Y(_10091_));
 NOR2x1_ASAP7_75t_R _18280_ (.A(_10089_),
    .B(_10091_),
    .Y(_10092_));
 AOI21x1_ASAP7_75t_R _18281_ (.A1(_10088_),
    .A2(_10092_),
    .B(net5953),
    .Y(_10093_));
 NAND2x1_ASAP7_75t_R _18282_ (.A(_09569_),
    .B(_10066_),
    .Y(_10094_));
 AO21x1_ASAP7_75t_R _18283_ (.A1(net6296),
    .A2(net6320),
    .B(net6293),
    .Y(_10095_));
 NOR2x1_ASAP7_75t_R _18284_ (.A(_09738_),
    .B(_09638_),
    .Y(_10096_));
 OAI21x1_ASAP7_75t_R _18285_ (.A1(_10095_),
    .A2(_10096_),
    .B(net6313),
    .Y(_10097_));
 AOI21x1_ASAP7_75t_R _18286_ (.A1(_09804_),
    .A2(_10094_),
    .B(_10097_),
    .Y(_10098_));
 AO21x1_ASAP7_75t_R _18287_ (.A1(net5961),
    .A2(_09729_),
    .B(_09982_),
    .Y(_10099_));
 AO21x1_ASAP7_75t_R _18288_ (.A1(_09828_),
    .A2(_09669_),
    .B(net5957),
    .Y(_10100_));
 AO21x1_ASAP7_75t_R _18289_ (.A1(_10100_),
    .A2(net5230),
    .B(net6293),
    .Y(_10101_));
 AOI21x1_ASAP7_75t_R _18290_ (.A1(_10099_),
    .A2(_10101_),
    .B(net6313),
    .Y(_10102_));
 OAI21x1_ASAP7_75t_R _18291_ (.A1(_10098_),
    .A2(_10102_),
    .B(_09653_),
    .Y(_10103_));
 AOI22x1_ASAP7_75t_R _18292_ (.A1(_10072_),
    .A2(_10084_),
    .B1(_10093_),
    .B2(_10103_),
    .Y(_00023_));
 OAI21x1_ASAP7_75t_R _18294_ (.A1(_09004_),
    .A2(_08798_),
    .B(net6679),
    .Y(_10104_));
 NAND2x1_ASAP7_75t_R _18295_ (.A(net6687),
    .B(net47),
    .Y(_10105_));
 OAI21x1_ASAP7_75t_R _18296_ (.A1(_09003_),
    .A2(_10104_),
    .B(_10105_),
    .Y(_10106_));
 NOR2x1_ASAP7_75t_R _18299_ (.A(_08985_),
    .B(_08787_),
    .Y(_10108_));
 OAI21x1_ASAP7_75t_R _18300_ (.A1(_08986_),
    .A2(_08988_),
    .B(_08030_),
    .Y(_10109_));
 INVx1_ASAP7_75t_R _18301_ (.A(_08991_),
    .Y(_10110_));
 OAI21x1_ASAP7_75t_R _18302_ (.A1(_10108_),
    .A2(_10109_),
    .B(_10110_),
    .Y(_10111_));
 NAND2x1_ASAP7_75t_R _18305_ (.A(net5565),
    .B(net6289),
    .Y(_10113_));
 OA21x2_ASAP7_75t_R _18306_ (.A1(_10113_),
    .A2(net5934),
    .B(net6297),
    .Y(_10114_));
 INVx1_ASAP7_75t_R _18307_ (.A(_10114_),
    .Y(_10115_));
 INVx1_ASAP7_75t_R _18310_ (.A(_01048_),
    .Y(_10118_));
 AO21x1_ASAP7_75t_R _18311_ (.A1(net6298),
    .A2(net6388),
    .B(net5228),
    .Y(_10119_));
 INVx1_ASAP7_75t_R _18313_ (.A(_01051_),
    .Y(_10121_));
 NAND2x1_ASAP7_75t_R _18314_ (.A(_10121_),
    .B(net6290),
    .Y(_10122_));
 INVx1_ASAP7_75t_R _18315_ (.A(_10122_),
    .Y(_10123_));
 NAND2x1_ASAP7_75t_R _18316_ (.A(net5934),
    .B(_10123_),
    .Y(_10124_));
 OAI21x1_ASAP7_75t_R _18317_ (.A1(net5934),
    .A2(net4965),
    .B(_10124_),
    .Y(_10125_));
 INVx2_ASAP7_75t_R _18318_ (.A(_09016_),
    .Y(_10126_));
 NAND2x1_ASAP7_75t_R _18320_ (.A(net5539),
    .B(_10123_),
    .Y(_10128_));
 INVx1_ASAP7_75t_R _18321_ (.A(_01049_),
    .Y(_10129_));
 NOR2x1_ASAP7_75t_R _18322_ (.A(_10129_),
    .B(net6292),
    .Y(_10130_));
 INVx1_ASAP7_75t_R _18323_ (.A(_10130_),
    .Y(_10131_));
 OA21x2_ASAP7_75t_R _18325_ (.A1(net5939),
    .A2(net5565),
    .B(net5934),
    .Y(_10133_));
 AOI21x1_ASAP7_75t_R _18326_ (.A1(_10131_),
    .A2(_10133_),
    .B(net6297),
    .Y(_10134_));
 AOI21x1_ASAP7_75t_R _18328_ (.A1(_10128_),
    .A2(_10134_),
    .B(net5933),
    .Y(_10136_));
 OAI21x1_ASAP7_75t_R _18329_ (.A1(_10115_),
    .A2(_10125_),
    .B(_10136_),
    .Y(_10137_));
 NAND2x1_ASAP7_75t_R _18330_ (.A(net6302),
    .B(_09007_),
    .Y(_10138_));
 AO21x1_ASAP7_75t_R _18331_ (.A1(_10138_),
    .A2(_10113_),
    .B(net5934),
    .Y(_10139_));
 INVx2_ASAP7_75t_R _18332_ (.A(_09021_),
    .Y(_10140_));
 NOR2x1_ASAP7_75t_R _18334_ (.A(net6301),
    .B(net6291),
    .Y(_10142_));
 NAND2x1_ASAP7_75t_R _18335_ (.A(_01050_),
    .B(_10106_),
    .Y(_10143_));
 INVx1_ASAP7_75t_R _18336_ (.A(_10143_),
    .Y(_10144_));
 OAI21x1_ASAP7_75t_R _18337_ (.A1(_10142_),
    .A2(_10144_),
    .B(net5935),
    .Y(_10145_));
 NAND3x1_ASAP7_75t_R _18338_ (.A(_10139_),
    .B(_10140_),
    .C(_10145_),
    .Y(_10146_));
 NOR2x1_ASAP7_75t_R _18339_ (.A(net5562),
    .B(net6292),
    .Y(_10147_));
 AO21x1_ASAP7_75t_R _18341_ (.A1(_10147_),
    .A2(net5539),
    .B(_10140_),
    .Y(_10149_));
 NOR2x1_ASAP7_75t_R _18343_ (.A(_01055_),
    .B(net5539),
    .Y(_10151_));
 OA21x2_ASAP7_75t_R _18344_ (.A1(_10149_),
    .A2(_10151_),
    .B(net5933),
    .Y(_10152_));
 AOI21x1_ASAP7_75t_R _18345_ (.A1(_10146_),
    .A2(_10152_),
    .B(net5932),
    .Y(_10153_));
 NAND2x1_ASAP7_75t_R _18346_ (.A(_10137_),
    .B(_10153_),
    .Y(_10154_));
 NAND2x1_ASAP7_75t_R _18347_ (.A(net6292),
    .B(_01042_),
    .Y(_10155_));
 NAND2x1p5_ASAP7_75t_R _18348_ (.A(_10155_),
    .B(net5937),
    .Y(_10156_));
 AO21x1_ASAP7_75t_R _18349_ (.A1(net6298),
    .A2(net6388),
    .B(_01046_),
    .Y(_10157_));
 NAND2x1_ASAP7_75t_R _18350_ (.A(_10129_),
    .B(net6290),
    .Y(_10158_));
 AO21x1_ASAP7_75t_R _18351_ (.A1(_10157_),
    .A2(net4962),
    .B(net5936),
    .Y(_10159_));
 AOI21x1_ASAP7_75t_R _18353_ (.A1(_10156_),
    .A2(_10159_),
    .B(net5917),
    .Y(_10161_));
 NOR2x1_ASAP7_75t_R _18354_ (.A(net5564),
    .B(net6289),
    .Y(_10162_));
 NAND2x1_ASAP7_75t_R _18355_ (.A(net5541),
    .B(_10162_),
    .Y(_10163_));
 NAND2x1_ASAP7_75t_R _18356_ (.A(net6287),
    .B(_09007_),
    .Y(_10164_));
 NAND2x1_ASAP7_75t_R _18357_ (.A(_01041_),
    .B(net6292),
    .Y(_10165_));
 AO21x1_ASAP7_75t_R _18358_ (.A1(_10164_),
    .A2(net5537),
    .B(net5541),
    .Y(_10166_));
 AOI21x1_ASAP7_75t_R _18360_ (.A1(_10163_),
    .A2(_10166_),
    .B(net6297),
    .Y(_10168_));
 OAI21x1_ASAP7_75t_R _18362_ (.A1(_10161_),
    .A2(_10168_),
    .B(net5933),
    .Y(_10170_));
 NAND2x1_ASAP7_75t_R _18363_ (.A(net6287),
    .B(net6289),
    .Y(_10171_));
 AO21x1_ASAP7_75t_R _18364_ (.A1(_10171_),
    .A2(_10119_),
    .B(net5539),
    .Y(_10172_));
 AO21x1_ASAP7_75t_R _18365_ (.A1(net6298),
    .A2(net6388),
    .B(_01042_),
    .Y(_10173_));
 AOI21x1_ASAP7_75t_R _18368_ (.A1(net6289),
    .A2(net6299),
    .B(net5937),
    .Y(_10176_));
 AOI21x1_ASAP7_75t_R _18370_ (.A1(net5262),
    .A2(_10176_),
    .B(net6297),
    .Y(_10178_));
 AOI21x1_ASAP7_75t_R _18371_ (.A1(_10172_),
    .A2(_10178_),
    .B(net5933),
    .Y(_10179_));
 INVx1_ASAP7_75t_R _18372_ (.A(_01050_),
    .Y(_10180_));
 AO21x1_ASAP7_75t_R _18373_ (.A1(net6298),
    .A2(net6388),
    .B(_10180_),
    .Y(_10181_));
 AO21x1_ASAP7_75t_R _18374_ (.A1(_10181_),
    .A2(net4964),
    .B(net5935),
    .Y(_10182_));
 NAND2x1_ASAP7_75t_R _18376_ (.A(net5564),
    .B(net6289),
    .Y(_10184_));
 NAND2x1_ASAP7_75t_R _18377_ (.A(net5936),
    .B(_10184_),
    .Y(_10185_));
 NAND3x1_ASAP7_75t_R _18378_ (.A(_10182_),
    .B(net6297),
    .C(_10185_),
    .Y(_10186_));
 INVx1_ASAP7_75t_R _18379_ (.A(_09030_),
    .Y(_10187_));
 AOI21x1_ASAP7_75t_R _18380_ (.A1(_10179_),
    .A2(_10186_),
    .B(net5536),
    .Y(_10188_));
 INVx1_ASAP7_75t_R _18381_ (.A(_09034_),
    .Y(_10189_));
 AOI21x1_ASAP7_75t_R _18382_ (.A1(_10170_),
    .A2(_10188_),
    .B(_10189_),
    .Y(_10190_));
 NAND2x1_ASAP7_75t_R _18383_ (.A(_10154_),
    .B(_10190_),
    .Y(_10191_));
 NOR2x1_ASAP7_75t_R _18384_ (.A(net6287),
    .B(net6300),
    .Y(_10192_));
 NOR2x1_ASAP7_75t_R _18385_ (.A(net6301),
    .B(_09007_),
    .Y(_10193_));
 OAI21x1_ASAP7_75t_R _18387_ (.A1(_10192_),
    .A2(_10193_),
    .B(net5935),
    .Y(_10195_));
 INVx1_ASAP7_75t_R _18388_ (.A(_10192_),
    .Y(_10196_));
 AOI21x1_ASAP7_75t_R _18389_ (.A1(net6287),
    .A2(net6289),
    .B(net5937),
    .Y(_10197_));
 NAND2x1_ASAP7_75t_R _18390_ (.A(_10196_),
    .B(_10197_),
    .Y(_10198_));
 AOI21x1_ASAP7_75t_R _18391_ (.A1(_10195_),
    .A2(_10198_),
    .B(net5913),
    .Y(_10199_));
 AO21x1_ASAP7_75t_R _18392_ (.A1(net6298),
    .A2(net6388),
    .B(net5567),
    .Y(_10200_));
 AOI21x1_ASAP7_75t_R _18393_ (.A1(net5562),
    .A2(net6292),
    .B(net5937),
    .Y(_10201_));
 NAND2x1_ASAP7_75t_R _18394_ (.A(_10200_),
    .B(_10201_),
    .Y(_10202_));
 NAND2x1_ASAP7_75t_R _18395_ (.A(_01048_),
    .B(_10106_),
    .Y(_10203_));
 AO21x1_ASAP7_75t_R _18396_ (.A1(_10181_),
    .A2(_10203_),
    .B(net5540),
    .Y(_10204_));
 AOI21x1_ASAP7_75t_R _18397_ (.A1(_10202_),
    .A2(_10204_),
    .B(net6297),
    .Y(_10205_));
 OAI21x1_ASAP7_75t_R _18398_ (.A1(_10199_),
    .A2(_10205_),
    .B(net5558),
    .Y(_10206_));
 NOR2x1_ASAP7_75t_R _18399_ (.A(net5224),
    .B(net6291),
    .Y(_10207_));
 INVx1_ASAP7_75t_R _18400_ (.A(_01042_),
    .Y(_10208_));
 NAND2x1p5_ASAP7_75t_R _18401_ (.A(_10208_),
    .B(net6291),
    .Y(_10209_));
 INVx2_ASAP7_75t_R _18402_ (.A(_10209_),
    .Y(_10210_));
 OAI21x1_ASAP7_75t_R _18404_ (.A1(_10207_),
    .A2(_10210_),
    .B(net5935),
    .Y(_10212_));
 NOR2x1_ASAP7_75t_R _18405_ (.A(_10118_),
    .B(net6291),
    .Y(_10213_));
 OAI21x1_ASAP7_75t_R _18407_ (.A1(net4961),
    .A2(_10144_),
    .B(net5540),
    .Y(_10215_));
 AOI21x1_ASAP7_75t_R _18408_ (.A1(_10212_),
    .A2(_10215_),
    .B(net6297),
    .Y(_10216_));
 NOR2x1p5_ASAP7_75t_R _18409_ (.A(net6291),
    .B(_10208_),
    .Y(_10217_));
 NAND2x1_ASAP7_75t_R _18410_ (.A(net5935),
    .B(_10217_),
    .Y(_10218_));
 NOR2x1_ASAP7_75t_R _18411_ (.A(net6291),
    .B(net5940),
    .Y(_10219_));
 OAI21x1_ASAP7_75t_R _18413_ (.A1(_10210_),
    .A2(_10219_),
    .B(net5540),
    .Y(_10221_));
 AOI21x1_ASAP7_75t_R _18414_ (.A1(_10218_),
    .A2(_10221_),
    .B(net5914),
    .Y(_10222_));
 OAI21x1_ASAP7_75t_R _18415_ (.A1(_10216_),
    .A2(_10222_),
    .B(net5933),
    .Y(_10223_));
 AOI21x1_ASAP7_75t_R _18416_ (.A1(_10206_),
    .A2(_10223_),
    .B(net5932),
    .Y(_10224_));
 INVx2_ASAP7_75t_R _18418_ (.A(_10155_),
    .Y(_10226_));
 INVx1_ASAP7_75t_R _18420_ (.A(_01043_),
    .Y(_10228_));
 AO21x1_ASAP7_75t_R _18421_ (.A1(net6298),
    .A2(net6388),
    .B(_10228_),
    .Y(_10229_));
 NAND2x1_ASAP7_75t_R _18422_ (.A(net5936),
    .B(_10229_),
    .Y(_10230_));
 NAND2x1_ASAP7_75t_R _18423_ (.A(net6302),
    .B(net6288),
    .Y(_10231_));
 AOI21x1_ASAP7_75t_R _18424_ (.A1(net6388),
    .A2(net6298),
    .B(net5565),
    .Y(_10232_));
 NOR2x1_ASAP7_75t_R _18425_ (.A(net5937),
    .B(_10232_),
    .Y(_10233_));
 NAND2x1_ASAP7_75t_R _18426_ (.A(_10231_),
    .B(_10233_),
    .Y(_10234_));
 OAI21x1_ASAP7_75t_R _18427_ (.A1(net5017),
    .A2(_10230_),
    .B(_10234_),
    .Y(_10235_));
 INVx1_ASAP7_75t_R _18428_ (.A(_01045_),
    .Y(_10236_));
 AO21x1_ASAP7_75t_R _18429_ (.A1(net6298),
    .A2(net6388),
    .B(_10236_),
    .Y(_10237_));
 INVx1_ASAP7_75t_R _18430_ (.A(_01046_),
    .Y(_10238_));
 NAND2x1_ASAP7_75t_R _18431_ (.A(_10238_),
    .B(net6289),
    .Y(_10239_));
 AO21x1_ASAP7_75t_R _18432_ (.A1(_10237_),
    .A2(_10239_),
    .B(net5541),
    .Y(_10240_));
 NOR2x1_ASAP7_75t_R _18433_ (.A(net6287),
    .B(net6289),
    .Y(_10241_));
 OA21x2_ASAP7_75t_R _18435_ (.A1(_10241_),
    .A2(net5936),
    .B(net5916),
    .Y(_10243_));
 AOI21x1_ASAP7_75t_R _18436_ (.A1(_10240_),
    .A2(_10243_),
    .B(net5933),
    .Y(_10244_));
 OAI21x1_ASAP7_75t_R _18437_ (.A1(net5912),
    .A2(_10235_),
    .B(_10244_),
    .Y(_10245_));
 NOR2x1_ASAP7_75t_R _18438_ (.A(net6292),
    .B(net6300),
    .Y(_10246_));
 OAI21x1_ASAP7_75t_R _18440_ (.A1(_10246_),
    .A2(_10123_),
    .B(net5541),
    .Y(_10248_));
 NAND2x1_ASAP7_75t_R _18441_ (.A(_10248_),
    .B(_10166_),
    .Y(_10249_));
 NAND2x1_ASAP7_75t_R _18442_ (.A(_10228_),
    .B(net6289),
    .Y(_10250_));
 AO21x1_ASAP7_75t_R _18443_ (.A1(_10164_),
    .A2(_10250_),
    .B(net5541),
    .Y(_10251_));
 INVx1_ASAP7_75t_R _18444_ (.A(_10232_),
    .Y(_10252_));
 AOI21x1_ASAP7_75t_R _18445_ (.A1(net6288),
    .A2(net5941),
    .B(net5937),
    .Y(_10253_));
 AOI21x1_ASAP7_75t_R _18446_ (.A1(_10252_),
    .A2(_10253_),
    .B(net5911),
    .Y(_10254_));
 AOI21x1_ASAP7_75t_R _18447_ (.A1(_10251_),
    .A2(_10254_),
    .B(net5558),
    .Y(_10255_));
 OAI21x1_ASAP7_75t_R _18448_ (.A1(net6297),
    .A2(_10249_),
    .B(_10255_),
    .Y(_10256_));
 AOI21x1_ASAP7_75t_R _18450_ (.A1(_10245_),
    .A2(_10256_),
    .B(net5536),
    .Y(_10258_));
 OAI21x1_ASAP7_75t_R _18451_ (.A1(_10224_),
    .A2(_10258_),
    .B(_10189_),
    .Y(_10259_));
 NAND2x1_ASAP7_75t_R _18452_ (.A(_10191_),
    .B(_10259_),
    .Y(_00024_));
 NAND2x1_ASAP7_75t_R _18454_ (.A(net5937),
    .B(net5538),
    .Y(_10261_));
 AO21x1_ASAP7_75t_R _18455_ (.A1(net5538),
    .A2(net5223),
    .B(net5937),
    .Y(_10262_));
 OA21x2_ASAP7_75t_R _18456_ (.A1(net5017),
    .A2(_10261_),
    .B(_10262_),
    .Y(_10263_));
 NOR2x1_ASAP7_75t_R _18457_ (.A(net5540),
    .B(_10237_),
    .Y(_10264_));
 NOR2x1_ASAP7_75t_R _18458_ (.A(net6297),
    .B(_10264_),
    .Y(_10265_));
 NAND2x1_ASAP7_75t_R _18459_ (.A(_10196_),
    .B(_10176_),
    .Y(_10266_));
 AO21x1_ASAP7_75t_R _18461_ (.A1(_10265_),
    .A2(_10266_),
    .B(net5933),
    .Y(_10268_));
 AOI21x1_ASAP7_75t_R _18462_ (.A1(net6297),
    .A2(_10263_),
    .B(_10268_),
    .Y(_10269_));
 OA21x2_ASAP7_75t_R _18463_ (.A1(_10157_),
    .A2(net5936),
    .B(net6297),
    .Y(_10270_));
 NAND2x1_ASAP7_75t_R _18464_ (.A(_01057_),
    .B(net5937),
    .Y(_10271_));
 NOR2x1_ASAP7_75t_R _18465_ (.A(net6300),
    .B(net5938),
    .Y(_10272_));
 NAND2x1_ASAP7_75t_R _18466_ (.A(net5541),
    .B(_10272_),
    .Y(_10273_));
 AND3x1_ASAP7_75t_R _18467_ (.A(_10270_),
    .B(_10271_),
    .C(_10273_),
    .Y(_10274_));
 AO21x1_ASAP7_75t_R _18468_ (.A1(net5263),
    .A2(_10250_),
    .B(net5539),
    .Y(_10275_));
 AO21x1_ASAP7_75t_R _18469_ (.A1(_10157_),
    .A2(_10113_),
    .B(net5934),
    .Y(_10276_));
 NAND2x1_ASAP7_75t_R _18470_ (.A(_10275_),
    .B(_10276_),
    .Y(_10277_));
 OAI21x1_ASAP7_75t_R _18471_ (.A1(net6297),
    .A2(_10277_),
    .B(net5933),
    .Y(_10278_));
 OAI21x1_ASAP7_75t_R _18472_ (.A1(_10274_),
    .A2(_10278_),
    .B(net5536),
    .Y(_10279_));
 NOR2x1_ASAP7_75t_R _18473_ (.A(_10269_),
    .B(_10279_),
    .Y(_10280_));
 NAND2x1_ASAP7_75t_R _18474_ (.A(net6290),
    .B(net6300),
    .Y(_10281_));
 AO21x1_ASAP7_75t_R _18475_ (.A1(net6298),
    .A2(net6388),
    .B(net5566),
    .Y(_10282_));
 AO21x1_ASAP7_75t_R _18476_ (.A1(_10281_),
    .A2(_10282_),
    .B(net5541),
    .Y(_10283_));
 OA21x2_ASAP7_75t_R _18477_ (.A1(net5937),
    .A2(net5537),
    .B(_10283_),
    .Y(_10284_));
 OA21x2_ASAP7_75t_R _18478_ (.A1(net5567),
    .A2(net6290),
    .B(net5937),
    .Y(_10285_));
 NAND2x1_ASAP7_75t_R _18479_ (.A(net5018),
    .B(_10285_),
    .Y(_10286_));
 OA21x2_ASAP7_75t_R _18480_ (.A1(net5223),
    .A2(net5937),
    .B(net5917),
    .Y(_10287_));
 AO21x1_ASAP7_75t_R _18481_ (.A1(_10286_),
    .A2(_10287_),
    .B(net5933),
    .Y(_10288_));
 AOI21x1_ASAP7_75t_R _18482_ (.A1(net6297),
    .A2(_10284_),
    .B(_10288_),
    .Y(_10289_));
 AOI21x1_ASAP7_75t_R _18483_ (.A1(net6301),
    .A2(net6290),
    .B(net5937),
    .Y(_10290_));
 INVx1_ASAP7_75t_R _18484_ (.A(_10290_),
    .Y(_10291_));
 NOR2x1_ASAP7_75t_R _18485_ (.A(net5265),
    .B(_10291_),
    .Y(_10292_));
 NOR2x1_ASAP7_75t_R _18486_ (.A(net6301),
    .B(net6300),
    .Y(_10293_));
 OAI21x1_ASAP7_75t_R _18488_ (.A1(_10293_),
    .A2(_10261_),
    .B(net5913),
    .Y(_10295_));
 OAI21x1_ASAP7_75t_R _18490_ (.A1(_10292_),
    .A2(_10295_),
    .B(net5933),
    .Y(_10297_));
 OA21x2_ASAP7_75t_R _18491_ (.A1(_10143_),
    .A2(net5937),
    .B(net6297),
    .Y(_10298_));
 AO21x1_ASAP7_75t_R _18492_ (.A1(_10157_),
    .A2(_10155_),
    .B(net5541),
    .Y(_10299_));
 NAND2x1_ASAP7_75t_R _18493_ (.A(net5540),
    .B(_10142_),
    .Y(_10300_));
 AND3x1_ASAP7_75t_R _18494_ (.A(_10298_),
    .B(_10299_),
    .C(_10300_),
    .Y(_10301_));
 OAI21x1_ASAP7_75t_R _18495_ (.A1(_10297_),
    .A2(_10301_),
    .B(net5932),
    .Y(_10302_));
 OAI21x1_ASAP7_75t_R _18496_ (.A1(_10289_),
    .A2(_10302_),
    .B(net5557),
    .Y(_10303_));
 AO21x1_ASAP7_75t_R _18497_ (.A1(net5263),
    .A2(net5225),
    .B(net5541),
    .Y(_10304_));
 AO21x1_ASAP7_75t_R _18498_ (.A1(_10164_),
    .A2(net4964),
    .B(net5937),
    .Y(_10305_));
 AOI21x1_ASAP7_75t_R _18499_ (.A1(_10304_),
    .A2(_10305_),
    .B(net5917),
    .Y(_10306_));
 AO21x1_ASAP7_75t_R _18500_ (.A1(net6298),
    .A2(net6388),
    .B(_01050_),
    .Y(_10307_));
 NAND2x1_ASAP7_75t_R _18501_ (.A(_10307_),
    .B(_10197_),
    .Y(_10308_));
 NAND2x1_ASAP7_75t_R _18502_ (.A(net6299),
    .B(_09007_),
    .Y(_10309_));
 AO21x1_ASAP7_75t_R _18503_ (.A1(_10309_),
    .A2(_10239_),
    .B(net5541),
    .Y(_10310_));
 AOI21x1_ASAP7_75t_R _18505_ (.A1(_10308_),
    .A2(_10310_),
    .B(net6297),
    .Y(_10312_));
 OAI21x1_ASAP7_75t_R _18506_ (.A1(_10306_),
    .A2(_10312_),
    .B(net5558),
    .Y(_10313_));
 AO21x1_ASAP7_75t_R _18507_ (.A1(net6298),
    .A2(net6388),
    .B(net5310),
    .Y(_10314_));
 AO21x1_ASAP7_75t_R _18508_ (.A1(_10314_),
    .A2(_10250_),
    .B(net5937),
    .Y(_10315_));
 AOI21x1_ASAP7_75t_R _18509_ (.A1(net5018),
    .A2(_10285_),
    .B(net5917),
    .Y(_10316_));
 NAND2x1_ASAP7_75t_R _18510_ (.A(_10315_),
    .B(_10316_),
    .Y(_10317_));
 OA21x2_ASAP7_75t_R _18511_ (.A1(net5537),
    .A2(net5937),
    .B(net5916),
    .Y(_10318_));
 AND2x2_ASAP7_75t_R _18512_ (.A(_10164_),
    .B(_10156_),
    .Y(_10319_));
 AOI21x1_ASAP7_75t_R _18514_ (.A1(_10318_),
    .A2(_10319_),
    .B(net5558),
    .Y(_10321_));
 AOI21x1_ASAP7_75t_R _18515_ (.A1(_10317_),
    .A2(_10321_),
    .B(net5536),
    .Y(_10322_));
 NAND2x1_ASAP7_75t_R _18516_ (.A(_10313_),
    .B(_10322_),
    .Y(_10323_));
 NAND2x1_ASAP7_75t_R _18517_ (.A(_01059_),
    .B(net5935),
    .Y(_10324_));
 INVx1_ASAP7_75t_R _18518_ (.A(_10165_),
    .Y(_10325_));
 OAI21x1_ASAP7_75t_R _18520_ (.A1(_10213_),
    .A2(_10325_),
    .B(net5540),
    .Y(_10327_));
 OAI21x1_ASAP7_75t_R _18521_ (.A1(net5558),
    .A2(_10324_),
    .B(_10327_),
    .Y(_10328_));
 AOI21x1_ASAP7_75t_R _18522_ (.A1(net5917),
    .A2(_10328_),
    .B(net5932),
    .Y(_10329_));
 NAND2x1_ASAP7_75t_R _18523_ (.A(_10309_),
    .B(_10197_),
    .Y(_10330_));
 NOR2x1_ASAP7_75t_R _18524_ (.A(net5541),
    .B(_10246_),
    .Y(_10331_));
 AOI21x1_ASAP7_75t_R _18525_ (.A1(_10184_),
    .A2(_10331_),
    .B(net5558),
    .Y(_10332_));
 NAND2x1_ASAP7_75t_R _18526_ (.A(_10330_),
    .B(_10332_),
    .Y(_10333_));
 AOI21x1_ASAP7_75t_R _18527_ (.A1(net5935),
    .A2(_10325_),
    .B(net5933),
    .Y(_10334_));
 AOI21x1_ASAP7_75t_R _18528_ (.A1(_10307_),
    .A2(_10290_),
    .B(_10264_),
    .Y(_10335_));
 AOI21x1_ASAP7_75t_R _18530_ (.A1(_10334_),
    .A2(_10335_),
    .B(net5913),
    .Y(_10337_));
 NAND2x1_ASAP7_75t_R _18531_ (.A(_10333_),
    .B(_10337_),
    .Y(_10338_));
 AOI21x1_ASAP7_75t_R _18532_ (.A1(_10329_),
    .A2(_10338_),
    .B(net5557),
    .Y(_10339_));
 NAND2x1_ASAP7_75t_R _18533_ (.A(_10323_),
    .B(_10339_),
    .Y(_10340_));
 OAI21x1_ASAP7_75t_R _18534_ (.A1(_10280_),
    .A2(_10303_),
    .B(_10340_),
    .Y(_00025_));
 AO21x1_ASAP7_75t_R _18535_ (.A1(_10282_),
    .A2(_10239_),
    .B(net5934),
    .Y(_10341_));
 NOR2x1_ASAP7_75t_R _18536_ (.A(_10232_),
    .B(_10126_),
    .Y(_10342_));
 NAND2x1_ASAP7_75t_R _18537_ (.A(_10281_),
    .B(_10342_),
    .Y(_10343_));
 AO21x1_ASAP7_75t_R _18538_ (.A1(_10341_),
    .A2(_10343_),
    .B(net5915),
    .Y(_10344_));
 AND2x2_ASAP7_75t_R _18539_ (.A(_10176_),
    .B(net5263),
    .Y(_10345_));
 NAND2x1_ASAP7_75t_R _18540_ (.A(net5534),
    .B(net6289),
    .Y(_10346_));
 AO21x1_ASAP7_75t_R _18541_ (.A1(net6298),
    .A2(net6388),
    .B(_10238_),
    .Y(_10347_));
 AOI21x1_ASAP7_75t_R _18542_ (.A1(_10346_),
    .A2(_10347_),
    .B(net5539),
    .Y(_10348_));
 OR3x1_ASAP7_75t_R _18543_ (.A(_10345_),
    .B(net6297),
    .C(_10348_),
    .Y(_10349_));
 NAND2x1_ASAP7_75t_R _18544_ (.A(_10344_),
    .B(_10349_),
    .Y(_10350_));
 OAI21x1_ASAP7_75t_R _18545_ (.A1(_10219_),
    .A2(_10226_),
    .B(net5540),
    .Y(_10351_));
 NAND2x1_ASAP7_75t_R _18546_ (.A(net5937),
    .B(_10171_),
    .Y(_10352_));
 INVx1_ASAP7_75t_R _18547_ (.A(_10352_),
    .Y(_10353_));
 NAND2x1_ASAP7_75t_R _18548_ (.A(_10314_),
    .B(_10353_),
    .Y(_10354_));
 AOI21x1_ASAP7_75t_R _18549_ (.A1(_10354_),
    .A2(_10351_),
    .B(net5916),
    .Y(_10355_));
 INVx1_ASAP7_75t_R _18550_ (.A(net5567),
    .Y(_10356_));
 NOR2x1_ASAP7_75t_R _18551_ (.A(_10356_),
    .B(net6289),
    .Y(_10357_));
 INVx1_ASAP7_75t_R _18552_ (.A(_10357_),
    .Y(_10358_));
 AO21x1_ASAP7_75t_R _18553_ (.A1(_10358_),
    .A2(_10250_),
    .B(net5539),
    .Y(_10359_));
 NOR2x1_ASAP7_75t_R _18554_ (.A(net6297),
    .B(_10233_),
    .Y(_10360_));
 AO21x1_ASAP7_75t_R _18555_ (.A1(_10359_),
    .A2(_10360_),
    .B(net5933),
    .Y(_10361_));
 OAI21x1_ASAP7_75t_R _18556_ (.A1(_10361_),
    .A2(_10355_),
    .B(net5536),
    .Y(_10362_));
 AOI21x1_ASAP7_75t_R _18557_ (.A1(net5933),
    .A2(_10350_),
    .B(_10362_),
    .Y(_10363_));
 AOI21x1_ASAP7_75t_R _18558_ (.A1(_10282_),
    .A2(net5535),
    .B(_10140_),
    .Y(_10364_));
 NAND2x1_ASAP7_75t_R _18559_ (.A(net4962),
    .B(_10331_),
    .Y(_10365_));
 NAND2x1_ASAP7_75t_R _18560_ (.A(_10364_),
    .B(_10365_),
    .Y(_10366_));
 NOR2x1p5_ASAP7_75t_R _18561_ (.A(net5265),
    .B(_10156_),
    .Y(_10367_));
 NOR2x1_ASAP7_75t_R _18562_ (.A(net4963),
    .B(_10291_),
    .Y(_10368_));
 OAI21x1_ASAP7_75t_R _18563_ (.A1(_10367_),
    .A2(_10368_),
    .B(_10140_),
    .Y(_10369_));
 AOI21x1_ASAP7_75t_R _18564_ (.A1(_10366_),
    .A2(_10369_),
    .B(net5933),
    .Y(_10370_));
 AO21x1_ASAP7_75t_R _18565_ (.A1(_10281_),
    .A2(_10157_),
    .B(net5541),
    .Y(_10371_));
 AND3x1_ASAP7_75t_R _18566_ (.A(_10371_),
    .B(net5917),
    .C(_10159_),
    .Y(_10372_));
 OA21x2_ASAP7_75t_R _18567_ (.A1(_10282_),
    .A2(net5937),
    .B(net6297),
    .Y(_10373_));
 AO21x1_ASAP7_75t_R _18568_ (.A1(_10171_),
    .A2(_10157_),
    .B(net5541),
    .Y(_10374_));
 INVx1_ASAP7_75t_R _18569_ (.A(_10158_),
    .Y(_10375_));
 NAND2x1_ASAP7_75t_R _18570_ (.A(net5541),
    .B(net4710),
    .Y(_10376_));
 AO31x2_ASAP7_75t_R _18571_ (.A1(_10373_),
    .A2(_10374_),
    .A3(_10376_),
    .B(net5558),
    .Y(_10377_));
 OAI21x1_ASAP7_75t_R _18572_ (.A1(_10372_),
    .A2(_10377_),
    .B(net5932),
    .Y(_10378_));
 OAI21x1_ASAP7_75t_R _18573_ (.A1(_10370_),
    .A2(_10378_),
    .B(_10189_),
    .Y(_10379_));
 AO21x1_ASAP7_75t_R _18574_ (.A1(net5263),
    .A2(_10203_),
    .B(net5540),
    .Y(_10380_));
 NAND2x1_ASAP7_75t_R _18575_ (.A(_10307_),
    .B(_10253_),
    .Y(_10381_));
 AO21x1_ASAP7_75t_R _18576_ (.A1(_10380_),
    .A2(_10381_),
    .B(net5911),
    .Y(_10382_));
 OAI21x1_ASAP7_75t_R _18577_ (.A1(_10293_),
    .A2(_10219_),
    .B(net5935),
    .Y(_10383_));
 NAND2x1_ASAP7_75t_R _18578_ (.A(_01059_),
    .B(net5540),
    .Y(_10384_));
 AO21x1_ASAP7_75t_R _18579_ (.A1(_10383_),
    .A2(_10384_),
    .B(net6297),
    .Y(_10385_));
 AOI21x1_ASAP7_75t_R _18580_ (.A1(_10382_),
    .A2(_10385_),
    .B(net5558),
    .Y(_10386_));
 OA21x2_ASAP7_75t_R _18581_ (.A1(_01055_),
    .A2(net5934),
    .B(net5911),
    .Y(_10387_));
 AO21x1_ASAP7_75t_R _18582_ (.A1(net5262),
    .A2(_10113_),
    .B(net5539),
    .Y(_10388_));
 AOI21x1_ASAP7_75t_R _18583_ (.A1(_10387_),
    .A2(_10388_),
    .B(net5933),
    .Y(_10389_));
 AOI21x1_ASAP7_75t_R _18584_ (.A1(net5262),
    .A2(_10176_),
    .B(net5916),
    .Y(_10390_));
 AO21x1_ASAP7_75t_R _18585_ (.A1(_10309_),
    .A2(_10171_),
    .B(net5539),
    .Y(_10391_));
 NAND2x1_ASAP7_75t_R _18586_ (.A(_10390_),
    .B(_10391_),
    .Y(_10392_));
 AO21x1_ASAP7_75t_R _18587_ (.A1(_10389_),
    .A2(_10392_),
    .B(net5536),
    .Y(_10393_));
 OA21x2_ASAP7_75t_R _18588_ (.A1(_01058_),
    .A2(net5934),
    .B(net6297),
    .Y(_10394_));
 NAND2x1_ASAP7_75t_R _18589_ (.A(_10394_),
    .B(_10343_),
    .Y(_10395_));
 NAND2x1_ASAP7_75t_R _18590_ (.A(_01053_),
    .B(net5934),
    .Y(_10396_));
 AOI21x1_ASAP7_75t_R _18591_ (.A1(_10396_),
    .A2(_10360_),
    .B(net5558),
    .Y(_10397_));
 AOI21x1_ASAP7_75t_R _18592_ (.A1(_10395_),
    .A2(_10397_),
    .B(net5932),
    .Y(_10398_));
 INVx1_ASAP7_75t_R _18593_ (.A(_10285_),
    .Y(_10399_));
 OAI21x1_ASAP7_75t_R _18594_ (.A1(_10193_),
    .A2(_10399_),
    .B(_10327_),
    .Y(_10400_));
 AO21x1_ASAP7_75t_R _18595_ (.A1(_10157_),
    .A2(_10209_),
    .B(net5541),
    .Y(_10401_));
 OA21x2_ASAP7_75t_R _18596_ (.A1(net5225),
    .A2(net5936),
    .B(net5917),
    .Y(_10402_));
 AOI21x1_ASAP7_75t_R _18597_ (.A1(_10401_),
    .A2(_10402_),
    .B(net5933),
    .Y(_10403_));
 OAI21x1_ASAP7_75t_R _18598_ (.A1(net5917),
    .A2(_10400_),
    .B(_10403_),
    .Y(_10404_));
 AOI21x1_ASAP7_75t_R _18599_ (.A1(_10398_),
    .A2(_10404_),
    .B(_10189_),
    .Y(_10405_));
 OAI21x1_ASAP7_75t_R _18600_ (.A1(_10386_),
    .A2(_10393_),
    .B(_10405_),
    .Y(_10406_));
 OAI21x1_ASAP7_75t_R _18601_ (.A1(_10379_),
    .A2(_10363_),
    .B(_10406_),
    .Y(_00026_));
 NOR2x1_ASAP7_75t_R _18602_ (.A(net5311),
    .B(net6290),
    .Y(_10407_));
 INVx1_ASAP7_75t_R _18603_ (.A(_10231_),
    .Y(_10408_));
 OAI21x1_ASAP7_75t_R _18604_ (.A1(_10407_),
    .A2(_10408_),
    .B(net5937),
    .Y(_10409_));
 AOI21x1_ASAP7_75t_R _18605_ (.A1(_10327_),
    .A2(_10409_),
    .B(net6297),
    .Y(_10410_));
 OAI21x1_ASAP7_75t_R _18606_ (.A1(_10364_),
    .A2(_10410_),
    .B(net5933),
    .Y(_10411_));
 NAND2x1_ASAP7_75t_R _18607_ (.A(_10229_),
    .B(_10201_),
    .Y(_10412_));
 OAI21x1_ASAP7_75t_R _18608_ (.A1(_10241_),
    .A2(_10375_),
    .B(net5936),
    .Y(_10413_));
 AOI21x1_ASAP7_75t_R _18609_ (.A1(_10412_),
    .A2(_10413_),
    .B(net5912),
    .Y(_10414_));
 AOI21x1_ASAP7_75t_R _18610_ (.A1(_10266_),
    .A2(_10145_),
    .B(net6297),
    .Y(_10415_));
 OAI21x1_ASAP7_75t_R _18611_ (.A1(_10414_),
    .A2(_10415_),
    .B(net5558),
    .Y(_10416_));
 AOI21x1_ASAP7_75t_R _18612_ (.A1(_10411_),
    .A2(_10416_),
    .B(net5536),
    .Y(_10417_));
 AOI21x1_ASAP7_75t_R _18613_ (.A1(net5936),
    .A2(net4710),
    .B(net5933),
    .Y(_10418_));
 OAI21x1_ASAP7_75t_R _18614_ (.A1(net4963),
    .A2(_10291_),
    .B(_10418_),
    .Y(_10419_));
 AOI21x1_ASAP7_75t_R _18615_ (.A1(net5538),
    .A2(_10201_),
    .B(net5558),
    .Y(_10420_));
 OAI21x1_ASAP7_75t_R _18616_ (.A1(_10193_),
    .A2(_10230_),
    .B(_10420_),
    .Y(_10421_));
 NAND2x1_ASAP7_75t_R _18617_ (.A(_10419_),
    .B(_10421_),
    .Y(_10422_));
 OAI21x1_ASAP7_75t_R _18618_ (.A1(net4961),
    .A2(_10272_),
    .B(net5540),
    .Y(_10423_));
 AOI21x1_ASAP7_75t_R _18619_ (.A1(_10218_),
    .A2(_10423_),
    .B(net5558),
    .Y(_10424_));
 NAND2x1p5_ASAP7_75t_R _18620_ (.A(_10226_),
    .B(net5540),
    .Y(_10425_));
 OA21x2_ASAP7_75t_R _18621_ (.A1(net4964),
    .A2(net5540),
    .B(net6297),
    .Y(_10426_));
 OAI21x1_ASAP7_75t_R _18622_ (.A1(net5933),
    .A2(_10425_),
    .B(_10426_),
    .Y(_10427_));
 OAI21x1_ASAP7_75t_R _18623_ (.A1(_10424_),
    .A2(_10427_),
    .B(net5536),
    .Y(_10428_));
 AOI21x1_ASAP7_75t_R _18624_ (.A1(net5917),
    .A2(_10422_),
    .B(_10428_),
    .Y(_10429_));
 OAI21x1_ASAP7_75t_R _18625_ (.A1(_10417_),
    .A2(_10429_),
    .B(_10189_),
    .Y(_10430_));
 OAI21x1_ASAP7_75t_R _18626_ (.A1(_10142_),
    .A2(_10192_),
    .B(net5540),
    .Y(_10431_));
 OAI21x1_ASAP7_75t_R _18627_ (.A1(_10156_),
    .A2(_10246_),
    .B(_10431_),
    .Y(_10432_));
 NAND2x1_ASAP7_75t_R _18628_ (.A(_09007_),
    .B(net5940),
    .Y(_10433_));
 NAND2x1_ASAP7_75t_R _18629_ (.A(_10433_),
    .B(_10290_),
    .Y(_10434_));
 INVx2_ASAP7_75t_R _18630_ (.A(_10217_),
    .Y(_10435_));
 AOI21x1_ASAP7_75t_R _18631_ (.A1(net5935),
    .A2(_10435_),
    .B(net5916),
    .Y(_10436_));
 AOI21x1_ASAP7_75t_R _18632_ (.A1(_10434_),
    .A2(_10436_),
    .B(net5558),
    .Y(_10437_));
 OAI21x1_ASAP7_75t_R _18633_ (.A1(net6297),
    .A2(_10432_),
    .B(_10437_),
    .Y(_10438_));
 OAI21x1_ASAP7_75t_R _18634_ (.A1(_10217_),
    .A2(_10144_),
    .B(net5935),
    .Y(_10439_));
 INVx1_ASAP7_75t_R _18635_ (.A(_10203_),
    .Y(_10440_));
 OAI21x1_ASAP7_75t_R _18636_ (.A1(_10142_),
    .A2(_10440_),
    .B(net5540),
    .Y(_10441_));
 AOI21x1_ASAP7_75t_R _18637_ (.A1(_10439_),
    .A2(_10441_),
    .B(net5914),
    .Y(_10442_));
 AO21x1_ASAP7_75t_R _18638_ (.A1(_10157_),
    .A2(_10250_),
    .B(net5540),
    .Y(_10443_));
 AOI21x1_ASAP7_75t_R _18639_ (.A1(_10443_),
    .A2(_10351_),
    .B(net6297),
    .Y(_10444_));
 OAI21x1_ASAP7_75t_R _18640_ (.A1(_10442_),
    .A2(_10444_),
    .B(net5558),
    .Y(_10445_));
 AOI21x1_ASAP7_75t_R _18641_ (.A1(_10438_),
    .A2(_10445_),
    .B(net5932),
    .Y(_10446_));
 OAI21x1_ASAP7_75t_R _18642_ (.A1(net4961),
    .A2(_10226_),
    .B(net5540),
    .Y(_10447_));
 NAND2x1_ASAP7_75t_R _18643_ (.A(net6301),
    .B(net6300),
    .Y(_10448_));
 INVx1_ASAP7_75t_R _18644_ (.A(_10448_),
    .Y(_10449_));
 OAI21x1_ASAP7_75t_R _18645_ (.A1(_10142_),
    .A2(_10449_),
    .B(net5935),
    .Y(_10450_));
 AOI21x1_ASAP7_75t_R _18646_ (.A1(_10447_),
    .A2(_10450_),
    .B(net5914),
    .Y(_10451_));
 AO21x1_ASAP7_75t_R _18647_ (.A1(net5263),
    .A2(net5537),
    .B(net5935),
    .Y(_10452_));
 AO21x1_ASAP7_75t_R _18648_ (.A1(_10237_),
    .A2(_10203_),
    .B(net5540),
    .Y(_10453_));
 AOI21x1_ASAP7_75t_R _18649_ (.A1(_10452_),
    .A2(_10453_),
    .B(net6297),
    .Y(_10454_));
 OAI21x1_ASAP7_75t_R _18650_ (.A1(_10451_),
    .A2(_10454_),
    .B(net5558),
    .Y(_10455_));
 INVx1_ASAP7_75t_R _18651_ (.A(_10342_),
    .Y(_10456_));
 AOI21x1_ASAP7_75t_R _18652_ (.A1(_10456_),
    .A2(_10431_),
    .B(net6297),
    .Y(_10457_));
 OAI21x1_ASAP7_75t_R _18653_ (.A1(_10407_),
    .A2(_10226_),
    .B(net5540),
    .Y(_10458_));
 AOI21x1_ASAP7_75t_R _18654_ (.A1(_10458_),
    .A2(_10283_),
    .B(net5913),
    .Y(_10459_));
 OAI21x1_ASAP7_75t_R _18655_ (.A1(_10457_),
    .A2(_10459_),
    .B(net5933),
    .Y(_10460_));
 AOI21x1_ASAP7_75t_R _18656_ (.A1(_10455_),
    .A2(_10460_),
    .B(net5536),
    .Y(_10461_));
 OAI21x1_ASAP7_75t_R _18657_ (.A1(_10446_),
    .A2(_10461_),
    .B(net5557),
    .Y(_10462_));
 NAND2x1_ASAP7_75t_R _18658_ (.A(_10430_),
    .B(_10462_),
    .Y(_00027_));
 NOR2x1_ASAP7_75t_R _18659_ (.A(net6289),
    .B(net5541),
    .Y(_10463_));
 AO21x1_ASAP7_75t_R _18660_ (.A1(net5535),
    .A2(_10229_),
    .B(_10463_),
    .Y(_10464_));
 OAI21x1_ASAP7_75t_R _18661_ (.A1(net6297),
    .A2(_10464_),
    .B(net5933),
    .Y(_10465_));
 NAND2x1_ASAP7_75t_R _18662_ (.A(net5541),
    .B(_10246_),
    .Y(_10466_));
 AND3x1_ASAP7_75t_R _18663_ (.A(_10310_),
    .B(_10466_),
    .C(_10298_),
    .Y(_10467_));
 NOR2x1_ASAP7_75t_R _18664_ (.A(_10465_),
    .B(_10467_),
    .Y(_10468_));
 NOR2x1_ASAP7_75t_R _18665_ (.A(net5917),
    .B(_10285_),
    .Y(_10469_));
 AO21x1_ASAP7_75t_R _18666_ (.A1(net5938),
    .A2(net5310),
    .B(net5937),
    .Y(_10470_));
 AO21x1_ASAP7_75t_R _18667_ (.A1(_10469_),
    .A2(_10470_),
    .B(net5933),
    .Y(_10471_));
 AO21x1_ASAP7_75t_R _18668_ (.A1(_10435_),
    .A2(net5223),
    .B(net5937),
    .Y(_10472_));
 AND3x1_ASAP7_75t_R _18669_ (.A(_10472_),
    .B(net5917),
    .C(_10166_),
    .Y(_10473_));
 OAI21x1_ASAP7_75t_R _18670_ (.A1(_10471_),
    .A2(_10473_),
    .B(net5932),
    .Y(_10474_));
 NOR2x1_ASAP7_75t_R _18671_ (.A(_10468_),
    .B(_10474_),
    .Y(_10475_));
 NAND2x1_ASAP7_75t_R _18672_ (.A(_10356_),
    .B(net5541),
    .Y(_10476_));
 OAI21x1_ASAP7_75t_R _18673_ (.A1(net5541),
    .A2(net5263),
    .B(_10476_),
    .Y(_10477_));
 INVx1_ASAP7_75t_R _18674_ (.A(_10281_),
    .Y(_10478_));
 OAI21x1_ASAP7_75t_R _18675_ (.A1(_10407_),
    .A2(_10478_),
    .B(net5936),
    .Y(_10479_));
 AOI221x1_ASAP7_75t_R _18676_ (.A1(_10140_),
    .A2(_10477_),
    .B1(_10479_),
    .B2(_10114_),
    .C(net5933),
    .Y(_10480_));
 AND3x1_ASAP7_75t_R _18677_ (.A(_10182_),
    .B(net5913),
    .C(_10195_),
    .Y(_10481_));
 INVx1_ASAP7_75t_R _18678_ (.A(_10409_),
    .Y(_10482_));
 NAND2x1_ASAP7_75t_R _18679_ (.A(_10448_),
    .B(_10433_),
    .Y(_10483_));
 OAI21x1_ASAP7_75t_R _18680_ (.A1(net5936),
    .A2(_10483_),
    .B(net6297),
    .Y(_10484_));
 OAI21x1_ASAP7_75t_R _18681_ (.A1(_10482_),
    .A2(_10484_),
    .B(net5933),
    .Y(_10485_));
 OAI21x1_ASAP7_75t_R _18682_ (.A1(_10481_),
    .A2(_10485_),
    .B(net5536),
    .Y(_10486_));
 OAI21x1_ASAP7_75t_R _18683_ (.A1(_10480_),
    .A2(_10486_),
    .B(_10189_),
    .Y(_10487_));
 AOI21x1_ASAP7_75t_R _18684_ (.A1(_10330_),
    .A2(_10383_),
    .B(net6297),
    .Y(_10488_));
 OAI21x1_ASAP7_75t_R _18685_ (.A1(_10246_),
    .A2(_10449_),
    .B(net5540),
    .Y(_10489_));
 AO21x1_ASAP7_75t_R _18686_ (.A1(_10281_),
    .A2(_10181_),
    .B(net5540),
    .Y(_10490_));
 AOI21x1_ASAP7_75t_R _18687_ (.A1(_10489_),
    .A2(_10490_),
    .B(net5914),
    .Y(_10491_));
 OAI21x1_ASAP7_75t_R _18688_ (.A1(_10488_),
    .A2(_10491_),
    .B(net5933),
    .Y(_10492_));
 AO21x1_ASAP7_75t_R _18689_ (.A1(net5311),
    .A2(net5938),
    .B(net5540),
    .Y(_10493_));
 NOR2x1_ASAP7_75t_R _18690_ (.A(net5916),
    .B(_10123_),
    .Y(_10494_));
 AOI21x1_ASAP7_75t_R _18691_ (.A1(_10493_),
    .A2(_10494_),
    .B(net5933),
    .Y(_10495_));
 AOI21x1_ASAP7_75t_R _18692_ (.A1(_10307_),
    .A2(_10290_),
    .B(net6297),
    .Y(_10496_));
 AO21x1_ASAP7_75t_R _18693_ (.A1(_10433_),
    .A2(_10171_),
    .B(net5540),
    .Y(_10497_));
 NAND2x1_ASAP7_75t_R _18694_ (.A(_10496_),
    .B(_10497_),
    .Y(_10498_));
 AOI21x1_ASAP7_75t_R _18695_ (.A1(_10495_),
    .A2(_10498_),
    .B(net5536),
    .Y(_10499_));
 AOI21x1_ASAP7_75t_R _18696_ (.A1(_10492_),
    .A2(_10499_),
    .B(_10189_),
    .Y(_10500_));
 AO21x1_ASAP7_75t_R _18697_ (.A1(_10309_),
    .A2(_10113_),
    .B(net5539),
    .Y(_10501_));
 AOI21x1_ASAP7_75t_R _18698_ (.A1(_10341_),
    .A2(_10501_),
    .B(net5915),
    .Y(_10502_));
 AO21x1_ASAP7_75t_R _18699_ (.A1(_10309_),
    .A2(net5226),
    .B(net5539),
    .Y(_10503_));
 AOI21x1_ASAP7_75t_R _18700_ (.A1(_10276_),
    .A2(_10503_),
    .B(net6297),
    .Y(_10504_));
 OAI21x1_ASAP7_75t_R _18701_ (.A1(_10502_),
    .A2(_10504_),
    .B(net5933),
    .Y(_10505_));
 AO21x1_ASAP7_75t_R _18702_ (.A1(_10147_),
    .A2(net5936),
    .B(_10140_),
    .Y(_10506_));
 NAND2x1_ASAP7_75t_R _18703_ (.A(net4962),
    .B(_10163_),
    .Y(_10507_));
 OR2x2_ASAP7_75t_R _18704_ (.A(_10506_),
    .B(_10507_),
    .Y(_10508_));
 AO21x1_ASAP7_75t_R _18705_ (.A1(net5263),
    .A2(_10250_),
    .B(net5934),
    .Y(_10509_));
 AOI21x1_ASAP7_75t_R _18706_ (.A1(_10509_),
    .A2(_10134_),
    .B(net5933),
    .Y(_10510_));
 AOI21x1_ASAP7_75t_R _18707_ (.A1(_10508_),
    .A2(_10510_),
    .B(net5932),
    .Y(_10511_));
 NAND2x1_ASAP7_75t_R _18708_ (.A(_10505_),
    .B(_10511_),
    .Y(_10512_));
 NAND2x1_ASAP7_75t_R _18709_ (.A(_10500_),
    .B(_10512_),
    .Y(_10513_));
 OAI21x1_ASAP7_75t_R _18710_ (.A1(_10475_),
    .A2(_10487_),
    .B(_10513_),
    .Y(_00028_));
 AO21x1_ASAP7_75t_R _18711_ (.A1(net5534),
    .A2(net6288),
    .B(net5937),
    .Y(_10514_));
 OAI21x1_ASAP7_75t_R _18712_ (.A1(net4963),
    .A2(_10514_),
    .B(net6297),
    .Y(_10515_));
 AOI21x1_ASAP7_75t_R _18713_ (.A1(_10347_),
    .A2(_10353_),
    .B(_10515_),
    .Y(_10516_));
 AO21x1_ASAP7_75t_R _18714_ (.A1(_10282_),
    .A2(_10239_),
    .B(net5541),
    .Y(_10517_));
 AND3x1_ASAP7_75t_R _18715_ (.A(_10517_),
    .B(net5912),
    .C(_10248_),
    .Y(_10518_));
 OAI21x1_ASAP7_75t_R _18716_ (.A1(_10516_),
    .A2(_10518_),
    .B(net5932),
    .Y(_10519_));
 NAND2x1_ASAP7_75t_R _18717_ (.A(net6287),
    .B(net6300),
    .Y(_10520_));
 AOI21x1_ASAP7_75t_R _18718_ (.A1(_10520_),
    .A2(_10138_),
    .B(net5937),
    .Y(_10521_));
 OA21x2_ASAP7_75t_R _18719_ (.A1(_10325_),
    .A2(net4961),
    .B(net5935),
    .Y(_10522_));
 OAI21x1_ASAP7_75t_R _18720_ (.A1(_10521_),
    .A2(_10522_),
    .B(net6297),
    .Y(_10523_));
 NOR2x1_ASAP7_75t_R _18721_ (.A(net5940),
    .B(net5540),
    .Y(_10524_));
 INVx1_ASAP7_75t_R _18722_ (.A(_10489_),
    .Y(_10525_));
 OAI21x1_ASAP7_75t_R _18723_ (.A1(_10524_),
    .A2(_10525_),
    .B(net5914),
    .Y(_10526_));
 NAND3x1_ASAP7_75t_R _18724_ (.A(_10523_),
    .B(_10526_),
    .C(net5536),
    .Y(_10527_));
 AOI21x1_ASAP7_75t_R _18725_ (.A1(_10519_),
    .A2(_10527_),
    .B(net5933),
    .Y(_10528_));
 NOR2x1_ASAP7_75t_R _18726_ (.A(net5534),
    .B(net6288),
    .Y(_10529_));
 AO21x1_ASAP7_75t_R _18727_ (.A1(_10184_),
    .A2(net5541),
    .B(_10529_),
    .Y(_10530_));
 OA21x2_ASAP7_75t_R _18728_ (.A1(_10530_),
    .A2(net5916),
    .B(net5932),
    .Y(_10531_));
 NOR2x1_ASAP7_75t_R _18729_ (.A(net6297),
    .B(_10201_),
    .Y(_10532_));
 NAND2x1_ASAP7_75t_R _18730_ (.A(_10532_),
    .B(_10413_),
    .Y(_10533_));
 AO21x1_ASAP7_75t_R _18731_ (.A1(_10531_),
    .A2(_10533_),
    .B(net5558),
    .Y(_10534_));
 AND3x1_ASAP7_75t_R _18732_ (.A(_10307_),
    .B(net5019),
    .C(net5936),
    .Y(_10535_));
 OAI21x1_ASAP7_75t_R _18733_ (.A1(net5934),
    .A2(_10282_),
    .B(_10140_),
    .Y(_10536_));
 NOR2x1_ASAP7_75t_R _18734_ (.A(_10478_),
    .B(_10470_),
    .Y(_10537_));
 OA21x2_ASAP7_75t_R _18735_ (.A1(_10537_),
    .A2(_10506_),
    .B(net5536),
    .Y(_10538_));
 OA21x2_ASAP7_75t_R _18736_ (.A1(_10535_),
    .A2(_10536_),
    .B(_10538_),
    .Y(_10539_));
 OAI21x1_ASAP7_75t_R _18737_ (.A1(_10534_),
    .A2(_10539_),
    .B(net5557),
    .Y(_10540_));
 AO21x1_ASAP7_75t_R _18738_ (.A1(_10171_),
    .A2(_10157_),
    .B(net5937),
    .Y(_10541_));
 AND3x1_ASAP7_75t_R _18739_ (.A(_10166_),
    .B(_10541_),
    .C(net5913),
    .Y(_10542_));
 NOR2x1_ASAP7_75t_R _18740_ (.A(net5540),
    .B(net4961),
    .Y(_10543_));
 AO21x1_ASAP7_75t_R _18741_ (.A1(net5540),
    .A2(net5537),
    .B(_10543_),
    .Y(_10544_));
 AO21x1_ASAP7_75t_R _18742_ (.A1(_10544_),
    .A2(_10373_),
    .B(net5558),
    .Y(_10545_));
 OA21x2_ASAP7_75t_R _18743_ (.A1(net6301),
    .A2(net5540),
    .B(net5916),
    .Y(_10546_));
 AOI21x1_ASAP7_75t_R _18744_ (.A1(_10198_),
    .A2(_10546_),
    .B(net5933),
    .Y(_10547_));
 AOI21x1_ASAP7_75t_R _18745_ (.A1(_10131_),
    .A2(_10253_),
    .B(net5911),
    .Y(_10548_));
 OAI21x1_ASAP7_75t_R _18746_ (.A1(net5017),
    .A2(_10456_),
    .B(_10548_),
    .Y(_10549_));
 AOI21x1_ASAP7_75t_R _18747_ (.A1(_10547_),
    .A2(_10549_),
    .B(net5536),
    .Y(_10550_));
 OAI21x1_ASAP7_75t_R _18748_ (.A1(_10542_),
    .A2(_10545_),
    .B(_10550_),
    .Y(_10551_));
 OA21x2_ASAP7_75t_R _18749_ (.A1(_10210_),
    .A2(net4961),
    .B(net5935),
    .Y(_10552_));
 NAND2x1p5_ASAP7_75t_R _18750_ (.A(_10425_),
    .B(_10373_),
    .Y(_10553_));
 NAND2x1_ASAP7_75t_R _18751_ (.A(net5227),
    .B(net5935),
    .Y(_10554_));
 OAI21x1_ASAP7_75t_R _18752_ (.A1(net5938),
    .A2(_10476_),
    .B(_10554_),
    .Y(_10555_));
 AOI21x1_ASAP7_75t_R _18753_ (.A1(net5914),
    .A2(_10555_),
    .B(net5558),
    .Y(_10556_));
 OAI21x1_ASAP7_75t_R _18754_ (.A1(_10552_),
    .A2(_10553_),
    .B(_10556_),
    .Y(_10557_));
 NAND2x1_ASAP7_75t_R _18755_ (.A(_10230_),
    .B(_10270_),
    .Y(_10558_));
 OA21x2_ASAP7_75t_R _18756_ (.A1(_10193_),
    .A2(net5540),
    .B(_10237_),
    .Y(_10559_));
 AOI21x1_ASAP7_75t_R _18757_ (.A1(_10318_),
    .A2(_10559_),
    .B(net5933),
    .Y(_10560_));
 AOI21x1_ASAP7_75t_R _18758_ (.A1(_10558_),
    .A2(_10560_),
    .B(net5932),
    .Y(_10561_));
 AOI21x1_ASAP7_75t_R _18759_ (.A1(_10561_),
    .A2(_10557_),
    .B(net5557),
    .Y(_10562_));
 NAND2x1_ASAP7_75t_R _18760_ (.A(_10562_),
    .B(_10551_),
    .Y(_10563_));
 OAI21x1_ASAP7_75t_R _18761_ (.A1(_10528_),
    .A2(_10540_),
    .B(_10563_),
    .Y(_00029_));
 AO21x1_ASAP7_75t_R _18762_ (.A1(_10138_),
    .A2(_10250_),
    .B(net5934),
    .Y(_10564_));
 AO21x1_ASAP7_75t_R _18763_ (.A1(_10448_),
    .A2(_10171_),
    .B(net5539),
    .Y(_10565_));
 AO21x1_ASAP7_75t_R _18764_ (.A1(_10564_),
    .A2(_10565_),
    .B(net5911),
    .Y(_10566_));
 OA21x2_ASAP7_75t_R _18765_ (.A1(_10272_),
    .A2(_10529_),
    .B(net5539),
    .Y(_10567_));
 AND3x1_ASAP7_75t_R _18766_ (.A(_10448_),
    .B(_10171_),
    .C(net5937),
    .Y(_10568_));
 OAI21x1_ASAP7_75t_R _18767_ (.A1(_10567_),
    .A2(_10568_),
    .B(net5911),
    .Y(_10569_));
 NAND3x1_ASAP7_75t_R _18768_ (.A(_10566_),
    .B(_10569_),
    .C(net5558),
    .Y(_10570_));
 OAI21x1_ASAP7_75t_R _18769_ (.A1(net5934),
    .A2(net5019),
    .B(_10413_),
    .Y(_10571_));
 AOI21x1_ASAP7_75t_R _18770_ (.A1(_10271_),
    .A2(_10234_),
    .B(net5911),
    .Y(_10572_));
 AOI21x1_ASAP7_75t_R _18771_ (.A1(net5911),
    .A2(_10571_),
    .B(_10572_),
    .Y(_10573_));
 AOI21x1_ASAP7_75t_R _18772_ (.A1(net5933),
    .A2(_10573_),
    .B(net5536),
    .Y(_10574_));
 OR2x2_ASAP7_75t_R _18773_ (.A(_01054_),
    .B(net5539),
    .Y(_10575_));
 NAND2x1_ASAP7_75t_R _18774_ (.A(_10131_),
    .B(_10253_),
    .Y(_10576_));
 AOI21x1_ASAP7_75t_R _18775_ (.A1(_10575_),
    .A2(_10576_),
    .B(net6297),
    .Y(_10577_));
 AOI21x1_ASAP7_75t_R _18776_ (.A1(net5019),
    .A2(_10229_),
    .B(net5541),
    .Y(_10578_));
 AO21x1_ASAP7_75t_R _18777_ (.A1(net5939),
    .A2(net6287),
    .B(net5934),
    .Y(_10579_));
 NAND2x1_ASAP7_75t_R _18778_ (.A(net6297),
    .B(_10579_),
    .Y(_10580_));
 OAI21x1_ASAP7_75t_R _18779_ (.A1(_10578_),
    .A2(_10580_),
    .B(net5558),
    .Y(_10581_));
 NOR2x1_ASAP7_75t_R _18780_ (.A(_10577_),
    .B(_10581_),
    .Y(_10582_));
 OAI21x1_ASAP7_75t_R _18781_ (.A1(net6297),
    .A2(_10348_),
    .B(net5933),
    .Y(_10583_));
 AO21x1_ASAP7_75t_R _18782_ (.A1(net5939),
    .A2(net5227),
    .B(net5934),
    .Y(_10584_));
 AOI21x1_ASAP7_75t_R _18783_ (.A1(_10584_),
    .A2(_10479_),
    .B(net5911),
    .Y(_10585_));
 OAI21x1_ASAP7_75t_R _18784_ (.A1(_10583_),
    .A2(_10585_),
    .B(net5536),
    .Y(_10586_));
 NOR2x1_ASAP7_75t_R _18785_ (.A(_10582_),
    .B(_10586_),
    .Y(_10587_));
 AOI21x1_ASAP7_75t_R _18786_ (.A1(_10570_),
    .A2(_10574_),
    .B(_10587_),
    .Y(_10588_));
 NAND2x1p5_ASAP7_75t_R _18787_ (.A(net5262),
    .B(net5535),
    .Y(_10589_));
 AND3x1_ASAP7_75t_R _18788_ (.A(_10413_),
    .B(_10589_),
    .C(net6297),
    .Y(_10590_));
 AO21x1_ASAP7_75t_R _18789_ (.A1(net5566),
    .A2(net6289),
    .B(net5934),
    .Y(_10591_));
 NOR2x1_ASAP7_75t_R _18790_ (.A(net4963),
    .B(_10591_),
    .Y(_10592_));
 NAND2x1_ASAP7_75t_R _18791_ (.A(net5934),
    .B(_10357_),
    .Y(_10593_));
 NAND3x1_ASAP7_75t_R _18792_ (.A(_10124_),
    .B(_10593_),
    .C(net5916),
    .Y(_10594_));
 OAI21x1_ASAP7_75t_R _18793_ (.A1(_10592_),
    .A2(_10594_),
    .B(net5933),
    .Y(_10595_));
 AO21x1_ASAP7_75t_R _18794_ (.A1(_10314_),
    .A2(net4962),
    .B(net5541),
    .Y(_10596_));
 AOI21x1_ASAP7_75t_R _18795_ (.A1(_10596_),
    .A2(_10298_),
    .B(net5933),
    .Y(_10597_));
 OA21x2_ASAP7_75t_R _18796_ (.A1(net6300),
    .A2(net5937),
    .B(net5911),
    .Y(_10598_));
 NAND2x1_ASAP7_75t_R _18797_ (.A(net6288),
    .B(net5941),
    .Y(_10599_));
 AO21x1_ASAP7_75t_R _18798_ (.A1(_10599_),
    .A2(_10520_),
    .B(net5539),
    .Y(_10600_));
 NAND2x1_ASAP7_75t_R _18799_ (.A(_10598_),
    .B(_10600_),
    .Y(_10601_));
 NAND2x1_ASAP7_75t_R _18800_ (.A(_10597_),
    .B(_10601_),
    .Y(_10602_));
 OAI21x1_ASAP7_75t_R _18801_ (.A1(_10590_),
    .A2(_10595_),
    .B(_10602_),
    .Y(_10603_));
 AOI21x1_ASAP7_75t_R _18802_ (.A1(net5262),
    .A2(net5535),
    .B(net6297),
    .Y(_10604_));
 AO21x1_ASAP7_75t_R _18803_ (.A1(_10138_),
    .A2(_10113_),
    .B(net5539),
    .Y(_10605_));
 NAND2x1_ASAP7_75t_R _18804_ (.A(_10604_),
    .B(_10605_),
    .Y(_10606_));
 OA21x2_ASAP7_75t_R _18805_ (.A1(_10119_),
    .A2(net5934),
    .B(net6297),
    .Y(_10607_));
 NAND2x1_ASAP7_75t_R _18806_ (.A(_10309_),
    .B(_10133_),
    .Y(_10608_));
 AOI21x1_ASAP7_75t_R _18807_ (.A1(_10607_),
    .A2(_10608_),
    .B(net5558),
    .Y(_10609_));
 NAND2x1_ASAP7_75t_R _18808_ (.A(_10606_),
    .B(_10609_),
    .Y(_10610_));
 NAND2x1_ASAP7_75t_R _18809_ (.A(_10233_),
    .B(net5264),
    .Y(_10611_));
 AND2x2_ASAP7_75t_R _18810_ (.A(_10396_),
    .B(net6297),
    .Y(_10612_));
 AOI21x1_ASAP7_75t_R _18811_ (.A1(_10612_),
    .A2(_10611_),
    .B(net5933),
    .Y(_10613_));
 AOI21x1_ASAP7_75t_R _18812_ (.A1(_10599_),
    .A2(_10342_),
    .B(net6297),
    .Y(_10614_));
 OAI21x1_ASAP7_75t_R _18813_ (.A1(_10210_),
    .A2(_10470_),
    .B(_10614_),
    .Y(_10615_));
 AOI21x1_ASAP7_75t_R _18814_ (.A1(_10615_),
    .A2(_10613_),
    .B(net5932),
    .Y(_10616_));
 AOI21x1_ASAP7_75t_R _18815_ (.A1(_10616_),
    .A2(_10610_),
    .B(_10189_),
    .Y(_10617_));
 OAI21x1_ASAP7_75t_R _18816_ (.A1(_10603_),
    .A2(net5536),
    .B(_10617_),
    .Y(_10618_));
 OAI21x1_ASAP7_75t_R _18817_ (.A1(net5557),
    .A2(_10588_),
    .B(_10618_),
    .Y(_00030_));
 OA21x2_ASAP7_75t_R _18818_ (.A1(net6287),
    .A2(net5937),
    .B(net6297),
    .Y(_10619_));
 NAND2x1_ASAP7_75t_R _18819_ (.A(_10619_),
    .B(_10497_),
    .Y(_10620_));
 NAND2x1_ASAP7_75t_R _18820_ (.A(_10200_),
    .B(_10253_),
    .Y(_10621_));
 AO21x1_ASAP7_75t_R _18821_ (.A1(_10383_),
    .A2(_10621_),
    .B(net6297),
    .Y(_10622_));
 AOI21x1_ASAP7_75t_R _18822_ (.A1(_10620_),
    .A2(_10622_),
    .B(net5933),
    .Y(_10623_));
 AO21x1_ASAP7_75t_R _18823_ (.A1(_10358_),
    .A2(net5264),
    .B(net5934),
    .Y(_10624_));
 NOR2x1_ASAP7_75t_R _18824_ (.A(net5916),
    .B(_10133_),
    .Y(_10625_));
 AOI21x1_ASAP7_75t_R _18825_ (.A1(net5935),
    .A2(_10325_),
    .B(net6297),
    .Y(_10626_));
 AO21x1_ASAP7_75t_R _18826_ (.A1(_10425_),
    .A2(_10626_),
    .B(net5558),
    .Y(_10627_));
 AOI21x1_ASAP7_75t_R _18827_ (.A1(_10624_),
    .A2(_10625_),
    .B(_10627_),
    .Y(_10628_));
 NOR3x1_ASAP7_75t_R _18828_ (.A(_10628_),
    .B(_10623_),
    .C(net5932),
    .Y(_10629_));
 OA21x2_ASAP7_75t_R _18829_ (.A1(net4963),
    .A2(_10591_),
    .B(_10391_),
    .Y(_10630_));
 NAND2x1_ASAP7_75t_R _18830_ (.A(net5538),
    .B(_10201_),
    .Y(_10631_));
 NAND2x1_ASAP7_75t_R _18831_ (.A(_10631_),
    .B(_10275_),
    .Y(_10632_));
 OAI21x1_ASAP7_75t_R _18832_ (.A1(net5915),
    .A2(_10632_),
    .B(net5933),
    .Y(_10633_));
 AOI21x1_ASAP7_75t_R _18833_ (.A1(net5915),
    .A2(_10630_),
    .B(_10633_),
    .Y(_10634_));
 AO21x1_ASAP7_75t_R _18834_ (.A1(_10164_),
    .A2(_10113_),
    .B(net5934),
    .Y(_10635_));
 OA21x2_ASAP7_75t_R _18835_ (.A1(net5226),
    .A2(net5539),
    .B(net6297),
    .Y(_10636_));
 AND3x1_ASAP7_75t_R _18836_ (.A(_10635_),
    .B(_10636_),
    .C(_10593_),
    .Y(_10637_));
 AND2x2_ASAP7_75t_R _18837_ (.A(_10591_),
    .B(net5916),
    .Y(_10638_));
 AO21x1_ASAP7_75t_R _18838_ (.A1(_10638_),
    .A2(_10479_),
    .B(net5933),
    .Y(_10639_));
 OAI21x1_ASAP7_75t_R _18839_ (.A1(_10637_),
    .A2(_10639_),
    .B(net5932),
    .Y(_10640_));
 OAI21x1_ASAP7_75t_R _18840_ (.A1(_10634_),
    .A2(_10640_),
    .B(_10189_),
    .Y(_10641_));
 NAND2x1_ASAP7_75t_R _18841_ (.A(_10200_),
    .B(_10176_),
    .Y(_10642_));
 AOI21x1_ASAP7_75t_R _18842_ (.A1(_10642_),
    .A2(_10409_),
    .B(net5911),
    .Y(_10643_));
 AO21x1_ASAP7_75t_R _18843_ (.A1(_10119_),
    .A2(net5264),
    .B(net5539),
    .Y(_10644_));
 AO21x1_ASAP7_75t_R _18844_ (.A1(_10358_),
    .A2(net5226),
    .B(net5934),
    .Y(_10645_));
 AOI21x1_ASAP7_75t_R _18845_ (.A1(_10644_),
    .A2(_10645_),
    .B(net6297),
    .Y(_10646_));
 OAI21x1_ASAP7_75t_R _18846_ (.A1(_10643_),
    .A2(_10646_),
    .B(net5558),
    .Y(_10647_));
 OA21x2_ASAP7_75t_R _18847_ (.A1(_10314_),
    .A2(net5936),
    .B(net5226),
    .Y(_10648_));
 AOI21x1_ASAP7_75t_R _18848_ (.A1(net5941),
    .A2(_10463_),
    .B(net6297),
    .Y(_10649_));
 NAND2x1_ASAP7_75t_R _18849_ (.A(_10648_),
    .B(_10649_),
    .Y(_10650_));
 OA21x2_ASAP7_75t_R _18850_ (.A1(_01046_),
    .A2(net5937),
    .B(net6297),
    .Y(_10651_));
 AOI21x1_ASAP7_75t_R _18851_ (.A1(_10651_),
    .A2(_10600_),
    .B(net5558),
    .Y(_10652_));
 AOI21x1_ASAP7_75t_R _18852_ (.A1(_10650_),
    .A2(_10652_),
    .B(net5536),
    .Y(_10653_));
 NAND2x1_ASAP7_75t_R _18853_ (.A(_10647_),
    .B(_10653_),
    .Y(_10654_));
 INVx1_ASAP7_75t_R _18854_ (.A(_10310_),
    .Y(_10655_));
 NAND2x1_ASAP7_75t_R _18855_ (.A(_10466_),
    .B(_10114_),
    .Y(_10656_));
 NAND2x1_ASAP7_75t_R _18856_ (.A(net5567),
    .B(net5936),
    .Y(_10657_));
 OA21x2_ASAP7_75t_R _18857_ (.A1(_10314_),
    .A2(net5936),
    .B(net5917),
    .Y(_10658_));
 AOI21x1_ASAP7_75t_R _18858_ (.A1(_10657_),
    .A2(_10658_),
    .B(net5933),
    .Y(_10659_));
 OAI21x1_ASAP7_75t_R _18859_ (.A1(_10655_),
    .A2(_10656_),
    .B(_10659_),
    .Y(_10660_));
 NAND2x1_ASAP7_75t_R _18860_ (.A(_01060_),
    .B(net5935),
    .Y(_10661_));
 OAI21x1_ASAP7_75t_R _18861_ (.A1(net5935),
    .A2(_10217_),
    .B(_10661_),
    .Y(_10662_));
 OA21x2_ASAP7_75t_R _18862_ (.A1(net4962),
    .A2(net5936),
    .B(net5917),
    .Y(_10663_));
 AOI21x1_ASAP7_75t_R _18863_ (.A1(_10662_),
    .A2(_10663_),
    .B(net5558),
    .Y(_10664_));
 INVx1_ASAP7_75t_R _18864_ (.A(_01055_),
    .Y(_10665_));
 NOR2x1_ASAP7_75t_R _18865_ (.A(_10665_),
    .B(_10579_),
    .Y(_10666_));
 OAI21x1_ASAP7_75t_R _18866_ (.A1(_10367_),
    .A2(_10666_),
    .B(net6297),
    .Y(_10667_));
 AOI21x1_ASAP7_75t_R _18867_ (.A1(_10664_),
    .A2(_10667_),
    .B(net5932),
    .Y(_10668_));
 AOI21x1_ASAP7_75t_R _18868_ (.A1(_10660_),
    .A2(_10668_),
    .B(_10189_),
    .Y(_10669_));
 NAND2x1_ASAP7_75t_R _18869_ (.A(_10654_),
    .B(_10669_),
    .Y(_10670_));
 OAI21x1_ASAP7_75t_R _18870_ (.A1(_10629_),
    .A2(_10641_),
    .B(_10670_),
    .Y(_00031_));
 NOR2x1_ASAP7_75t_R _18875_ (.A(_00444_),
    .B(net6666),
    .Y(_10675_));
 INVx4_ASAP7_75t_R _18876_ (.A(_00574_),
    .Y(_10676_));
 XOR2x2_ASAP7_75t_R _18879_ (.A(_00582_),
    .B(net6652),
    .Y(_10679_));
 XOR2x2_ASAP7_75t_R _18880_ (.A(net6621),
    .B(net6597),
    .Y(_10680_));
 XOR2x2_ASAP7_75t_R _18881_ (.A(_10680_),
    .B(_10679_),
    .Y(_10681_));
 XOR2x2_ASAP7_75t_R _18882_ (.A(net6623),
    .B(net6618),
    .Y(_10682_));
 XOR2x2_ASAP7_75t_R _18883_ (.A(net6450),
    .B(net6565),
    .Y(_10683_));
 XOR2x2_ASAP7_75t_R _18884_ (.A(_10681_),
    .B(_10683_),
    .Y(_10684_));
 NOR2x1p5_ASAP7_75t_R _18885_ (.A(net6461),
    .B(_10684_),
    .Y(_10685_));
 OAI21x1_ASAP7_75t_R _18886_ (.A1(_10675_),
    .A2(net6366),
    .B(net6527),
    .Y(_10686_));
 AND2x2_ASAP7_75t_R _18889_ (.A(net6461),
    .B(_00444_),
    .Y(_10689_));
 XNOR2x2_ASAP7_75t_R _18891_ (.A(_10683_),
    .B(_10681_),
    .Y(_10691_));
 NOR2x1p5_ASAP7_75t_R _18892_ (.A(net6461),
    .B(_10691_),
    .Y(_10692_));
 INVx1_ASAP7_75t_R _18893_ (.A(net6527),
    .Y(_10693_));
 OAI21x1_ASAP7_75t_R _18894_ (.A1(_10689_),
    .A2(net6365),
    .B(_10693_),
    .Y(_10694_));
 NAND2x1p5_ASAP7_75t_R _18895_ (.A(_10686_),
    .B(_10694_),
    .Y(_10695_));
 INVx1_ASAP7_75t_R _18897_ (.A(net6567),
    .Y(_10696_));
 XOR2x2_ASAP7_75t_R _18898_ (.A(net6644),
    .B(net6617),
    .Y(_10697_));
 NAND2x1_ASAP7_75t_R _18899_ (.A(net6449),
    .B(_10697_),
    .Y(_10698_));
 XNOR2x2_ASAP7_75t_R _18900_ (.A(net6644),
    .B(net6617),
    .Y(_10699_));
 NAND2x1_ASAP7_75t_R _18901_ (.A(net6567),
    .B(_10699_),
    .Y(_10700_));
 XOR2x2_ASAP7_75t_R _18902_ (.A(net6598),
    .B(net6622),
    .Y(_10701_));
 INVx2_ASAP7_75t_R _18903_ (.A(_10701_),
    .Y(_10702_));
 AOI21x1_ASAP7_75t_R _18904_ (.A1(_10698_),
    .A2(_10700_),
    .B(_10702_),
    .Y(_10703_));
 NAND2x1_ASAP7_75t_R _18905_ (.A(net6567),
    .B(_10697_),
    .Y(_10704_));
 NAND2x1_ASAP7_75t_R _18906_ (.A(net6449),
    .B(_10699_),
    .Y(_10705_));
 AOI21x1_ASAP7_75t_R _18907_ (.A1(_10704_),
    .A2(_10705_),
    .B(net6448),
    .Y(_10706_));
 OAI21x1_ASAP7_75t_R _18908_ (.A1(_10703_),
    .A2(_10706_),
    .B(net6668),
    .Y(_10707_));
 INVx1_ASAP7_75t_R _18909_ (.A(net6528),
    .Y(_10708_));
 NOR2x1_ASAP7_75t_R _18912_ (.A(net6668),
    .B(_00445_),
    .Y(_10711_));
 INVx1_ASAP7_75t_R _18913_ (.A(_10711_),
    .Y(_10712_));
 NAND3x1_ASAP7_75t_R _18914_ (.A(net6364),
    .B(_10708_),
    .C(_10712_),
    .Y(_10713_));
 AO21x1_ASAP7_75t_R _18915_ (.A1(net6364),
    .A2(_10712_),
    .B(_10708_),
    .Y(_10714_));
 NAND2x1_ASAP7_75t_R _18916_ (.A(_10713_),
    .B(_10714_),
    .Y(_10715_));
 INVx1_ASAP7_75t_R _18918_ (.A(net6620),
    .Y(_10716_));
 XOR2x2_ASAP7_75t_R _18919_ (.A(net6649),
    .B(net6621),
    .Y(_10717_));
 NAND2x1_ASAP7_75t_R _18920_ (.A(_10716_),
    .B(net6447),
    .Y(_10718_));
 XNOR2x2_ASAP7_75t_R _18921_ (.A(net6621),
    .B(net6649),
    .Y(_10719_));
 NAND2x1_ASAP7_75t_R _18922_ (.A(net6620),
    .B(net6446),
    .Y(_10720_));
 XNOR2x2_ASAP7_75t_R _18923_ (.A(_00641_),
    .B(_00673_),
    .Y(_10721_));
 AOI21x1_ASAP7_75t_R _18924_ (.A1(_10718_),
    .A2(_10720_),
    .B(_10721_),
    .Y(_10722_));
 NAND2x1_ASAP7_75t_R _18925_ (.A(net6620),
    .B(net6447),
    .Y(_10723_));
 NAND2x1_ASAP7_75t_R _18926_ (.A(_10716_),
    .B(net6446),
    .Y(_10724_));
 XOR2x2_ASAP7_75t_R _18927_ (.A(_00641_),
    .B(_00673_),
    .Y(_10725_));
 AOI21x1_ASAP7_75t_R _18928_ (.A1(_10723_),
    .A2(_10724_),
    .B(_10725_),
    .Y(_10726_));
 OAI21x1_ASAP7_75t_R _18929_ (.A1(_10722_),
    .A2(_10726_),
    .B(net6668),
    .Y(_10727_));
 NOR2x1_ASAP7_75t_R _18930_ (.A(net6667),
    .B(_00446_),
    .Y(_10728_));
 INVx1_ASAP7_75t_R _18931_ (.A(_10728_),
    .Y(_10729_));
 NAND3x1_ASAP7_75t_R _18932_ (.A(_10727_),
    .B(net6526),
    .C(_10729_),
    .Y(_10730_));
 AO21x1_ASAP7_75t_R _18933_ (.A1(_10727_),
    .A2(_10729_),
    .B(net6526),
    .Y(_10731_));
 NAND2x1_ASAP7_75t_R _18934_ (.A(_10730_),
    .B(_10731_),
    .Y(_10732_));
 NAND3x1_ASAP7_75t_R _18937_ (.A(_10707_),
    .B(net6528),
    .C(_10712_),
    .Y(_10734_));
 AO21x1_ASAP7_75t_R _18938_ (.A1(_10707_),
    .A2(_10712_),
    .B(net6528),
    .Y(_10735_));
 NAND2x1p5_ASAP7_75t_R _18939_ (.A(_10734_),
    .B(_10735_),
    .Y(_10736_));
 INVx1_ASAP7_75t_R _18941_ (.A(net6526),
    .Y(_10737_));
 NAND3x1_ASAP7_75t_R _18942_ (.A(_10727_),
    .B(_10737_),
    .C(_10729_),
    .Y(_10738_));
 AO21x1_ASAP7_75t_R _18943_ (.A1(_10727_),
    .A2(_10729_),
    .B(_10737_),
    .Y(_10739_));
 NAND2x1_ASAP7_75t_R _18945_ (.A(_10738_),
    .B(_10739_),
    .Y(_10741_));
 XOR2x2_ASAP7_75t_R _18948_ (.A(_00580_),
    .B(_00612_),
    .Y(_10743_));
 XOR2x2_ASAP7_75t_R _18949_ (.A(_00613_),
    .B(_00645_),
    .Y(_10744_));
 XOR2x2_ASAP7_75t_R _18950_ (.A(_10744_),
    .B(_00677_),
    .Y(_10745_));
 XNOR2x2_ASAP7_75t_R _18951_ (.A(_10743_),
    .B(_10745_),
    .Y(_10746_));
 NOR2x1_ASAP7_75t_R _18955_ (.A(net6665),
    .B(_00550_),
    .Y(_10750_));
 AO21x1_ASAP7_75t_R _18956_ (.A1(_10746_),
    .A2(net6665),
    .B(_10750_),
    .Y(_10751_));
 XOR2x2_ASAP7_75t_R _18957_ (.A(_10751_),
    .B(net6521),
    .Y(_10752_));
 INVx1_ASAP7_75t_R _18958_ (.A(_10752_),
    .Y(_10753_));
 NOR2x1_ASAP7_75t_R _18961_ (.A(net5309),
    .B(net5903),
    .Y(_10756_));
 XOR2x2_ASAP7_75t_R _18962_ (.A(_00577_),
    .B(net6643),
    .Y(_10757_));
 INVx1_ASAP7_75t_R _18963_ (.A(net6619),
    .Y(_10758_));
 XOR2x2_ASAP7_75t_R _18964_ (.A(_10757_),
    .B(_10758_),
    .Y(_10759_));
 XNOR2x2_ASAP7_75t_R _18965_ (.A(_00642_),
    .B(_00674_),
    .Y(_10760_));
 XOR2x2_ASAP7_75t_R _18966_ (.A(_00609_),
    .B(net6617),
    .Y(_10761_));
 XOR2x2_ASAP7_75t_R _18967_ (.A(_10760_),
    .B(_10761_),
    .Y(_10762_));
 NOR2x1_ASAP7_75t_R _18968_ (.A(_10759_),
    .B(_10762_),
    .Y(_10763_));
 AO21x1_ASAP7_75t_R _18970_ (.A1(_10762_),
    .A2(_10759_),
    .B(net6461),
    .Y(_10765_));
 NAND2x1_ASAP7_75t_R _18972_ (.A(_00553_),
    .B(net6461),
    .Y(_10767_));
 OAI21x1_ASAP7_75t_R _18973_ (.A1(_10763_),
    .A2(_10765_),
    .B(_10767_),
    .Y(_10768_));
 INVx1_ASAP7_75t_R _18974_ (.A(net6525),
    .Y(_10769_));
 XOR2x2_ASAP7_75t_R _18975_ (.A(_10768_),
    .B(_10769_),
    .Y(_10770_));
 XOR2x2_ASAP7_75t_R _18978_ (.A(net6645),
    .B(net6643),
    .Y(_10773_));
 XNOR2x2_ASAP7_75t_R _18979_ (.A(_00611_),
    .B(_10773_),
    .Y(_10774_));
 XOR2x2_ASAP7_75t_R _18980_ (.A(net6619),
    .B(net6617),
    .Y(_10775_));
 XOR2x2_ASAP7_75t_R _18981_ (.A(_00643_),
    .B(_00675_),
    .Y(_10776_));
 XNOR2x2_ASAP7_75t_R _18982_ (.A(_10775_),
    .B(_10776_),
    .Y(_10777_));
 NOR2x1_ASAP7_75t_R _18983_ (.A(_10774_),
    .B(_10777_),
    .Y(_10778_));
 AO21x1_ASAP7_75t_R _18985_ (.A1(_10777_),
    .A2(_10774_),
    .B(net6461),
    .Y(_10780_));
 NAND2x1_ASAP7_75t_R _18987_ (.A(_00552_),
    .B(net6461),
    .Y(_10782_));
 OAI21x1_ASAP7_75t_R _18988_ (.A1(_10778_),
    .A2(_10780_),
    .B(_10782_),
    .Y(_10783_));
 XOR2x2_ASAP7_75t_R _18989_ (.A(_10783_),
    .B(net6524),
    .Y(_10784_));
 AO21x1_ASAP7_75t_R _18992_ (.A1(_10756_),
    .A2(net6274),
    .B(net6272),
    .Y(_10787_));
 INVx1_ASAP7_75t_R _18995_ (.A(_01070_),
    .Y(_10790_));
 AOI21x1_ASAP7_75t_R _18996_ (.A1(net6284),
    .A2(net6283),
    .B(_10790_),
    .Y(_10791_));
 NOR2x1_ASAP7_75t_R _18998_ (.A(_10791_),
    .B(_10770_),
    .Y(_10793_));
 INVx1_ASAP7_75t_R _18999_ (.A(_10793_),
    .Y(_10794_));
 AOI211x1_ASAP7_75t_R _19001_ (.A1(net6285),
    .A2(net6286),
    .B(net5904),
    .C(net5906),
    .Y(_10796_));
 NOR2x1_ASAP7_75t_R _19002_ (.A(_10794_),
    .B(_10796_),
    .Y(_10797_));
 INVx1_ASAP7_75t_R _19003_ (.A(_00551_),
    .Y(_10798_));
 NAND2x1_ASAP7_75t_R _19004_ (.A(net6461),
    .B(_10798_),
    .Y(_10799_));
 XOR2x2_ASAP7_75t_R _19005_ (.A(_00579_),
    .B(_00611_),
    .Y(_10800_));
 INVx1_ASAP7_75t_R _19006_ (.A(_10800_),
    .Y(_10801_));
 XOR2x2_ASAP7_75t_R _19007_ (.A(_00612_),
    .B(_00644_),
    .Y(_10802_));
 INVx1_ASAP7_75t_R _19008_ (.A(_00676_),
    .Y(_10803_));
 XOR2x2_ASAP7_75t_R _19009_ (.A(_10802_),
    .B(_10803_),
    .Y(_10804_));
 NAND2x1_ASAP7_75t_R _19010_ (.A(_10801_),
    .B(_10804_),
    .Y(_10805_));
 XOR2x2_ASAP7_75t_R _19011_ (.A(_10802_),
    .B(net6561),
    .Y(_10806_));
 NAND2x1_ASAP7_75t_R _19012_ (.A(_10800_),
    .B(_10806_),
    .Y(_10807_));
 AOI21x1_ASAP7_75t_R _19013_ (.A1(_10805_),
    .A2(_10807_),
    .B(net6461),
    .Y(_10808_));
 INVx1_ASAP7_75t_R _19014_ (.A(_10808_),
    .Y(_10809_));
 INVx1_ASAP7_75t_R _19015_ (.A(net6523),
    .Y(_10810_));
 AOI21x1_ASAP7_75t_R _19016_ (.A1(_10799_),
    .A2(_10809_),
    .B(_10810_),
    .Y(_10811_));
 AOI211x1_ASAP7_75t_R _19017_ (.A1(net6461),
    .A2(_10798_),
    .B(_10808_),
    .C(net6523),
    .Y(_10812_));
 NOR2x1_ASAP7_75t_R _19018_ (.A(_10811_),
    .B(_10812_),
    .Y(_10813_));
 INVx1_ASAP7_75t_R _19019_ (.A(_10813_),
    .Y(_10814_));
 OAI21x1_ASAP7_75t_R _19022_ (.A1(_10787_),
    .A2(_10797_),
    .B(net5219),
    .Y(_10817_));
 XNOR2x2_ASAP7_75t_R _19023_ (.A(net6524),
    .B(_10783_),
    .Y(_10818_));
 AOI21x1_ASAP7_75t_R _19026_ (.A1(net6284),
    .A2(net6283),
    .B(net5305),
    .Y(_10821_));
 XOR2x2_ASAP7_75t_R _19027_ (.A(_10768_),
    .B(net6525),
    .Y(_10822_));
 NOR2x1_ASAP7_75t_R _19029_ (.A(_10821_),
    .B(net6264),
    .Y(_10824_));
 INVx1_ASAP7_75t_R _19030_ (.A(_10824_),
    .Y(_10825_));
 AO21x1_ASAP7_75t_R _19031_ (.A1(net6279),
    .A2(net6280),
    .B(net5309),
    .Y(_10826_));
 NOR2x1_ASAP7_75t_R _19032_ (.A(net6273),
    .B(_10826_),
    .Y(_10827_));
 INVx1_ASAP7_75t_R _19033_ (.A(_10827_),
    .Y(_10828_));
 OAI21x1_ASAP7_75t_R _19034_ (.A1(_10825_),
    .A2(_10796_),
    .B(_10828_),
    .Y(_10829_));
 NOR2x1_ASAP7_75t_R _19035_ (.A(net6268),
    .B(_10829_),
    .Y(_10830_));
 AOI21x1_ASAP7_75t_R _19036_ (.A1(net6284),
    .A2(net6283),
    .B(net5308),
    .Y(_10831_));
 AOI21x1_ASAP7_75t_R _19037_ (.A1(net5907),
    .A2(net5899),
    .B(net5217),
    .Y(_10832_));
 OAI21x1_ASAP7_75t_R _19038_ (.A1(_10675_),
    .A2(_10685_),
    .B(_10693_),
    .Y(_10833_));
 OAI21x1_ASAP7_75t_R _19039_ (.A1(_10689_),
    .A2(_10692_),
    .B(net6527),
    .Y(_10834_));
 NAND2x1p5_ASAP7_75t_R _19040_ (.A(_10834_),
    .B(_10833_),
    .Y(_10835_));
 NAND2x1_ASAP7_75t_R _19041_ (.A(net5899),
    .B(net5893),
    .Y(_10836_));
 AOI21x1_ASAP7_75t_R _19044_ (.A1(_10832_),
    .A2(net5532),
    .B(net6266),
    .Y(_10839_));
 INVx1_ASAP7_75t_R _19045_ (.A(_01063_),
    .Y(_10840_));
 NOR2x1_ASAP7_75t_R _19046_ (.A(_10840_),
    .B(net5905),
    .Y(_10841_));
 NOR2x1_ASAP7_75t_R _19047_ (.A(net5901),
    .B(net5899),
    .Y(_10842_));
 NOR2x1_ASAP7_75t_R _19048_ (.A(_10841_),
    .B(_10842_),
    .Y(_10843_));
 AOI21x1_ASAP7_75t_R _19049_ (.A1(net6284),
    .A2(net6283),
    .B(net5309),
    .Y(_10844_));
 AOI21x1_ASAP7_75t_R _19052_ (.A1(_10844_),
    .A2(net6274),
    .B(_10784_),
    .Y(_10847_));
 OAI21x1_ASAP7_75t_R _19053_ (.A1(net6274),
    .A2(_10843_),
    .B(_10847_),
    .Y(_10848_));
 AOI21x1_ASAP7_75t_R _19054_ (.A1(net6284),
    .A2(net6283),
    .B(net5259),
    .Y(_10849_));
 AOI21x1_ASAP7_75t_R _19055_ (.A1(net5016),
    .A2(net6274),
    .B(net6268),
    .Y(_10850_));
 OR2x2_ASAP7_75t_R _19057_ (.A(_01077_),
    .B(net6274),
    .Y(_10852_));
 AOI21x1_ASAP7_75t_R _19059_ (.A1(_10850_),
    .A2(_10852_),
    .B(net5219),
    .Y(_10854_));
 OAI21x1_ASAP7_75t_R _19060_ (.A1(_10839_),
    .A2(_10848_),
    .B(_10854_),
    .Y(_10855_));
 OAI21x1_ASAP7_75t_R _19061_ (.A1(_10817_),
    .A2(_10830_),
    .B(_10855_),
    .Y(_10856_));
 XNOR2x2_ASAP7_75t_R _19062_ (.A(_00581_),
    .B(_00613_),
    .Y(_10857_));
 INVx1_ASAP7_75t_R _19063_ (.A(net6560),
    .Y(_10858_));
 XOR2x2_ASAP7_75t_R _19064_ (.A(_10857_),
    .B(net6445),
    .Y(_10859_));
 XNOR2x2_ASAP7_75t_R _19065_ (.A(net6617),
    .B(net6593),
    .Y(_10860_));
 XOR2x2_ASAP7_75t_R _19066_ (.A(_10859_),
    .B(_10860_),
    .Y(_10861_));
 NOR2x1_ASAP7_75t_R _19070_ (.A(net6665),
    .B(_00549_),
    .Y(_10865_));
 AO21x1_ASAP7_75t_R _19071_ (.A1(_10861_),
    .A2(net6668),
    .B(_10865_),
    .Y(_10866_));
 XOR2x2_ASAP7_75t_R _19072_ (.A(_10866_),
    .B(net6520),
    .Y(_10867_));
 INVx1_ASAP7_75t_R _19073_ (.A(_10867_),
    .Y(_10868_));
 OAI21x1_ASAP7_75t_R _19074_ (.A1(net5895),
    .A2(_10856_),
    .B(_10868_),
    .Y(_10869_));
 NAND2x1_ASAP7_75t_R _19075_ (.A(net5906),
    .B(net5898),
    .Y(_10870_));
 INVx1_ASAP7_75t_R _19076_ (.A(_01069_),
    .Y(_10871_));
 AO21x1_ASAP7_75t_R _19077_ (.A1(net6283),
    .A2(net6284),
    .B(_10871_),
    .Y(_10872_));
 AO21x1_ASAP7_75t_R _19078_ (.A1(net5530),
    .A2(_10872_),
    .B(net6276),
    .Y(_10873_));
 NOR2x1_ASAP7_75t_R _19079_ (.A(_10784_),
    .B(_10813_),
    .Y(_10874_));
 INVx1_ASAP7_75t_R _19080_ (.A(_10874_),
    .Y(_10875_));
 OAI21x1_ASAP7_75t_R _19082_ (.A1(net5903),
    .A2(net5893),
    .B(net6276),
    .Y(_10876_));
 NOR2x1_ASAP7_75t_R _19083_ (.A(net5016),
    .B(_10876_),
    .Y(_10877_));
 NOR2x1_ASAP7_75t_R _19084_ (.A(_10875_),
    .B(_10877_),
    .Y(_10878_));
 AOI21x1_ASAP7_75t_R _19085_ (.A1(net6284),
    .A2(net6283),
    .B(_10840_),
    .Y(_10879_));
 OA21x2_ASAP7_75t_R _19087_ (.A1(_10756_),
    .A2(net4960),
    .B(net6276),
    .Y(_10881_));
 INVx1_ASAP7_75t_R _19088_ (.A(_01067_),
    .Y(_10882_));
 OAI21x1_ASAP7_75t_R _19090_ (.A1(net5213),
    .A2(net5902),
    .B(net6266),
    .Y(_10884_));
 OAI21x1_ASAP7_75t_R _19091_ (.A1(_10812_),
    .A2(_10811_),
    .B(_10784_),
    .Y(_10885_));
 INVx1_ASAP7_75t_R _19092_ (.A(_10885_),
    .Y(_10886_));
 NAND2x1_ASAP7_75t_R _19093_ (.A(_10884_),
    .B(_10886_),
    .Y(_10887_));
 NOR2x1_ASAP7_75t_R _19094_ (.A(_10881_),
    .B(_10887_),
    .Y(_10888_));
 AOI21x1_ASAP7_75t_R _19095_ (.A1(_10873_),
    .A2(_10878_),
    .B(_10888_),
    .Y(_10889_));
 NAND2x1_ASAP7_75t_R _19097_ (.A(net5905),
    .B(net5900),
    .Y(_10891_));
 NAND2x1_ASAP7_75t_R _19098_ (.A(net6265),
    .B(_10891_),
    .Y(_10892_));
 AOI211x1_ASAP7_75t_R _19099_ (.A1(net6285),
    .A2(net6286),
    .B(net5904),
    .C(net5900),
    .Y(_10893_));
 AOI21x1_ASAP7_75t_R _19100_ (.A1(net5216),
    .A2(net6277),
    .B(net6271),
    .Y(_10894_));
 OAI21x1_ASAP7_75t_R _19101_ (.A1(_10892_),
    .A2(_10893_),
    .B(_10894_),
    .Y(_10895_));
 INVx1_ASAP7_75t_R _19102_ (.A(_10895_),
    .Y(_10896_));
 INVx1_ASAP7_75t_R _19103_ (.A(_10831_),
    .Y(_10897_));
 AO21x1_ASAP7_75t_R _19104_ (.A1(_10739_),
    .A2(net6280),
    .B(_01070_),
    .Y(_10898_));
 NAND2x1_ASAP7_75t_R _19106_ (.A(_10897_),
    .B(_10898_),
    .Y(_10900_));
 INVx1_ASAP7_75t_R _19107_ (.A(_01064_),
    .Y(_10901_));
 AO21x1_ASAP7_75t_R _19108_ (.A1(_10739_),
    .A2(net6280),
    .B(_10901_),
    .Y(_10902_));
 NAND2x2_ASAP7_75t_R _19110_ (.A(_10902_),
    .B(net6265),
    .Y(_10904_));
 INVx2_ASAP7_75t_R _19111_ (.A(_10904_),
    .Y(_10905_));
 AOI211x1_ASAP7_75t_R _19112_ (.A1(net4708),
    .A2(net6276),
    .B(_10905_),
    .C(net6268),
    .Y(_10906_));
 OAI21x1_ASAP7_75t_R _19114_ (.A1(_10896_),
    .A2(_10906_),
    .B(net5533),
    .Y(_10908_));
 AOI21x1_ASAP7_75t_R _19116_ (.A1(_10889_),
    .A2(_10908_),
    .B(net6278),
    .Y(_10910_));
 AO21x1_ASAP7_75t_R _19117_ (.A1(_10841_),
    .A2(net6274),
    .B(net6272),
    .Y(_10911_));
 AOI21x1_ASAP7_75t_R _19118_ (.A1(net6280),
    .A2(net6279),
    .B(net5259),
    .Y(_10912_));
 INVx2_ASAP7_75t_R _19119_ (.A(_10912_),
    .Y(_10913_));
 INVx1_ASAP7_75t_R _19120_ (.A(_10879_),
    .Y(_10914_));
 AO21x1_ASAP7_75t_R _19121_ (.A1(_10913_),
    .A2(_10914_),
    .B(net6276),
    .Y(_10915_));
 OAI21x1_ASAP7_75t_R _19122_ (.A1(net6266),
    .A2(_10872_),
    .B(_10915_),
    .Y(_10916_));
 OAI21x1_ASAP7_75t_R _19123_ (.A1(_10911_),
    .A2(_10916_),
    .B(net6278),
    .Y(_10917_));
 NOR2x1_ASAP7_75t_R _19124_ (.A(net5014),
    .B(net5905),
    .Y(_10918_));
 AOI21x1_ASAP7_75t_R _19125_ (.A1(net6284),
    .A2(net6283),
    .B(net5015),
    .Y(_10919_));
 NOR2x2_ASAP7_75t_R _19126_ (.A(net6274),
    .B(_10919_),
    .Y(_10920_));
 AO21x1_ASAP7_75t_R _19127_ (.A1(net6274),
    .A2(_10918_),
    .B(_10920_),
    .Y(_10921_));
 NAND2x1_ASAP7_75t_R _19129_ (.A(net5905),
    .B(net5892),
    .Y(_10923_));
 NOR2x1_ASAP7_75t_R _19130_ (.A(net6265),
    .B(_10923_),
    .Y(_10924_));
 OA21x2_ASAP7_75t_R _19132_ (.A1(_10921_),
    .A2(_10924_),
    .B(net6271),
    .Y(_10926_));
 NOR2x1_ASAP7_75t_R _19133_ (.A(_10917_),
    .B(_10926_),
    .Y(_10927_));
 OAI21x1_ASAP7_75t_R _19135_ (.A1(_10892_),
    .A2(_10893_),
    .B(net6267),
    .Y(_10929_));
 NOR2x1_ASAP7_75t_R _19137_ (.A(net5897),
    .B(net5910),
    .Y(_10931_));
 OA21x2_ASAP7_75t_R _19138_ (.A1(_10931_),
    .A2(_10756_),
    .B(net6277),
    .Y(_10932_));
 NOR2x1_ASAP7_75t_R _19139_ (.A(_10929_),
    .B(_10932_),
    .Y(_10933_));
 INVx1_ASAP7_75t_R _19140_ (.A(_01072_),
    .Y(_10934_));
 NOR2x1_ASAP7_75t_R _19141_ (.A(_10934_),
    .B(net5902),
    .Y(_10935_));
 OAI21x1_ASAP7_75t_R _19143_ (.A1(net4958),
    .A2(_10892_),
    .B(net6271),
    .Y(_10937_));
 OAI21x1_ASAP7_75t_R _19144_ (.A1(net5904),
    .A2(net5908),
    .B(net6277),
    .Y(_10938_));
 NOR3x1_ASAP7_75t_R _19145_ (.A(net5892),
    .B(net5906),
    .C(net5897),
    .Y(_10939_));
 NOR2x1_ASAP7_75t_R _19146_ (.A(_10938_),
    .B(_10939_),
    .Y(_10940_));
 OAI21x1_ASAP7_75t_R _19147_ (.A1(_10937_),
    .A2(_10940_),
    .B(net5895),
    .Y(_10941_));
 OAI21x1_ASAP7_75t_R _19148_ (.A1(_10933_),
    .A2(_10941_),
    .B(net5533),
    .Y(_10942_));
 NOR2x1_ASAP7_75t_R _19149_ (.A(_10942_),
    .B(_10927_),
    .Y(_10943_));
 NOR2x1_ASAP7_75t_R _19150_ (.A(net5906),
    .B(net5910),
    .Y(_10944_));
 NAND2x1_ASAP7_75t_R _19151_ (.A(net6277),
    .B(_10870_),
    .Y(_10945_));
 NOR2x1_ASAP7_75t_R _19152_ (.A(_10944_),
    .B(_10945_),
    .Y(_10946_));
 OAI21x1_ASAP7_75t_R _19153_ (.A1(net5907),
    .A2(net5893),
    .B(net6266),
    .Y(_10947_));
 OAI21x1_ASAP7_75t_R _19154_ (.A1(_10842_),
    .A2(_10947_),
    .B(net6272),
    .Y(_10948_));
 NOR2x1_ASAP7_75t_R _19155_ (.A(_10946_),
    .B(_10948_),
    .Y(_10949_));
 INVx1_ASAP7_75t_R _19156_ (.A(net6286),
    .Y(_10950_));
 INVx1_ASAP7_75t_R _19157_ (.A(net6285),
    .Y(_10951_));
 OAI21x1_ASAP7_75t_R _19158_ (.A1(_10950_),
    .A2(_10951_),
    .B(net5906),
    .Y(_10952_));
 INVx1_ASAP7_75t_R _19159_ (.A(_10952_),
    .Y(_10953_));
 NAND2x1_ASAP7_75t_R _19160_ (.A(net6275),
    .B(net4781),
    .Y(_10954_));
 AOI21x1_ASAP7_75t_R _19161_ (.A1(net5902),
    .A2(_10953_),
    .B(_10954_),
    .Y(_10955_));
 NOR2x1_ASAP7_75t_R _19162_ (.A(net5215),
    .B(net5903),
    .Y(_10956_));
 OAI21x1_ASAP7_75t_R _19163_ (.A1(net4960),
    .A2(_10956_),
    .B(net6265),
    .Y(_10957_));
 NAND2x1_ASAP7_75t_R _19164_ (.A(net6267),
    .B(_10957_),
    .Y(_10958_));
 OAI21x1_ASAP7_75t_R _19165_ (.A1(_10955_),
    .A2(_10958_),
    .B(net6278),
    .Y(_10959_));
 NOR2x1_ASAP7_75t_R _19166_ (.A(_10949_),
    .B(_10959_),
    .Y(_10960_));
 NOR2x1_ASAP7_75t_R _19167_ (.A(_10934_),
    .B(net5898),
    .Y(_10961_));
 OAI21x1_ASAP7_75t_R _19168_ (.A1(net4957),
    .A2(net4595),
    .B(net6271),
    .Y(_10962_));
 NAND2x1_ASAP7_75t_R _19169_ (.A(net6277),
    .B(net5892),
    .Y(_10963_));
 NAND2x1_ASAP7_75t_R _19170_ (.A(net6277),
    .B(_10891_),
    .Y(_10964_));
 NOR2x1_ASAP7_75t_R _19171_ (.A(net5904),
    .B(net5906),
    .Y(_10965_));
 AOI21x1_ASAP7_75t_R _19172_ (.A1(_10963_),
    .A2(_10964_),
    .B(_10965_),
    .Y(_10966_));
 NOR2x1_ASAP7_75t_R _19173_ (.A(_10962_),
    .B(_10966_),
    .Y(_10967_));
 AO21x1_ASAP7_75t_R _19174_ (.A1(_10891_),
    .A2(net6277),
    .B(net6271),
    .Y(_10968_));
 NOR2x1_ASAP7_75t_R _19175_ (.A(net5906),
    .B(net5892),
    .Y(_10969_));
 AOI21x1_ASAP7_75t_R _19176_ (.A1(net5902),
    .A2(_10969_),
    .B(_10884_),
    .Y(_10970_));
 OAI21x1_ASAP7_75t_R _19177_ (.A1(_10968_),
    .A2(_10970_),
    .B(net5895),
    .Y(_10971_));
 OAI21x1_ASAP7_75t_R _19178_ (.A1(_10967_),
    .A2(_10971_),
    .B(net5220),
    .Y(_10972_));
 OAI21x1_ASAP7_75t_R _19179_ (.A1(_10960_),
    .A2(_10972_),
    .B(net6263),
    .Y(_10973_));
 OAI22x1_ASAP7_75t_R _19180_ (.A1(_10869_),
    .A2(_10910_),
    .B1(_10943_),
    .B2(_10973_),
    .Y(_00032_));
 OAI21x1_ASAP7_75t_R _19182_ (.A1(net5900),
    .A2(net5892),
    .B(net5897),
    .Y(_10975_));
 NOR2x1_ASAP7_75t_R _19183_ (.A(net6265),
    .B(_10975_),
    .Y(_10976_));
 NOR2x1_ASAP7_75t_R _19184_ (.A(net5903),
    .B(net5910),
    .Y(_10977_));
 AO21x1_ASAP7_75t_R _19185_ (.A1(net5304),
    .A2(net5903),
    .B(net6277),
    .Y(_10978_));
 OAI21x1_ASAP7_75t_R _19186_ (.A1(_10977_),
    .A2(_10978_),
    .B(net6271),
    .Y(_10979_));
 NOR2x1_ASAP7_75t_R _19187_ (.A(_10976_),
    .B(_10979_),
    .Y(_10980_));
 OAI21x1_ASAP7_75t_R _19188_ (.A1(net5896),
    .A2(_10952_),
    .B(net6264),
    .Y(_10981_));
 AO21x1_ASAP7_75t_R _19189_ (.A1(net6279),
    .A2(net6280),
    .B(net5307),
    .Y(_10982_));
 OA21x2_ASAP7_75t_R _19190_ (.A1(_10982_),
    .A2(net6265),
    .B(_10818_),
    .Y(_10983_));
 OA21x2_ASAP7_75t_R _19191_ (.A1(_10981_),
    .A2(net5013),
    .B(_10983_),
    .Y(_10984_));
 OAI21x1_ASAP7_75t_R _19192_ (.A1(_10980_),
    .A2(_10984_),
    .B(net5221),
    .Y(_10985_));
 AO21x1_ASAP7_75t_R _19193_ (.A1(net6279),
    .A2(net6280),
    .B(_10840_),
    .Y(_10986_));
 NAND2x1_ASAP7_75t_R _19194_ (.A(net5902),
    .B(net5906),
    .Y(_10987_));
 NAND2x1_ASAP7_75t_R _19195_ (.A(_10986_),
    .B(_10987_),
    .Y(_10988_));
 OA21x2_ASAP7_75t_R _19196_ (.A1(net4595),
    .A2(net5216),
    .B(net6271),
    .Y(_10989_));
 OAI21x1_ASAP7_75t_R _19197_ (.A1(net6265),
    .A2(_10988_),
    .B(_10989_),
    .Y(_10990_));
 NOR2x1_ASAP7_75t_R _19198_ (.A(net5900),
    .B(net5910),
    .Y(_10991_));
 NAND2x1_ASAP7_75t_R _19199_ (.A(net5901),
    .B(net5899),
    .Y(_10992_));
 NOR2x1_ASAP7_75t_R _19200_ (.A(net5016),
    .B(net6265),
    .Y(_10993_));
 NAND2x1_ASAP7_75t_R _19201_ (.A(_10992_),
    .B(_10993_),
    .Y(_10994_));
 OAI21x1_ASAP7_75t_R _19202_ (.A1(_10892_),
    .A2(_10991_),
    .B(_10994_),
    .Y(_10995_));
 AOI21x1_ASAP7_75t_R _19203_ (.A1(net6267),
    .A2(_10995_),
    .B(net5220),
    .Y(_10996_));
 AOI21x1_ASAP7_75t_R _19204_ (.A1(_10990_),
    .A2(_10996_),
    .B(net6278),
    .Y(_10997_));
 NAND2x1_ASAP7_75t_R _19205_ (.A(_10985_),
    .B(_10997_),
    .Y(_10998_));
 NAND2x1_ASAP7_75t_R _19206_ (.A(net5903),
    .B(net5910),
    .Y(_10999_));
 AOI21x1_ASAP7_75t_R _19207_ (.A1(net6265),
    .A2(net5525),
    .B(_10977_),
    .Y(_11000_));
 OA21x2_ASAP7_75t_R _19208_ (.A1(net4959),
    .A2(net6265),
    .B(net6272),
    .Y(_11001_));
 AO21x1_ASAP7_75t_R _19209_ (.A1(_11000_),
    .A2(_11001_),
    .B(net5220),
    .Y(_11002_));
 INVx1_ASAP7_75t_R _19210_ (.A(_10935_),
    .Y(_11003_));
 AOI211x1_ASAP7_75t_R _19211_ (.A1(net4593),
    .A2(net4707),
    .B(_10839_),
    .C(net6272),
    .Y(_11004_));
 NAND2x1_ASAP7_75t_R _19212_ (.A(net5903),
    .B(net6265),
    .Y(_11005_));
 OAI22x1_ASAP7_75t_R _19213_ (.A1(_10876_),
    .A2(net5527),
    .B1(_11005_),
    .B2(_10969_),
    .Y(_11006_));
 OAI21x1_ASAP7_75t_R _19214_ (.A1(net5012),
    .A2(_10842_),
    .B(net6266),
    .Y(_11007_));
 AOI21x1_ASAP7_75t_R _19215_ (.A1(net6280),
    .A2(net6279),
    .B(_10882_),
    .Y(_11008_));
 NOR2x1p5_ASAP7_75t_R _19216_ (.A(_11008_),
    .B(net6266),
    .Y(_11009_));
 NAND2x1_ASAP7_75t_R _19217_ (.A(_10987_),
    .B(net4706),
    .Y(_11010_));
 AOI21x1_ASAP7_75t_R _19218_ (.A1(_11007_),
    .A2(_11010_),
    .B(net5529),
    .Y(_11011_));
 AOI21x1_ASAP7_75t_R _19219_ (.A1(net5214),
    .A2(_11006_),
    .B(_11011_),
    .Y(_11012_));
 OAI21x1_ASAP7_75t_R _19220_ (.A1(_11002_),
    .A2(_11004_),
    .B(_11012_),
    .Y(_11013_));
 AOI21x1_ASAP7_75t_R _19221_ (.A1(net6278),
    .A2(_11013_),
    .B(net6263),
    .Y(_11014_));
 INVx1_ASAP7_75t_R _19222_ (.A(_10945_),
    .Y(_11015_));
 AOI21x1_ASAP7_75t_R _19223_ (.A1(net5525),
    .A2(_11015_),
    .B(net5220),
    .Y(_11016_));
 NOR2x1p5_ASAP7_75t_R _19224_ (.A(_11008_),
    .B(net6277),
    .Y(_11017_));
 AOI21x1_ASAP7_75t_R _19225_ (.A1(_11017_),
    .A2(_10923_),
    .B(net6267),
    .Y(_11018_));
 AND2x2_ASAP7_75t_R _19226_ (.A(_11016_),
    .B(_11018_),
    .Y(_11019_));
 AO21x1_ASAP7_75t_R _19227_ (.A1(net6283),
    .A2(net6284),
    .B(_01063_),
    .Y(_11020_));
 NAND2x1_ASAP7_75t_R _19228_ (.A(net6277),
    .B(_11020_),
    .Y(_11021_));
 NOR2x1_ASAP7_75t_R _19229_ (.A(_10965_),
    .B(_11021_),
    .Y(_11022_));
 NOR2x1_ASAP7_75t_R _19230_ (.A(net5904),
    .B(net6277),
    .Y(_11023_));
 NAND2x1_ASAP7_75t_R _19231_ (.A(_10952_),
    .B(_11023_),
    .Y(_11024_));
 NOR2x1_ASAP7_75t_R _19232_ (.A(net5899),
    .B(net6274),
    .Y(_11025_));
 NAND2x1_ASAP7_75t_R _19233_ (.A(net5900),
    .B(net5910),
    .Y(_11026_));
 AOI21x1_ASAP7_75t_R _19234_ (.A1(_11025_),
    .A2(_11026_),
    .B(net5529),
    .Y(_11027_));
 NAND2x1_ASAP7_75t_R _19235_ (.A(_11024_),
    .B(_11027_),
    .Y(_11028_));
 OAI21x1_ASAP7_75t_R _19236_ (.A1(net5905),
    .A2(_10952_),
    .B(_10824_),
    .Y(_11029_));
 INVx1_ASAP7_75t_R _19238_ (.A(_01079_),
    .Y(_11031_));
 NOR2x1_ASAP7_75t_R _19239_ (.A(_11031_),
    .B(net6273),
    .Y(_11032_));
 AOI21x1_ASAP7_75t_R _19240_ (.A1(net5533),
    .A2(_11032_),
    .B(net6271),
    .Y(_11033_));
 AOI21x1_ASAP7_75t_R _19241_ (.A1(_11029_),
    .A2(_11033_),
    .B(net5895),
    .Y(_11034_));
 OAI21x1_ASAP7_75t_R _19242_ (.A1(_11022_),
    .A2(_11028_),
    .B(_11034_),
    .Y(_11035_));
 OAI21x1_ASAP7_75t_R _19243_ (.A1(_11019_),
    .A2(_11035_),
    .B(net6263),
    .Y(_11036_));
 OAI21x1_ASAP7_75t_R _19244_ (.A1(_10756_),
    .A2(_10842_),
    .B(net6277),
    .Y(_11037_));
 INVx2_ASAP7_75t_R _19245_ (.A(net5016),
    .Y(_11038_));
 AO21x1_ASAP7_75t_R _19246_ (.A1(_10986_),
    .A2(_11038_),
    .B(net6277),
    .Y(_11039_));
 AOI21x1_ASAP7_75t_R _19247_ (.A1(_11037_),
    .A2(_11039_),
    .B(net6267),
    .Y(_11040_));
 OAI21x1_ASAP7_75t_R _19248_ (.A1(net4960),
    .A2(_10965_),
    .B(net6277),
    .Y(_11041_));
 NAND2x1_ASAP7_75t_R _19249_ (.A(_11017_),
    .B(_10923_),
    .Y(_11042_));
 AOI21x1_ASAP7_75t_R _19250_ (.A1(_11041_),
    .A2(_11042_),
    .B(net6271),
    .Y(_11043_));
 OAI21x1_ASAP7_75t_R _19251_ (.A1(_11040_),
    .A2(_11043_),
    .B(net5221),
    .Y(_11044_));
 INVx1_ASAP7_75t_R _19252_ (.A(net5309),
    .Y(_11045_));
 AO21x1_ASAP7_75t_R _19253_ (.A1(net6283),
    .A2(net6284),
    .B(_11045_),
    .Y(_11046_));
 AOI21x1_ASAP7_75t_R _19254_ (.A1(net5304),
    .A2(net5897),
    .B(net6265),
    .Y(_11047_));
 AOI21x1_ASAP7_75t_R _19255_ (.A1(net4955),
    .A2(_11047_),
    .B(net6267),
    .Y(_11048_));
 OAI21x1_ASAP7_75t_R _19256_ (.A1(net5013),
    .A2(_10981_),
    .B(_11048_),
    .Y(_11049_));
 NAND2x1_ASAP7_75t_R _19257_ (.A(net5896),
    .B(net5910),
    .Y(_11050_));
 AOI21x1_ASAP7_75t_R _19258_ (.A1(net5901),
    .A2(net5902),
    .B(net6266),
    .Y(_11051_));
 OAI21x1_ASAP7_75t_R _19259_ (.A1(net5900),
    .A2(_11050_),
    .B(_11051_),
    .Y(_11052_));
 NOR2x1_ASAP7_75t_R _19260_ (.A(net6271),
    .B(_10905_),
    .Y(_11053_));
 AOI21x1_ASAP7_75t_R _19261_ (.A1(_11052_),
    .A2(_11053_),
    .B(net5221),
    .Y(_11054_));
 NAND2x1_ASAP7_75t_R _19262_ (.A(_11049_),
    .B(_11054_),
    .Y(_11055_));
 AOI21x1_ASAP7_75t_R _19263_ (.A1(_11044_),
    .A2(_11055_),
    .B(net6278),
    .Y(_11056_));
 NOR2x1_ASAP7_75t_R _19264_ (.A(_11036_),
    .B(_11056_),
    .Y(_11057_));
 AOI21x1_ASAP7_75t_R _19265_ (.A1(_10998_),
    .A2(_11014_),
    .B(_11057_),
    .Y(_00033_));
 NAND2x1_ASAP7_75t_R _19266_ (.A(net6272),
    .B(_11029_),
    .Y(_11058_));
 NAND2x1_ASAP7_75t_R _19267_ (.A(net5528),
    .B(_10923_),
    .Y(_11059_));
 NAND2x1_ASAP7_75t_R _19268_ (.A(net5309),
    .B(net5307),
    .Y(_11060_));
 AND3x1_ASAP7_75t_R _19269_ (.A(net6283),
    .B(net6284),
    .C(_11060_),
    .Y(_11061_));
 OA21x2_ASAP7_75t_R _19270_ (.A1(_11059_),
    .A2(_11061_),
    .B(net6264),
    .Y(_11062_));
 OA21x2_ASAP7_75t_R _19271_ (.A1(net5216),
    .A2(_10912_),
    .B(net6264),
    .Y(_11063_));
 OA21x2_ASAP7_75t_R _19272_ (.A1(_10911_),
    .A2(_11063_),
    .B(net5219),
    .Y(_11064_));
 OAI21x1_ASAP7_75t_R _19273_ (.A1(_11058_),
    .A2(_11062_),
    .B(_11064_),
    .Y(_11065_));
 OA21x2_ASAP7_75t_R _19274_ (.A1(net6264),
    .A2(_01081_),
    .B(net6272),
    .Y(_11066_));
 OAI21x1_ASAP7_75t_R _19275_ (.A1(net5901),
    .A2(net5899),
    .B(net5909),
    .Y(_11067_));
 NAND2x1_ASAP7_75t_R _19276_ (.A(net6264),
    .B(_11067_),
    .Y(_11068_));
 AOI21x1_ASAP7_75t_R _19277_ (.A1(_11066_),
    .A2(_11068_),
    .B(net5219),
    .Y(_11069_));
 AOI22x1_ASAP7_75t_R _19278_ (.A1(net6281),
    .A2(net6282),
    .B1(net6283),
    .B2(net6284),
    .Y(_11070_));
 AOI21x1_ASAP7_75t_R _19279_ (.A1(net5909),
    .A2(_11070_),
    .B(net6264),
    .Y(_11071_));
 AND2x2_ASAP7_75t_R _19280_ (.A(net6264),
    .B(_01076_),
    .Y(_11072_));
 OR3x1_ASAP7_75t_R _19281_ (.A(_11071_),
    .B(net6272),
    .C(_11072_),
    .Y(_11073_));
 AOI21x1_ASAP7_75t_R _19282_ (.A1(_11069_),
    .A2(_11073_),
    .B(net5895),
    .Y(_11074_));
 NAND2x1_ASAP7_75t_R _19283_ (.A(_11065_),
    .B(_11074_),
    .Y(_11075_));
 NOR3x1_ASAP7_75t_R _19284_ (.A(_10956_),
    .B(net6277),
    .C(net5016),
    .Y(_11076_));
 NOR2x1_ASAP7_75t_R _19285_ (.A(net4960),
    .B(_10876_),
    .Y(_11077_));
 OAI21x1_ASAP7_75t_R _19286_ (.A1(_11076_),
    .A2(_11077_),
    .B(net6272),
    .Y(_11078_));
 NAND2x1_ASAP7_75t_R _19287_ (.A(_01079_),
    .B(net6273),
    .Y(_11079_));
 AOI21x1_ASAP7_75t_R _19288_ (.A1(net5900),
    .A2(net5892),
    .B(net6277),
    .Y(_11080_));
 AOI21x1_ASAP7_75t_R _19289_ (.A1(_11050_),
    .A2(_11080_),
    .B(net6271),
    .Y(_11081_));
 AOI21x1_ASAP7_75t_R _19290_ (.A1(_11079_),
    .A2(_11081_),
    .B(net5221),
    .Y(_11082_));
 NAND2x1_ASAP7_75t_R _19291_ (.A(_11078_),
    .B(_11082_),
    .Y(_11083_));
 AOI21x1_ASAP7_75t_R _19292_ (.A1(net5905),
    .A2(net5893),
    .B(net6274),
    .Y(_11084_));
 NAND2x1_ASAP7_75t_R _19293_ (.A(_10992_),
    .B(_11084_),
    .Y(_11085_));
 AOI21x1_ASAP7_75t_R _19294_ (.A1(net5896),
    .A2(net5910),
    .B(net6265),
    .Y(_11086_));
 AOI21x1_ASAP7_75t_R _19295_ (.A1(_11038_),
    .A2(_11086_),
    .B(net6267),
    .Y(_11087_));
 NAND2x1_ASAP7_75t_R _19296_ (.A(_11085_),
    .B(_11087_),
    .Y(_11088_));
 OA21x2_ASAP7_75t_R _19297_ (.A1(net6264),
    .A2(_01077_),
    .B(net6268),
    .Y(_11089_));
 OAI21x1_ASAP7_75t_R _19298_ (.A1(net5905),
    .A2(_11026_),
    .B(_10920_),
    .Y(_11090_));
 AOI21x1_ASAP7_75t_R _19299_ (.A1(_11090_),
    .A2(_11089_),
    .B(net5533),
    .Y(_11091_));
 AOI21x1_ASAP7_75t_R _19300_ (.A1(_11088_),
    .A2(_11091_),
    .B(net6278),
    .Y(_11092_));
 AOI21x1_ASAP7_75t_R _19301_ (.A1(_11092_),
    .A2(_11083_),
    .B(net6263),
    .Y(_11093_));
 NAND2x1_ASAP7_75t_R _19302_ (.A(_11093_),
    .B(_11075_),
    .Y(_11094_));
 NOR2x1_ASAP7_75t_R _19303_ (.A(_10791_),
    .B(net6264),
    .Y(_11095_));
 NAND2x1_ASAP7_75t_R _19304_ (.A(_10992_),
    .B(_11095_),
    .Y(_11096_));
 INVx2_ASAP7_75t_R _19305_ (.A(net4778),
    .Y(_11097_));
 AO21x1_ASAP7_75t_R _19306_ (.A1(_11097_),
    .A2(_10913_),
    .B(net6277),
    .Y(_11098_));
 AOI21x1_ASAP7_75t_R _19307_ (.A1(_11096_),
    .A2(_11098_),
    .B(_10875_),
    .Y(_11099_));
 NOR2x1_ASAP7_75t_R _19308_ (.A(net5903),
    .B(net5901),
    .Y(_11100_));
 AO21x1_ASAP7_75t_R _19309_ (.A1(net6283),
    .A2(net6284),
    .B(net5304),
    .Y(_11101_));
 NAND2x1_ASAP7_75t_R _19310_ (.A(net6276),
    .B(_11101_),
    .Y(_11102_));
 OAI21x1_ASAP7_75t_R _19311_ (.A1(_11100_),
    .A2(_11102_),
    .B(net6272),
    .Y(_11103_));
 NAND2x1_ASAP7_75t_R _19312_ (.A(net6265),
    .B(_10898_),
    .Y(_11104_));
 OAI21x1_ASAP7_75t_R _19313_ (.A1(_10931_),
    .A2(_11104_),
    .B(net5219),
    .Y(_11105_));
 OAI21x1_ASAP7_75t_R _19314_ (.A1(_11103_),
    .A2(_11105_),
    .B(net5895),
    .Y(_11106_));
 NOR2x1_ASAP7_75t_R _19315_ (.A(_11099_),
    .B(_11106_),
    .Y(_11107_));
 AO21x1_ASAP7_75t_R _19316_ (.A1(_10898_),
    .A2(net4959),
    .B(net6266),
    .Y(_11108_));
 AOI21x1_ASAP7_75t_R _19317_ (.A1(net5307),
    .A2(net5903),
    .B(net6274),
    .Y(_11109_));
 NAND2x1_ASAP7_75t_R _19318_ (.A(net5532),
    .B(_11109_),
    .Y(_11110_));
 AOI21x1_ASAP7_75t_R _19319_ (.A1(_11108_),
    .A2(_11110_),
    .B(_10784_),
    .Y(_11111_));
 AO21x1_ASAP7_75t_R _19320_ (.A1(_11101_),
    .A2(_10898_),
    .B(net6265),
    .Y(_11112_));
 AO21x1_ASAP7_75t_R _19321_ (.A1(net5530),
    .A2(net4959),
    .B(net6276),
    .Y(_11113_));
 AOI21x1_ASAP7_75t_R _19322_ (.A1(_11112_),
    .A2(_11113_),
    .B(net6268),
    .Y(_11114_));
 OAI21x1_ASAP7_75t_R _19323_ (.A1(_11111_),
    .A2(_11114_),
    .B(net5533),
    .Y(_11115_));
 AOI21x1_ASAP7_75t_R _19324_ (.A1(_11107_),
    .A2(_11115_),
    .B(_10868_),
    .Y(_11116_));
 INVx1_ASAP7_75t_R _19325_ (.A(_10961_),
    .Y(_11117_));
 AND2x2_ASAP7_75t_R _19326_ (.A(_11009_),
    .B(_11117_),
    .Y(_11118_));
 INVx1_ASAP7_75t_R _19327_ (.A(_11118_),
    .Y(_11119_));
 AOI21x1_ASAP7_75t_R _19328_ (.A1(_11068_),
    .A2(_11119_),
    .B(net6268),
    .Y(_11120_));
 OAI21x1_ASAP7_75t_R _19329_ (.A1(net5902),
    .A2(net5910),
    .B(net6266),
    .Y(_11121_));
 INVx1_ASAP7_75t_R _19330_ (.A(_10832_),
    .Y(_11122_));
 OAI21x1_ASAP7_75t_R _19331_ (.A1(_11121_),
    .A2(_11122_),
    .B(net6268),
    .Y(_11123_));
 OAI21x1_ASAP7_75t_R _19332_ (.A1(_10877_),
    .A2(_11123_),
    .B(net5533),
    .Y(_11124_));
 NOR2x1_ASAP7_75t_R _19333_ (.A(_11120_),
    .B(_11124_),
    .Y(_11125_));
 OAI21x1_ASAP7_75t_R _19334_ (.A1(net5309),
    .A2(net5899),
    .B(net6264),
    .Y(_11126_));
 NOR2x1_ASAP7_75t_R _19335_ (.A(_11100_),
    .B(_11126_),
    .Y(_11127_));
 AOI21x1_ASAP7_75t_R _19336_ (.A1(net4781),
    .A2(net5525),
    .B(net6266),
    .Y(_11128_));
 OAI21x1_ASAP7_75t_R _19337_ (.A1(_11127_),
    .A2(_11128_),
    .B(net6272),
    .Y(_11129_));
 NOR2x1_ASAP7_75t_R _19338_ (.A(net6272),
    .B(_11071_),
    .Y(_11130_));
 OAI21x1_ASAP7_75t_R _19339_ (.A1(net4958),
    .A2(_10981_),
    .B(_11130_),
    .Y(_11131_));
 AOI21x1_ASAP7_75t_R _19340_ (.A1(_11129_),
    .A2(_11131_),
    .B(net5533),
    .Y(_11132_));
 OAI21x1_ASAP7_75t_R _19341_ (.A1(_11125_),
    .A2(_11132_),
    .B(net6278),
    .Y(_11133_));
 NAND2x1_ASAP7_75t_R _19342_ (.A(_11116_),
    .B(_11133_),
    .Y(_11134_));
 NAND2x1_ASAP7_75t_R _19343_ (.A(_11134_),
    .B(_11094_),
    .Y(_00034_));
 NOR2x1_ASAP7_75t_R _19344_ (.A(_10956_),
    .B(_10842_),
    .Y(_11135_));
 AO21x1_ASAP7_75t_R _19345_ (.A1(_11135_),
    .A2(_11084_),
    .B(net6272),
    .Y(_11136_));
 AND2x2_ASAP7_75t_R _19346_ (.A(_10975_),
    .B(_10993_),
    .Y(_11137_));
 INVx1_ASAP7_75t_R _19347_ (.A(_10872_),
    .Y(_11138_));
 NOR2x1_ASAP7_75t_R _19348_ (.A(net4704),
    .B(net4592),
    .Y(_11139_));
 OAI22x1_ASAP7_75t_R _19349_ (.A1(_11136_),
    .A2(_11137_),
    .B1(_10948_),
    .B2(_11139_),
    .Y(_11140_));
 NOR2x1p5_ASAP7_75t_R _19350_ (.A(_10822_),
    .B(_10912_),
    .Y(_11141_));
 OA21x2_ASAP7_75t_R _19351_ (.A1(net5222),
    .A2(net5896),
    .B(_11141_),
    .Y(_11142_));
 NOR2x1_ASAP7_75t_R _19352_ (.A(_11142_),
    .B(_10979_),
    .Y(_11143_));
 OAI21x1_ASAP7_75t_R _19353_ (.A1(net5900),
    .A2(net5896),
    .B(_10818_),
    .Y(_11144_));
 NOR2x1_ASAP7_75t_R _19354_ (.A(_11144_),
    .B(_10944_),
    .Y(_11145_));
 INVx1_ASAP7_75t_R _19355_ (.A(_11023_),
    .Y(_11146_));
 AO21x1_ASAP7_75t_R _19356_ (.A1(_11145_),
    .A2(_11146_),
    .B(net5220),
    .Y(_11147_));
 OAI21x1_ASAP7_75t_R _19357_ (.A1(_11143_),
    .A2(_11147_),
    .B(net5895),
    .Y(_11148_));
 AOI21x1_ASAP7_75t_R _19358_ (.A1(net5220),
    .A2(_11140_),
    .B(_11148_),
    .Y(_11149_));
 AOI21x1_ASAP7_75t_R _19359_ (.A1(net4707),
    .A2(_11109_),
    .B(_11128_),
    .Y(_11150_));
 OAI21x1_ASAP7_75t_R _19360_ (.A1(_10875_),
    .A2(_11150_),
    .B(net6278),
    .Y(_11151_));
 NAND2x1_ASAP7_75t_R _19361_ (.A(net4956),
    .B(net4593),
    .Y(_11152_));
 AOI21x1_ASAP7_75t_R _19362_ (.A1(net6276),
    .A2(_11135_),
    .B(net5529),
    .Y(_11153_));
 NAND2x1_ASAP7_75t_R _19363_ (.A(_11152_),
    .B(_11153_),
    .Y(_11154_));
 NOR2x1p5_ASAP7_75t_R _19364_ (.A(_10931_),
    .B(net4595),
    .Y(_11155_));
 NOR2x1_ASAP7_75t_R _19365_ (.A(_10969_),
    .B(_10945_),
    .Y(_11156_));
 NOR2x1_ASAP7_75t_R _19366_ (.A(_10784_),
    .B(_10814_),
    .Y(_11157_));
 OAI21x1_ASAP7_75t_R _19367_ (.A1(_11155_),
    .A2(_11156_),
    .B(_11157_),
    .Y(_11158_));
 AOI21x1_ASAP7_75t_R _19368_ (.A1(net5530),
    .A2(net5525),
    .B(net6265),
    .Y(_11159_));
 NOR2x1_ASAP7_75t_R _19369_ (.A(_10818_),
    .B(_10814_),
    .Y(_11160_));
 OAI21x1_ASAP7_75t_R _19370_ (.A1(net4593),
    .A2(_11159_),
    .B(net4954),
    .Y(_11161_));
 NAND3x1_ASAP7_75t_R _19371_ (.A(_11158_),
    .B(_11154_),
    .C(_11161_),
    .Y(_11162_));
 OAI21x1_ASAP7_75t_R _19372_ (.A1(_11151_),
    .A2(_11162_),
    .B(_10868_),
    .Y(_11163_));
 AO21x1_ASAP7_75t_R _19373_ (.A1(net5211),
    .A2(net6265),
    .B(_11017_),
    .Y(_11164_));
 AO21x1_ASAP7_75t_R _19374_ (.A1(_11051_),
    .A2(net4781),
    .B(net5220),
    .Y(_11165_));
 AOI21x1_ASAP7_75t_R _19375_ (.A1(net4705),
    .A2(_11164_),
    .B(_11165_),
    .Y(_11166_));
 NOR2x1_ASAP7_75t_R _19376_ (.A(net6277),
    .B(_10898_),
    .Y(_11167_));
 NOR2x1_ASAP7_75t_R _19377_ (.A(net5533),
    .B(_11167_),
    .Y(_11168_));
 AO21x1_ASAP7_75t_R _19378_ (.A1(_11168_),
    .A2(_11096_),
    .B(_10784_),
    .Y(_11169_));
 NAND2x1_ASAP7_75t_R _19379_ (.A(net4778),
    .B(net6264),
    .Y(_11170_));
 NAND2x1_ASAP7_75t_R _19380_ (.A(_10824_),
    .B(_11050_),
    .Y(_11171_));
 INVx1_ASAP7_75t_R _19381_ (.A(_11160_),
    .Y(_11172_));
 AOI21x1_ASAP7_75t_R _19382_ (.A1(_11170_),
    .A2(_11171_),
    .B(_11172_),
    .Y(_11173_));
 NOR2x2_ASAP7_75t_R _19383_ (.A(net6264),
    .B(net4779),
    .Y(_11174_));
 AOI21x1_ASAP7_75t_R _19384_ (.A1(net5220),
    .A2(_11174_),
    .B(_10827_),
    .Y(_11175_));
 OAI21x1_ASAP7_75t_R _19385_ (.A1(_11175_),
    .A2(net6268),
    .B(net6278),
    .Y(_11176_));
 NOR2x1_ASAP7_75t_R _19386_ (.A(_11173_),
    .B(_11176_),
    .Y(_11177_));
 OAI21x1_ASAP7_75t_R _19387_ (.A1(_11166_),
    .A2(_11169_),
    .B(_11177_),
    .Y(_11178_));
 OAI21x1_ASAP7_75t_R _19388_ (.A1(net5905),
    .A2(net5210),
    .B(net4709),
    .Y(_11179_));
 INVx1_ASAP7_75t_R _19389_ (.A(_11157_),
    .Y(_11180_));
 AOI21x1_ASAP7_75t_R _19390_ (.A1(_11179_),
    .A2(_11029_),
    .B(_11180_),
    .Y(_11181_));
 OAI21x1_ASAP7_75t_R _19391_ (.A1(net5219),
    .A2(_11103_),
    .B(net5895),
    .Y(_11182_));
 NOR2x1_ASAP7_75t_R _19392_ (.A(_11181_),
    .B(_11182_),
    .Y(_11183_));
 AO21x1_ASAP7_75t_R _19393_ (.A1(_10891_),
    .A2(net5212),
    .B(net6275),
    .Y(_11184_));
 AO21x1_ASAP7_75t_R _19394_ (.A1(_11101_),
    .A2(_10913_),
    .B(net6265),
    .Y(_11185_));
 NAND3x1_ASAP7_75t_R _19395_ (.A(_11184_),
    .B(net6270),
    .C(_11185_),
    .Y(_11186_));
 OAI21x1_ASAP7_75t_R _19396_ (.A1(net5910),
    .A2(net5906),
    .B(_11086_),
    .Y(_11187_));
 AOI21x1_ASAP7_75t_R _19397_ (.A1(net6265),
    .A2(_10988_),
    .B(net6271),
    .Y(_11188_));
 AOI21x1_ASAP7_75t_R _19398_ (.A1(_11187_),
    .A2(_11188_),
    .B(net5533),
    .Y(_11189_));
 NAND2x1_ASAP7_75t_R _19399_ (.A(_11186_),
    .B(_11189_),
    .Y(_11190_));
 AOI21x1_ASAP7_75t_R _19400_ (.A1(_11183_),
    .A2(_11190_),
    .B(_10868_),
    .Y(_11191_));
 NAND2x1_ASAP7_75t_R _19401_ (.A(_11191_),
    .B(_11178_),
    .Y(_11192_));
 OAI21x1_ASAP7_75t_R _19402_ (.A1(_11149_),
    .A2(_11163_),
    .B(_11192_),
    .Y(_00035_));
 NOR2x1_ASAP7_75t_R _19403_ (.A(net6277),
    .B(_10796_),
    .Y(_11193_));
 AOI21x1_ASAP7_75t_R _19404_ (.A1(_10923_),
    .A2(_11193_),
    .B(net4527),
    .Y(_11194_));
 OAI21x1_ASAP7_75t_R _19405_ (.A1(_11172_),
    .A2(_11194_),
    .B(net6278),
    .Y(_11195_));
 OA21x2_ASAP7_75t_R _19406_ (.A1(_11038_),
    .A2(net6275),
    .B(net5212),
    .Y(_11196_));
 AO21x1_ASAP7_75t_R _19407_ (.A1(_11196_),
    .A2(_11001_),
    .B(net5533),
    .Y(_11197_));
 AO21x1_ASAP7_75t_R _19408_ (.A1(_11047_),
    .A2(_11097_),
    .B(net6272),
    .Y(_11198_));
 NOR2x1_ASAP7_75t_R _19409_ (.A(_10797_),
    .B(_11198_),
    .Y(_11199_));
 AOI21x1_ASAP7_75t_R _19410_ (.A1(net4956),
    .A2(net5525),
    .B(net6276),
    .Y(_11200_));
 OAI21x1_ASAP7_75t_R _19411_ (.A1(_11200_),
    .A2(_10839_),
    .B(_11157_),
    .Y(_11201_));
 OAI21x1_ASAP7_75t_R _19412_ (.A1(_11199_),
    .A2(_11197_),
    .B(_11201_),
    .Y(_11202_));
 OAI21x1_ASAP7_75t_R _19413_ (.A1(_11195_),
    .A2(_11202_),
    .B(_10868_),
    .Y(_11203_));
 AND3x1_ASAP7_75t_R _19414_ (.A(_10794_),
    .B(net6271),
    .C(_10826_),
    .Y(_11204_));
 AOI21x1_ASAP7_75t_R _19415_ (.A1(net5530),
    .A2(_10923_),
    .B(net6275),
    .Y(_11205_));
 OAI21x1_ASAP7_75t_R _19416_ (.A1(_10965_),
    .A2(_11021_),
    .B(net6267),
    .Y(_11206_));
 NOR2x1_ASAP7_75t_R _19417_ (.A(_11205_),
    .B(_11206_),
    .Y(_11207_));
 OAI21x1_ASAP7_75t_R _19418_ (.A1(_11204_),
    .A2(_11207_),
    .B(net5221),
    .Y(_11208_));
 OA21x2_ASAP7_75t_R _19419_ (.A1(_10938_),
    .A2(_10953_),
    .B(net4954),
    .Y(_11209_));
 INVx1_ASAP7_75t_R _19420_ (.A(_11121_),
    .Y(_11210_));
 NAND2x1_ASAP7_75t_R _19421_ (.A(_11020_),
    .B(_11210_),
    .Y(_11211_));
 AOI22x1_ASAP7_75t_R _19422_ (.A1(_11209_),
    .A2(_11211_),
    .B1(_11016_),
    .B2(_11081_),
    .Y(_11212_));
 AOI21x1_ASAP7_75t_R _19423_ (.A1(_11208_),
    .A2(_11212_),
    .B(net6278),
    .Y(_11213_));
 AOI21x1_ASAP7_75t_R _19424_ (.A1(net4777),
    .A2(net4706),
    .B(_10929_),
    .Y(_11214_));
 NAND2x1_ASAP7_75t_R _19425_ (.A(net6275),
    .B(_11046_),
    .Y(_11215_));
 AND2x2_ASAP7_75t_R _19426_ (.A(_11215_),
    .B(net6269),
    .Y(_11216_));
 AO21x1_ASAP7_75t_R _19427_ (.A1(_11216_),
    .A2(_10981_),
    .B(net5533),
    .Y(_11217_));
 OAI21x1_ASAP7_75t_R _19428_ (.A1(net5896),
    .A2(net5910),
    .B(_10986_),
    .Y(_11218_));
 NAND2x1_ASAP7_75t_R _19429_ (.A(net6275),
    .B(_11218_),
    .Y(_11219_));
 NAND2x1_ASAP7_75t_R _19430_ (.A(_11018_),
    .B(_11219_),
    .Y(_11220_));
 NOR2x1_ASAP7_75t_R _19431_ (.A(net6270),
    .B(_11025_),
    .Y(_11221_));
 AO21x1_ASAP7_75t_R _19432_ (.A1(_10992_),
    .A2(_11101_),
    .B(net6265),
    .Y(_11222_));
 AOI21x1_ASAP7_75t_R _19433_ (.A1(_11221_),
    .A2(_11222_),
    .B(net5221),
    .Y(_11223_));
 AOI21x1_ASAP7_75t_R _19434_ (.A1(_11220_),
    .A2(_11223_),
    .B(net6278),
    .Y(_11224_));
 OA21x2_ASAP7_75t_R _19435_ (.A1(_11214_),
    .A2(_11217_),
    .B(_11224_),
    .Y(_11225_));
 NOR2x1_ASAP7_75t_R _19436_ (.A(_10842_),
    .B(_10947_),
    .Y(_11226_));
 OAI21x1_ASAP7_75t_R _19437_ (.A1(_10881_),
    .A2(_11226_),
    .B(_11157_),
    .Y(_11227_));
 AOI21x1_ASAP7_75t_R _19438_ (.A1(net5530),
    .A2(net5532),
    .B(net6266),
    .Y(_11228_));
 NAND2x1_ASAP7_75t_R _19439_ (.A(_10793_),
    .B(net5531),
    .Y(_11229_));
 INVx1_ASAP7_75t_R _19440_ (.A(_11229_),
    .Y(_11230_));
 OAI21x1_ASAP7_75t_R _19441_ (.A1(_11228_),
    .A2(_11230_),
    .B(_10886_),
    .Y(_11231_));
 NAND2x1_ASAP7_75t_R _19442_ (.A(_11227_),
    .B(_11231_),
    .Y(_11232_));
 NOR2x1_ASAP7_75t_R _19443_ (.A(_11100_),
    .B(_10794_),
    .Y(_11233_));
 AOI21x1_ASAP7_75t_R _19444_ (.A1(net5526),
    .A2(net5531),
    .B(net6266),
    .Y(_11234_));
 OAI21x1_ASAP7_75t_R _19445_ (.A1(_11233_),
    .A2(_11234_),
    .B(net4954),
    .Y(_11235_));
 NAND2x1_ASAP7_75t_R _19446_ (.A(net5016),
    .B(net6265),
    .Y(_11236_));
 OA21x2_ASAP7_75t_R _19447_ (.A1(_01071_),
    .A2(net6266),
    .B(net5214),
    .Y(_11237_));
 AOI21x1_ASAP7_75t_R _19448_ (.A1(_11236_),
    .A2(_11237_),
    .B(net5895),
    .Y(_11238_));
 NAND2x1_ASAP7_75t_R _19449_ (.A(_11235_),
    .B(_11238_),
    .Y(_11239_));
 OAI21x1_ASAP7_75t_R _19450_ (.A1(_11232_),
    .A2(_11239_),
    .B(net6263),
    .Y(_11240_));
 OAI22x1_ASAP7_75t_R _19451_ (.A1(_11203_),
    .A2(_11213_),
    .B1(_11225_),
    .B2(_11240_),
    .Y(_00036_));
 NOR2x1_ASAP7_75t_R _19452_ (.A(net6265),
    .B(net5530),
    .Y(_11241_));
 NOR2x1_ASAP7_75t_R _19453_ (.A(_11241_),
    .B(_10895_),
    .Y(_11242_));
 AO21x1_ASAP7_75t_R _19454_ (.A1(_11138_),
    .A2(net6265),
    .B(net6268),
    .Y(_11243_));
 AOI21x1_ASAP7_75t_R _19455_ (.A1(net5209),
    .A2(_10975_),
    .B(net6265),
    .Y(_11244_));
 OAI21x1_ASAP7_75t_R _19456_ (.A1(_11243_),
    .A2(_11244_),
    .B(net5533),
    .Y(_11245_));
 NOR2x1_ASAP7_75t_R _19457_ (.A(_11242_),
    .B(_11245_),
    .Y(_11246_));
 AO21x1_ASAP7_75t_R _19458_ (.A1(net6265),
    .A2(net5906),
    .B(net6271),
    .Y(_11247_));
 OAI21x1_ASAP7_75t_R _19459_ (.A1(_11247_),
    .A2(_10946_),
    .B(net5220),
    .Y(_11248_));
 AO21x1_ASAP7_75t_R _19460_ (.A1(net5532),
    .A2(_11095_),
    .B(net6268),
    .Y(_11249_));
 NOR2x1_ASAP7_75t_R _19461_ (.A(net4595),
    .B(_10939_),
    .Y(_11250_));
 NOR2x1_ASAP7_75t_R _19462_ (.A(_11249_),
    .B(_11250_),
    .Y(_11251_));
 OAI21x1_ASAP7_75t_R _19463_ (.A1(_11248_),
    .A2(_11251_),
    .B(net5895),
    .Y(_11252_));
 OAI21x1_ASAP7_75t_R _19464_ (.A1(_11246_),
    .A2(_11252_),
    .B(net6263),
    .Y(_11253_));
 NOR2x1_ASAP7_75t_R _19465_ (.A(net6271),
    .B(_11164_),
    .Y(_11254_));
 AO21x1_ASAP7_75t_R _19466_ (.A1(_10964_),
    .A2(_10963_),
    .B(_10893_),
    .Y(_11255_));
 AO21x1_ASAP7_75t_R _19467_ (.A1(_11001_),
    .A2(_10978_),
    .B(net5533),
    .Y(_11256_));
 AOI21x1_ASAP7_75t_R _19468_ (.A1(_11254_),
    .A2(_11255_),
    .B(_11256_),
    .Y(_11257_));
 NOR2x1_ASAP7_75t_R _19469_ (.A(net5906),
    .B(net6265),
    .Y(_11258_));
 NOR2x1_ASAP7_75t_R _19470_ (.A(_11258_),
    .B(_11086_),
    .Y(_11259_));
 NAND2x1_ASAP7_75t_R _19471_ (.A(net5306),
    .B(net6265),
    .Y(_11260_));
 AO21x1_ASAP7_75t_R _19472_ (.A1(_11259_),
    .A2(_11260_),
    .B(_11180_),
    .Y(_11261_));
 NAND2x1_ASAP7_75t_R _19473_ (.A(net4705),
    .B(_11141_),
    .Y(_11262_));
 OAI21x1_ASAP7_75t_R _19474_ (.A1(net4594),
    .A2(net5218),
    .B(_11262_),
    .Y(_11263_));
 AOI21x1_ASAP7_75t_R _19475_ (.A1(net4954),
    .A2(_11263_),
    .B(net5895),
    .Y(_11264_));
 NAND2x1_ASAP7_75t_R _19476_ (.A(_11261_),
    .B(_11264_),
    .Y(_11265_));
 NOR2x1_ASAP7_75t_R _19477_ (.A(_11257_),
    .B(_11265_),
    .Y(_11266_));
 NAND2x1_ASAP7_75t_R _19478_ (.A(_10952_),
    .B(_11051_),
    .Y(_11267_));
 OAI21x1_ASAP7_75t_R _19479_ (.A1(net5218),
    .A2(_10893_),
    .B(net6265),
    .Y(_11268_));
 NAND2x1_ASAP7_75t_R _19480_ (.A(_11267_),
    .B(_11268_),
    .Y(_11269_));
 AO21x1_ASAP7_75t_R _19481_ (.A1(net5908),
    .A2(net6265),
    .B(net6269),
    .Y(_11270_));
 NOR2x1_ASAP7_75t_R _19482_ (.A(_10953_),
    .B(_10938_),
    .Y(_11271_));
 OAI21x1_ASAP7_75t_R _19483_ (.A1(_11270_),
    .A2(_11271_),
    .B(net5221),
    .Y(_11272_));
 AOI21x1_ASAP7_75t_R _19484_ (.A1(net6269),
    .A2(_11269_),
    .B(_11272_),
    .Y(_11273_));
 INVx1_ASAP7_75t_R _19485_ (.A(_11050_),
    .Y(_11274_));
 OAI21x1_ASAP7_75t_R _19486_ (.A1(_11215_),
    .A2(_11274_),
    .B(_11236_),
    .Y(_11275_));
 NAND2x1_ASAP7_75t_R _19487_ (.A(net4954),
    .B(_11275_),
    .Y(_11276_));
 NAND2x1p5_ASAP7_75t_R _19488_ (.A(_10914_),
    .B(_10905_),
    .Y(_11277_));
 AND2x2_ASAP7_75t_R _19489_ (.A(_11157_),
    .B(_11102_),
    .Y(_11278_));
 AOI21x1_ASAP7_75t_R _19490_ (.A1(_11277_),
    .A2(_11278_),
    .B(net5895),
    .Y(_11279_));
 NAND2x1_ASAP7_75t_R _19491_ (.A(_11276_),
    .B(_11279_),
    .Y(_11280_));
 OAI21x1_ASAP7_75t_R _19492_ (.A1(_11273_),
    .A2(_11280_),
    .B(_10868_),
    .Y(_11281_));
 AO21x1_ASAP7_75t_R _19493_ (.A1(_11026_),
    .A2(_11025_),
    .B(net4706),
    .Y(_11282_));
 NAND2x1_ASAP7_75t_R _19494_ (.A(net6270),
    .B(_11282_),
    .Y(_11283_));
 AO21x1_ASAP7_75t_R _19495_ (.A1(_11184_),
    .A2(_10954_),
    .B(net6270),
    .Y(_11284_));
 AOI21x1_ASAP7_75t_R _19496_ (.A1(_11283_),
    .A2(_11284_),
    .B(net5220),
    .Y(_11285_));
 NOR2x1_ASAP7_75t_R _19497_ (.A(net4957),
    .B(_10884_),
    .Y(_11286_));
 NOR2x1_ASAP7_75t_R _19498_ (.A(_11286_),
    .B(_10932_),
    .Y(_11287_));
 INVx1_ASAP7_75t_R _19499_ (.A(_11095_),
    .Y(_11288_));
 OAI21x1_ASAP7_75t_R _19500_ (.A1(net5213),
    .A2(_10756_),
    .B(net6266),
    .Y(_11289_));
 OAI21x1_ASAP7_75t_R _19501_ (.A1(_11288_),
    .A2(_10796_),
    .B(_11289_),
    .Y(_11290_));
 AOI21x1_ASAP7_75t_R _19502_ (.A1(_10886_),
    .A2(_11290_),
    .B(net6278),
    .Y(_11291_));
 OAI21x1_ASAP7_75t_R _19503_ (.A1(_10875_),
    .A2(_11287_),
    .B(_11291_),
    .Y(_11292_));
 NOR2x1_ASAP7_75t_R _19504_ (.A(_11285_),
    .B(_11292_),
    .Y(_11293_));
 OAI22x1_ASAP7_75t_R _19505_ (.A1(_11253_),
    .A2(_11266_),
    .B1(_11281_),
    .B2(_11293_),
    .Y(_00037_));
 AO21x1_ASAP7_75t_R _19506_ (.A1(_10842_),
    .A2(net6274),
    .B(net6268),
    .Y(_11294_));
 NOR2x1_ASAP7_75t_R _19507_ (.A(net5012),
    .B(_10978_),
    .Y(_11295_));
 AOI21x1_ASAP7_75t_R _19508_ (.A1(_01075_),
    .A2(net6264),
    .B(net6272),
    .Y(_11296_));
 NAND2x1_ASAP7_75t_R _19509_ (.A(_11095_),
    .B(net5532),
    .Y(_11297_));
 AOI21x1_ASAP7_75t_R _19510_ (.A1(_11296_),
    .A2(_11297_),
    .B(net5533),
    .Y(_11298_));
 OAI21x1_ASAP7_75t_R _19511_ (.A1(_11294_),
    .A2(_11295_),
    .B(_11298_),
    .Y(_11299_));
 INVx1_ASAP7_75t_R _19512_ (.A(_11123_),
    .Y(_11300_));
 AOI21x1_ASAP7_75t_R _19513_ (.A1(_10825_),
    .A2(_11229_),
    .B(net6268),
    .Y(_11301_));
 OAI21x1_ASAP7_75t_R _19514_ (.A1(_11300_),
    .A2(_11301_),
    .B(net5533),
    .Y(_11302_));
 AOI21x1_ASAP7_75t_R _19515_ (.A1(_11299_),
    .A2(_11302_),
    .B(net5895),
    .Y(_11303_));
 OA21x2_ASAP7_75t_R _19516_ (.A1(_11080_),
    .A2(_11047_),
    .B(_10987_),
    .Y(_11304_));
 AOI21x1_ASAP7_75t_R _19517_ (.A1(_10963_),
    .A2(_11145_),
    .B(net5533),
    .Y(_11305_));
 OAI21x1_ASAP7_75t_R _19518_ (.A1(net6267),
    .A2(_11304_),
    .B(_11305_),
    .Y(_11306_));
 AOI21x1_ASAP7_75t_R _19519_ (.A1(net6277),
    .A2(net5012),
    .B(_11167_),
    .Y(_11307_));
 OA21x2_ASAP7_75t_R _19520_ (.A1(_11005_),
    .A2(net5907),
    .B(net6268),
    .Y(_11308_));
 NAND2x1_ASAP7_75t_R _19521_ (.A(_11307_),
    .B(_11308_),
    .Y(_11309_));
 AOI21x1_ASAP7_75t_R _19522_ (.A1(net6266),
    .A2(net5525),
    .B(net6268),
    .Y(_11310_));
 NOR2x1_ASAP7_75t_R _19523_ (.A(net6266),
    .B(net5910),
    .Y(_11311_));
 OAI21x1_ASAP7_75t_R _19524_ (.A1(_11311_),
    .A2(_11051_),
    .B(_10992_),
    .Y(_11312_));
 AOI21x1_ASAP7_75t_R _19525_ (.A1(_11310_),
    .A2(_11312_),
    .B(net5219),
    .Y(_11313_));
 NAND2x1_ASAP7_75t_R _19526_ (.A(_11309_),
    .B(_11313_),
    .Y(_11314_));
 AOI21x1_ASAP7_75t_R _19527_ (.A1(_11306_),
    .A2(_11314_),
    .B(net6278),
    .Y(_11315_));
 OAI21x1_ASAP7_75t_R _19528_ (.A1(_11303_),
    .A2(_11315_),
    .B(net6263),
    .Y(_11316_));
 INVx1_ASAP7_75t_R _19529_ (.A(_11308_),
    .Y(_11317_));
 OAI21x1_ASAP7_75t_R _19530_ (.A1(net4778),
    .A2(_11061_),
    .B(net6274),
    .Y(_11318_));
 OAI21x1_ASAP7_75t_R _19531_ (.A1(_10842_),
    .A2(_10947_),
    .B(_11318_),
    .Y(_11319_));
 OA21x2_ASAP7_75t_R _19532_ (.A1(_10872_),
    .A2(net6266),
    .B(_10784_),
    .Y(_11320_));
 AO21x1_ASAP7_75t_R _19533_ (.A1(net5530),
    .A2(net5910),
    .B(net6277),
    .Y(_11321_));
 AOI21x1_ASAP7_75t_R _19534_ (.A1(_11320_),
    .A2(_11321_),
    .B(net5219),
    .Y(_11322_));
 OAI21x1_ASAP7_75t_R _19535_ (.A1(_11317_),
    .A2(_11319_),
    .B(_11322_),
    .Y(_11323_));
 NAND2x1p5_ASAP7_75t_R _19536_ (.A(_11046_),
    .B(_11141_),
    .Y(_11324_));
 OAI21x1_ASAP7_75t_R _19537_ (.A1(_11121_),
    .A2(_10939_),
    .B(_11324_),
    .Y(_11325_));
 AOI21x1_ASAP7_75t_R _19538_ (.A1(net5214),
    .A2(_11325_),
    .B(net5895),
    .Y(_11326_));
 NOR2x1p5_ASAP7_75t_R _19539_ (.A(net5529),
    .B(_11174_),
    .Y(_11327_));
 OAI21x1_ASAP7_75t_R _19540_ (.A1(_11071_),
    .A2(_11072_),
    .B(_11327_),
    .Y(_11328_));
 NAND3x1_ASAP7_75t_R _19541_ (.A(_11323_),
    .B(_11326_),
    .C(_11328_),
    .Y(_11329_));
 INVx1_ASAP7_75t_R _19542_ (.A(net5212),
    .Y(_11330_));
 AO21x1_ASAP7_75t_R _19543_ (.A1(_11330_),
    .A2(net6264),
    .B(net6268),
    .Y(_11331_));
 AO22x1_ASAP7_75t_R _19544_ (.A1(net6274),
    .A2(_10841_),
    .B1(_11025_),
    .B2(net5211),
    .Y(_11332_));
 AND2x2_ASAP7_75t_R _19545_ (.A(_01074_),
    .B(_01080_),
    .Y(_11333_));
 OA21x2_ASAP7_75t_R _19546_ (.A1(net6264),
    .A2(_11333_),
    .B(net6268),
    .Y(_11334_));
 NAND2x1_ASAP7_75t_R _19547_ (.A(_11026_),
    .B(_11084_),
    .Y(_11335_));
 AOI21x1_ASAP7_75t_R _19548_ (.A1(_11334_),
    .A2(_11335_),
    .B(net5533),
    .Y(_11336_));
 OAI21x1_ASAP7_75t_R _19549_ (.A1(_11331_),
    .A2(_11332_),
    .B(_11336_),
    .Y(_11337_));
 NAND2x1_ASAP7_75t_R _19550_ (.A(_11003_),
    .B(_11095_),
    .Y(_11338_));
 AOI21x1_ASAP7_75t_R _19551_ (.A1(net5526),
    .A2(_11025_),
    .B(_10827_),
    .Y(_11339_));
 AOI21x1_ASAP7_75t_R _19552_ (.A1(_11338_),
    .A2(_11339_),
    .B(_11180_),
    .Y(_11340_));
 NOR2x1_ASAP7_75t_R _19553_ (.A(_11126_),
    .B(_10900_),
    .Y(_11341_));
 AOI21x1_ASAP7_75t_R _19554_ (.A1(net6274),
    .A2(_11100_),
    .B(net5219),
    .Y(_11342_));
 NAND2x1_ASAP7_75t_R _19555_ (.A(_10850_),
    .B(_11342_),
    .Y(_11343_));
 OAI21x1_ASAP7_75t_R _19556_ (.A1(_11341_),
    .A2(_11343_),
    .B(net5895),
    .Y(_11344_));
 NOR2x1_ASAP7_75t_R _19557_ (.A(_11340_),
    .B(_11344_),
    .Y(_11345_));
 AOI21x1_ASAP7_75t_R _19558_ (.A1(_11337_),
    .A2(_11345_),
    .B(net6263),
    .Y(_11346_));
 NAND2x1_ASAP7_75t_R _19559_ (.A(_11329_),
    .B(_11346_),
    .Y(_11347_));
 NAND2x1_ASAP7_75t_R _19560_ (.A(_11316_),
    .B(_11347_),
    .Y(_00038_));
 OAI21x1_ASAP7_75t_R _19561_ (.A1(_11070_),
    .A2(_11218_),
    .B(net6264),
    .Y(_11348_));
 OA21x2_ASAP7_75t_R _19562_ (.A1(_10796_),
    .A2(_10964_),
    .B(net6271),
    .Y(_11349_));
 NOR2x1_ASAP7_75t_R _19563_ (.A(net6271),
    .B(_11047_),
    .Y(_11350_));
 AO21x1_ASAP7_75t_R _19564_ (.A1(_11350_),
    .A2(_11229_),
    .B(net5533),
    .Y(_11351_));
 AOI21x1_ASAP7_75t_R _19565_ (.A1(_11348_),
    .A2(_11349_),
    .B(_11351_),
    .Y(_11352_));
 AO21x1_ASAP7_75t_R _19566_ (.A1(_11085_),
    .A2(_11338_),
    .B(_11180_),
    .Y(_11353_));
 AOI22x1_ASAP7_75t_R _19567_ (.A1(_11051_),
    .A2(net4780),
    .B1(_10920_),
    .B2(_11003_),
    .Y(_11354_));
 OA21x2_ASAP7_75t_R _19568_ (.A1(_11354_),
    .A2(_11172_),
    .B(net5895),
    .Y(_11355_));
 NAND2x1_ASAP7_75t_R _19569_ (.A(_11353_),
    .B(_11355_),
    .Y(_11356_));
 NOR2x1_ASAP7_75t_R _19570_ (.A(_11352_),
    .B(_11356_),
    .Y(_11357_));
 AO21x1_ASAP7_75t_R _19571_ (.A1(net5904),
    .A2(_10953_),
    .B(_10938_),
    .Y(_11358_));
 AND2x2_ASAP7_75t_R _19572_ (.A(_11358_),
    .B(_11081_),
    .Y(_11359_));
 OAI21x1_ASAP7_75t_R _19573_ (.A1(_11258_),
    .A2(_11205_),
    .B(net6269),
    .Y(_11360_));
 NAND2x1_ASAP7_75t_R _19574_ (.A(net5221),
    .B(_11360_),
    .Y(_11361_));
 NOR2x1_ASAP7_75t_R _19575_ (.A(_11359_),
    .B(_11361_),
    .Y(_11362_));
 NOR2x1_ASAP7_75t_R _19576_ (.A(net6271),
    .B(_11174_),
    .Y(_11363_));
 AO21x1_ASAP7_75t_R _19577_ (.A1(_11363_),
    .A2(_11024_),
    .B(net5221),
    .Y(_11364_));
 NAND2x1_ASAP7_75t_R _19578_ (.A(net5904),
    .B(_10953_),
    .Y(_11365_));
 AOI211x1_ASAP7_75t_R _19579_ (.A1(_11365_),
    .A2(net4776),
    .B(_11193_),
    .C(net6267),
    .Y(_11366_));
 OAI21x1_ASAP7_75t_R _19580_ (.A1(_11364_),
    .A2(_11366_),
    .B(net6278),
    .Y(_11367_));
 OAI21x1_ASAP7_75t_R _19581_ (.A1(_11362_),
    .A2(_11367_),
    .B(net6263),
    .Y(_11368_));
 INVx1_ASAP7_75t_R _19582_ (.A(_01071_),
    .Y(_11369_));
 OAI21x1_ASAP7_75t_R _19583_ (.A1(_11369_),
    .A2(net6274),
    .B(_10847_),
    .Y(_11370_));
 AO21x1_ASAP7_75t_R _19584_ (.A1(net5530),
    .A2(net5910),
    .B(net6266),
    .Y(_11371_));
 NAND2x1_ASAP7_75t_R _19585_ (.A(_11371_),
    .B(_11018_),
    .Y(_11372_));
 AOI21x1_ASAP7_75t_R _19586_ (.A1(_11370_),
    .A2(_11372_),
    .B(net5533),
    .Y(_11373_));
 OA21x2_ASAP7_75t_R _19587_ (.A1(_01080_),
    .A2(net6274),
    .B(net5533),
    .Y(_11374_));
 AO21x1_ASAP7_75t_R _19588_ (.A1(net5212),
    .A2(_11097_),
    .B(net6264),
    .Y(_11375_));
 AOI21x1_ASAP7_75t_R _19589_ (.A1(_11374_),
    .A2(_11375_),
    .B(net4954),
    .Y(_11376_));
 NAND2x1_ASAP7_75t_R _19590_ (.A(_10913_),
    .B(_10920_),
    .Y(_11377_));
 NAND2x1_ASAP7_75t_R _19591_ (.A(net5531),
    .B(_11051_),
    .Y(_11378_));
 AOI21x1_ASAP7_75t_R _19592_ (.A1(_11377_),
    .A2(_11378_),
    .B(net6268),
    .Y(_11379_));
 OAI21x1_ASAP7_75t_R _19593_ (.A1(_11376_),
    .A2(_11379_),
    .B(net6278),
    .Y(_11380_));
 NOR2x1_ASAP7_75t_R _19594_ (.A(_11373_),
    .B(_11380_),
    .Y(_11381_));
 AO21x1_ASAP7_75t_R _19595_ (.A1(net6274),
    .A2(net5213),
    .B(net6268),
    .Y(_11382_));
 AO21x1_ASAP7_75t_R _19596_ (.A1(_11026_),
    .A2(_11084_),
    .B(_11382_),
    .Y(_11383_));
 AOI21x1_ASAP7_75t_R _19597_ (.A1(net5893),
    .A2(_11025_),
    .B(_10841_),
    .Y(_11384_));
 AOI21x1_ASAP7_75t_R _19598_ (.A1(_10847_),
    .A2(_11384_),
    .B(net5220),
    .Y(_11385_));
 NAND2x1_ASAP7_75t_R _19599_ (.A(_11383_),
    .B(_11385_),
    .Y(_11386_));
 AO21x1_ASAP7_75t_R _19600_ (.A1(net5528),
    .A2(net5910),
    .B(net6265),
    .Y(_11387_));
 AOI21x1_ASAP7_75t_R _19601_ (.A1(_11179_),
    .A2(_11387_),
    .B(net5529),
    .Y(_11388_));
 OAI21x1_ASAP7_75t_R _19602_ (.A1(net4594),
    .A2(_11138_),
    .B(net5214),
    .Y(_11389_));
 NOR2x1_ASAP7_75t_R _19603_ (.A(_10964_),
    .B(_11218_),
    .Y(_11390_));
 NOR2x1_ASAP7_75t_R _19604_ (.A(_11390_),
    .B(_11389_),
    .Y(_11391_));
 NOR2x1_ASAP7_75t_R _19605_ (.A(_11388_),
    .B(_11391_),
    .Y(_11392_));
 AOI21x1_ASAP7_75t_R _19606_ (.A1(_11386_),
    .A2(_11392_),
    .B(net6278),
    .Y(_11393_));
 OAI21x1_ASAP7_75t_R _19607_ (.A1(_11393_),
    .A2(_11381_),
    .B(_10868_),
    .Y(_11394_));
 OAI21x1_ASAP7_75t_R _19608_ (.A1(_11357_),
    .A2(_11368_),
    .B(_11394_),
    .Y(_00039_));
 NOR2x1_ASAP7_75t_R _19609_ (.A(net6669),
    .B(_00447_),
    .Y(_11395_));
 XOR2x2_ASAP7_75t_R _19610_ (.A(_00590_),
    .B(_00583_),
    .Y(_11396_));
 XOR2x2_ASAP7_75t_R _19611_ (.A(net6615),
    .B(net6591),
    .Y(_11397_));
 XOR2x2_ASAP7_75t_R _19612_ (.A(_11396_),
    .B(_11397_),
    .Y(_11398_));
 XOR2x2_ASAP7_75t_R _19613_ (.A(_00615_),
    .B(_00622_),
    .Y(_11399_));
 XOR2x2_ASAP7_75t_R _19614_ (.A(_11399_),
    .B(net6558),
    .Y(_11400_));
 XOR2x2_ASAP7_75t_R _19615_ (.A(_11398_),
    .B(_11400_),
    .Y(_11401_));
 NOR2x1p5_ASAP7_75t_R _19616_ (.A(net6463),
    .B(_11401_),
    .Y(_11402_));
 OAI21x1_ASAP7_75t_R _19617_ (.A1(_11395_),
    .A2(net6363),
    .B(net6502),
    .Y(_11403_));
 AND2x2_ASAP7_75t_R _19618_ (.A(net6463),
    .B(_00447_),
    .Y(_11404_));
 XNOR2x2_ASAP7_75t_R _19619_ (.A(_11400_),
    .B(_11398_),
    .Y(_11405_));
 NOR2x1p5_ASAP7_75t_R _19620_ (.A(net6463),
    .B(_11405_),
    .Y(_11406_));
 INVx1_ASAP7_75t_R _19621_ (.A(net6502),
    .Y(_11407_));
 OAI21x1_ASAP7_75t_R _19622_ (.A1(_11404_),
    .A2(net6362),
    .B(_11407_),
    .Y(_11408_));
 NAND2x1_ASAP7_75t_R _19623_ (.A(_11403_),
    .B(_11408_),
    .Y(_11409_));
 INVx1_ASAP7_75t_R _19625_ (.A(net6559),
    .Y(_11410_));
 XOR2x2_ASAP7_75t_R _19626_ (.A(net6640),
    .B(net6614),
    .Y(_11411_));
 NAND2x1_ASAP7_75t_R _19627_ (.A(_11410_),
    .B(_11411_),
    .Y(_11412_));
 XNOR2x2_ASAP7_75t_R _19628_ (.A(net6640),
    .B(net6614),
    .Y(_11413_));
 NAND2x1_ASAP7_75t_R _19629_ (.A(net6559),
    .B(_11413_),
    .Y(_11414_));
 XOR2x2_ASAP7_75t_R _19630_ (.A(_00647_),
    .B(_00615_),
    .Y(_11415_));
 INVx1_ASAP7_75t_R _19631_ (.A(net6442),
    .Y(_11416_));
 AOI21x1_ASAP7_75t_R _19632_ (.A1(_11412_),
    .A2(_11414_),
    .B(_11416_),
    .Y(_11417_));
 NAND2x1_ASAP7_75t_R _19633_ (.A(net6559),
    .B(_11411_),
    .Y(_11418_));
 NAND2x1_ASAP7_75t_R _19634_ (.A(_11410_),
    .B(_11413_),
    .Y(_11419_));
 AOI21x1_ASAP7_75t_R _19635_ (.A1(_11418_),
    .A2(_11419_),
    .B(net6442),
    .Y(_11420_));
 OAI21x1_ASAP7_75t_R _19636_ (.A1(_11417_),
    .A2(_11420_),
    .B(net6669),
    .Y(_11421_));
 NOR2x1_ASAP7_75t_R _19637_ (.A(net6668),
    .B(_00448_),
    .Y(_11422_));
 INVx1_ASAP7_75t_R _19638_ (.A(_11422_),
    .Y(_11423_));
 NAND3x1_ASAP7_75t_R _19639_ (.A(_11421_),
    .B(_08987_),
    .C(_11423_),
    .Y(_11424_));
 AO21x1_ASAP7_75t_R _19640_ (.A1(_11421_),
    .A2(_11423_),
    .B(_08987_),
    .Y(_11425_));
 NAND2x1_ASAP7_75t_R _19641_ (.A(_11424_),
    .B(_11425_),
    .Y(_11426_));
 INVx1_ASAP7_75t_R _19643_ (.A(_00617_),
    .Y(_11427_));
 XOR2x2_ASAP7_75t_R _19644_ (.A(_00584_),
    .B(_00616_),
    .Y(_11428_));
 NAND2x1_ASAP7_75t_R _19645_ (.A(_11427_),
    .B(net6441),
    .Y(_11429_));
 XNOR2x2_ASAP7_75t_R _19646_ (.A(_00616_),
    .B(_00584_),
    .Y(_11430_));
 NAND2x1_ASAP7_75t_R _19647_ (.A(_00617_),
    .B(_11430_),
    .Y(_11431_));
 XNOR2x2_ASAP7_75t_R _19648_ (.A(net6589),
    .B(net6557),
    .Y(_11432_));
 AOI21x1_ASAP7_75t_R _19649_ (.A1(_11429_),
    .A2(_11431_),
    .B(_11432_),
    .Y(_11433_));
 NAND2x1_ASAP7_75t_R _19650_ (.A(_00617_),
    .B(net6441),
    .Y(_11434_));
 NAND2x1_ASAP7_75t_R _19651_ (.A(_11427_),
    .B(_11430_),
    .Y(_11435_));
 XOR2x2_ASAP7_75t_R _19652_ (.A(_00649_),
    .B(_00681_),
    .Y(_11436_));
 AOI21x1_ASAP7_75t_R _19653_ (.A1(_11434_),
    .A2(_11435_),
    .B(_11436_),
    .Y(_11437_));
 OAI21x1_ASAP7_75t_R _19654_ (.A1(_11433_),
    .A2(_11437_),
    .B(net6669),
    .Y(_11438_));
 NOR2x1_ASAP7_75t_R _19655_ (.A(net6669),
    .B(_00449_),
    .Y(_11439_));
 INVx1_ASAP7_75t_R _19656_ (.A(_11439_),
    .Y(_11440_));
 NAND3x1_ASAP7_75t_R _19657_ (.A(_11438_),
    .B(net6501),
    .C(_11440_),
    .Y(_11441_));
 AO21x1_ASAP7_75t_R _19658_ (.A1(_11438_),
    .A2(_11440_),
    .B(net6501),
    .Y(_11442_));
 NAND2x2_ASAP7_75t_R _19659_ (.A(_11441_),
    .B(_11442_),
    .Y(_11443_));
 NAND3x1_ASAP7_75t_R _19661_ (.A(_11421_),
    .B(net6503),
    .C(_11423_),
    .Y(_11444_));
 AO21x1_ASAP7_75t_R _19662_ (.A1(_11421_),
    .A2(_11423_),
    .B(net6503),
    .Y(_11445_));
 NAND2x1p5_ASAP7_75t_R _19663_ (.A(_11444_),
    .B(_11445_),
    .Y(_11446_));
 INVx1_ASAP7_75t_R _19665_ (.A(_11438_),
    .Y(_11447_));
 OAI21x1_ASAP7_75t_R _19666_ (.A1(_11439_),
    .A2(_11447_),
    .B(net6501),
    .Y(_11448_));
 NAND3x1_ASAP7_75t_R _19668_ (.A(_11438_),
    .B(_08797_),
    .C(_11440_),
    .Y(_11450_));
 NAND2x1_ASAP7_75t_R _19670_ (.A(_11448_),
    .B(_11450_),
    .Y(_11452_));
 XOR2x2_ASAP7_75t_R _19673_ (.A(_00588_),
    .B(_00620_),
    .Y(_11454_));
 XOR2x2_ASAP7_75t_R _19674_ (.A(_00621_),
    .B(_00653_),
    .Y(_11455_));
 XOR2x2_ASAP7_75t_R _19675_ (.A(_11455_),
    .B(_00685_),
    .Y(_11456_));
 XNOR2x2_ASAP7_75t_R _19676_ (.A(_11454_),
    .B(_11456_),
    .Y(_11457_));
 NOR2x1_ASAP7_75t_R _19681_ (.A(net6667),
    .B(_00491_),
    .Y(_11462_));
 AO21x1_ASAP7_75t_R _19682_ (.A1(_11457_),
    .A2(net6667),
    .B(_11462_),
    .Y(_11463_));
 XOR2x2_ASAP7_75t_R _19683_ (.A(_11463_),
    .B(_00893_),
    .Y(_11464_));
 INVx1_ASAP7_75t_R _19684_ (.A(_11464_),
    .Y(_11465_));
 NOR2x1_ASAP7_75t_R _19686_ (.A(net5303),
    .B(_11443_),
    .Y(_11467_));
 XOR2x2_ASAP7_75t_R _19687_ (.A(_00585_),
    .B(net6640),
    .Y(_11468_));
 XNOR2x2_ASAP7_75t_R _19688_ (.A(_00618_),
    .B(_11468_),
    .Y(_11469_));
 XNOR2x2_ASAP7_75t_R _19689_ (.A(_00650_),
    .B(_00682_),
    .Y(_11470_));
 XOR2x2_ASAP7_75t_R _19690_ (.A(_00617_),
    .B(net6614),
    .Y(_11471_));
 XOR2x2_ASAP7_75t_R _19691_ (.A(_11470_),
    .B(_11471_),
    .Y(_11472_));
 NOR2x1_ASAP7_75t_R _19692_ (.A(_11469_),
    .B(_11472_),
    .Y(_11473_));
 AO21x1_ASAP7_75t_R _19693_ (.A1(_11472_),
    .A2(_11469_),
    .B(net6463),
    .Y(_11474_));
 NAND2x1_ASAP7_75t_R _19694_ (.A(_00494_),
    .B(net6463),
    .Y(_11475_));
 OAI21x1_ASAP7_75t_R _19695_ (.A1(_11473_),
    .A2(_11474_),
    .B(_11475_),
    .Y(_11476_));
 XNOR2x2_ASAP7_75t_R _19696_ (.A(net6500),
    .B(_11476_),
    .Y(_11477_));
 XOR2x2_ASAP7_75t_R _19699_ (.A(_00586_),
    .B(net6640),
    .Y(_11480_));
 XNOR2x2_ASAP7_75t_R _19700_ (.A(_00619_),
    .B(_11480_),
    .Y(_11481_));
 XOR2x2_ASAP7_75t_R _19701_ (.A(_00618_),
    .B(net6614),
    .Y(_11482_));
 XOR2x2_ASAP7_75t_R _19702_ (.A(_00651_),
    .B(_00683_),
    .Y(_11483_));
 XNOR2x2_ASAP7_75t_R _19703_ (.A(_11482_),
    .B(_11483_),
    .Y(_11484_));
 NOR2x1_ASAP7_75t_R _19704_ (.A(_11481_),
    .B(_11484_),
    .Y(_11485_));
 AO21x1_ASAP7_75t_R _19705_ (.A1(_11484_),
    .A2(_11481_),
    .B(net6463),
    .Y(_11486_));
 AND2x2_ASAP7_75t_R _19706_ (.A(net6461),
    .B(_00493_),
    .Y(_11487_));
 INVx1_ASAP7_75t_R _19707_ (.A(_11487_),
    .Y(_11488_));
 OAI21x1_ASAP7_75t_R _19708_ (.A1(_11485_),
    .A2(_11486_),
    .B(_11488_),
    .Y(_11489_));
 XOR2x2_ASAP7_75t_R _19709_ (.A(_11489_),
    .B(_00890_),
    .Y(_11490_));
 AO21x1_ASAP7_75t_R _19712_ (.A1(_11467_),
    .A2(net6252),
    .B(net6249),
    .Y(_11493_));
 INVx1_ASAP7_75t_R _19715_ (.A(_01091_),
    .Y(_11496_));
 AOI21x1_ASAP7_75t_R _19716_ (.A1(net6260),
    .A2(net6259),
    .B(_11496_),
    .Y(_11497_));
 NOR2x1_ASAP7_75t_R _19717_ (.A(_11497_),
    .B(net6252),
    .Y(_11498_));
 INVx1_ASAP7_75t_R _19718_ (.A(_11498_),
    .Y(_11499_));
 AOI211x1_ASAP7_75t_R _19720_ (.A1(net6261),
    .A2(net6262),
    .B(_11443_),
    .C(net5887),
    .Y(_11501_));
 NOR2x1_ASAP7_75t_R _19721_ (.A(_11499_),
    .B(_11501_),
    .Y(_11502_));
 XOR2x2_ASAP7_75t_R _19722_ (.A(_00587_),
    .B(_00619_),
    .Y(_11503_));
 XOR2x2_ASAP7_75t_R _19723_ (.A(_00620_),
    .B(_00652_),
    .Y(_11504_));
 XOR2x2_ASAP7_75t_R _19724_ (.A(_11504_),
    .B(net6555),
    .Y(_11505_));
 NOR2x1_ASAP7_75t_R _19725_ (.A(_11503_),
    .B(_11505_),
    .Y(_11506_));
 XNOR2x2_ASAP7_75t_R _19726_ (.A(_00587_),
    .B(_00619_),
    .Y(_11507_));
 INVx1_ASAP7_75t_R _19727_ (.A(_00684_),
    .Y(_11508_));
 XOR2x2_ASAP7_75t_R _19728_ (.A(_11504_),
    .B(_11508_),
    .Y(_11509_));
 NOR2x1_ASAP7_75t_R _19729_ (.A(_11507_),
    .B(_11509_),
    .Y(_11510_));
 OAI21x1_ASAP7_75t_R _19732_ (.A1(_11506_),
    .A2(_11510_),
    .B(net6667),
    .Y(_11513_));
 INVx1_ASAP7_75t_R _19733_ (.A(_00891_),
    .Y(_11514_));
 NOR2x1_ASAP7_75t_R _19734_ (.A(net6667),
    .B(_00492_),
    .Y(_11515_));
 INVx1_ASAP7_75t_R _19735_ (.A(_11515_),
    .Y(_11516_));
 NAND3x1_ASAP7_75t_R _19736_ (.A(_11513_),
    .B(_11514_),
    .C(_11516_),
    .Y(_11517_));
 AO21x1_ASAP7_75t_R _19737_ (.A1(_11513_),
    .A2(_11516_),
    .B(_11514_),
    .Y(_11518_));
 NAND2x1_ASAP7_75t_R _19738_ (.A(_11517_),
    .B(_11518_),
    .Y(_11519_));
 OAI21x1_ASAP7_75t_R _19741_ (.A1(_11493_),
    .A2(_11502_),
    .B(net5879),
    .Y(_11522_));
 XNOR2x2_ASAP7_75t_R _19742_ (.A(_00890_),
    .B(_11489_),
    .Y(_11523_));
 AOI21x1_ASAP7_75t_R _19746_ (.A1(net6260),
    .A2(net6259),
    .B(_01090_),
    .Y(_11527_));
 XOR2x2_ASAP7_75t_R _19747_ (.A(_11476_),
    .B(net6500),
    .Y(_11528_));
 NOR2x1_ASAP7_75t_R _19749_ (.A(_11527_),
    .B(net6246),
    .Y(_11530_));
 INVx1_ASAP7_75t_R _19750_ (.A(_11530_),
    .Y(_11531_));
 AO21x1_ASAP7_75t_R _19752_ (.A1(net6258),
    .A2(net5881),
    .B(net5303),
    .Y(_11533_));
 NOR2x1_ASAP7_75t_R _19753_ (.A(net6253),
    .B(_11533_),
    .Y(_11534_));
 INVx1_ASAP7_75t_R _19754_ (.A(_11534_),
    .Y(_11535_));
 OAI21x1_ASAP7_75t_R _19755_ (.A1(_11531_),
    .A2(_11501_),
    .B(_11535_),
    .Y(_11536_));
 NOR2x1_ASAP7_75t_R _19756_ (.A(net6248),
    .B(_11536_),
    .Y(_11537_));
 INVx1_ASAP7_75t_R _19759_ (.A(_01084_),
    .Y(_11540_));
 AOI21x1_ASAP7_75t_R _19760_ (.A1(net5881),
    .A2(net6258),
    .B(_11540_),
    .Y(_11541_));
 AOI21x1_ASAP7_75t_R _19761_ (.A1(net5888),
    .A2(net5885),
    .B(net4952),
    .Y(_11542_));
 AOI21x1_ASAP7_75t_R _19762_ (.A1(net6260),
    .A2(net6259),
    .B(net5303),
    .Y(_11543_));
 AOI21x1_ASAP7_75t_R _19765_ (.A1(net5208),
    .A2(net6253),
    .B(net6249),
    .Y(_11546_));
 OAI21x1_ASAP7_75t_R _19766_ (.A1(net6252),
    .A2(_11542_),
    .B(_11546_),
    .Y(_11547_));
 AOI21x1_ASAP7_75t_R _19768_ (.A1(net6260),
    .A2(net6259),
    .B(net5302),
    .Y(_11549_));
 AOI21x1_ASAP7_75t_R _19769_ (.A1(net5887),
    .A2(net5524),
    .B(_11549_),
    .Y(_11550_));
 OAI21x1_ASAP7_75t_R _19770_ (.A1(_11395_),
    .A2(_11402_),
    .B(_11407_),
    .Y(_11551_));
 OAI21x1_ASAP7_75t_R _19771_ (.A1(_11404_),
    .A2(_11406_),
    .B(net6502),
    .Y(_11552_));
 NAND2x1p5_ASAP7_75t_R _19772_ (.A(_11551_),
    .B(_11552_),
    .Y(_11553_));
 NAND2x1_ASAP7_75t_R _19773_ (.A(net5524),
    .B(net5877),
    .Y(_11554_));
 AOI21x1_ASAP7_75t_R _19775_ (.A1(_11550_),
    .A2(net5206),
    .B(net6244),
    .Y(_11556_));
 AOI21x1_ASAP7_75t_R _19776_ (.A1(net6260),
    .A2(net6259),
    .B(net5258),
    .Y(_11557_));
 AOI21x1_ASAP7_75t_R _19777_ (.A1(net5011),
    .A2(net6254),
    .B(net6247),
    .Y(_11558_));
 OR2x2_ASAP7_75t_R _19778_ (.A(_01098_),
    .B(net6254),
    .Y(_11559_));
 AOI21x1_ASAP7_75t_R _19780_ (.A1(_11558_),
    .A2(_11559_),
    .B(_11519_),
    .Y(_11561_));
 OAI21x1_ASAP7_75t_R _19781_ (.A1(_11547_),
    .A2(_11556_),
    .B(_11561_),
    .Y(_11562_));
 OAI21x1_ASAP7_75t_R _19782_ (.A1(_11522_),
    .A2(_11537_),
    .B(_11562_),
    .Y(_11563_));
 XNOR2x2_ASAP7_75t_R _19783_ (.A(_00589_),
    .B(_00621_),
    .Y(_11564_));
 INVx1_ASAP7_75t_R _19784_ (.A(net6554),
    .Y(_11565_));
 XOR2x2_ASAP7_75t_R _19785_ (.A(_11564_),
    .B(net6440),
    .Y(_11566_));
 XNOR2x2_ASAP7_75t_R _19786_ (.A(net6614),
    .B(net6587),
    .Y(_11567_));
 XOR2x2_ASAP7_75t_R _19787_ (.A(_11566_),
    .B(_11567_),
    .Y(_11568_));
 NOR2x1_ASAP7_75t_R _19788_ (.A(net6667),
    .B(_00490_),
    .Y(_11569_));
 AO21x1_ASAP7_75t_R _19789_ (.A1(_11568_),
    .A2(net6667),
    .B(_11569_),
    .Y(_11570_));
 XOR2x2_ASAP7_75t_R _19790_ (.A(_11570_),
    .B(_00894_),
    .Y(_11571_));
 INVx1_ASAP7_75t_R _19791_ (.A(_11571_),
    .Y(_11572_));
 OAI21x1_ASAP7_75t_R _19792_ (.A1(net5880),
    .A2(_11563_),
    .B(_11572_),
    .Y(_11573_));
 NAND3x1_ASAP7_75t_R _19793_ (.A(_11513_),
    .B(_00891_),
    .C(_11516_),
    .Y(_11574_));
 AO21x1_ASAP7_75t_R _19794_ (.A1(_11513_),
    .A2(_11516_),
    .B(_00891_),
    .Y(_11575_));
 NAND2x1_ASAP7_75t_R _19795_ (.A(_11574_),
    .B(_11575_),
    .Y(_11576_));
 OAI21x1_ASAP7_75t_R _19797_ (.A1(net5887),
    .A2(net5524),
    .B(net6244),
    .Y(_11578_));
 INVx1_ASAP7_75t_R _19798_ (.A(_11578_),
    .Y(_11579_));
 NAND3x1_ASAP7_75t_R _19799_ (.A(net5889),
    .B(net5888),
    .C(net5524),
    .Y(_11580_));
 AO21x1_ASAP7_75t_R _19800_ (.A1(net6256),
    .A2(_11549_),
    .B(net6249),
    .Y(_11581_));
 AOI21x1_ASAP7_75t_R _19801_ (.A1(_11579_),
    .A2(_11580_),
    .B(_11581_),
    .Y(_11582_));
 NAND2x1_ASAP7_75t_R _19802_ (.A(net5875),
    .B(_11582_),
    .Y(_11583_));
 OAI21x1_ASAP7_75t_R _19804_ (.A1(net5883),
    .A2(net5877),
    .B(net6252),
    .Y(_11584_));
 NOR2x1_ASAP7_75t_R _19805_ (.A(net5010),
    .B(_11584_),
    .Y(_11585_));
 NOR2x1_ASAP7_75t_R _19806_ (.A(net5882),
    .B(_11443_),
    .Y(_11586_));
 INVx1_ASAP7_75t_R _19807_ (.A(_01090_),
    .Y(_11587_));
 AO21x1_ASAP7_75t_R _19808_ (.A1(net6259),
    .A2(net6260),
    .B(_11587_),
    .Y(_11588_));
 INVx1_ASAP7_75t_R _19809_ (.A(_11588_),
    .Y(_11589_));
 NOR2x1_ASAP7_75t_R _19810_ (.A(net5522),
    .B(_11589_),
    .Y(_11590_));
 NOR2x1_ASAP7_75t_R _19811_ (.A(_11490_),
    .B(_11576_),
    .Y(_11591_));
 OAI21x1_ASAP7_75t_R _19812_ (.A1(net6253),
    .A2(_11590_),
    .B(_11591_),
    .Y(_11592_));
 NOR2x1_ASAP7_75t_R _19813_ (.A(_11585_),
    .B(_11592_),
    .Y(_11593_));
 INVx1_ASAP7_75t_R _19814_ (.A(_01085_),
    .Y(_11594_));
 AOI21x1_ASAP7_75t_R _19815_ (.A1(net5881),
    .A2(net6258),
    .B(_11594_),
    .Y(_11595_));
 INVx2_ASAP7_75t_R _19816_ (.A(_11595_),
    .Y(_11596_));
 NAND2x2_ASAP7_75t_R _19817_ (.A(_11596_),
    .B(net6246),
    .Y(_11597_));
 AOI21x1_ASAP7_75t_R _19818_ (.A1(_11549_),
    .A2(net6252),
    .B(net6248),
    .Y(_11598_));
 NAND2x1p5_ASAP7_75t_R _19819_ (.A(_11598_),
    .B(net4481),
    .Y(_11599_));
 NOR2x1_ASAP7_75t_R _19820_ (.A(net5300),
    .B(net5886),
    .Y(_11600_));
 AO21x1_ASAP7_75t_R _19822_ (.A1(_11600_),
    .A2(net6254),
    .B(net5879),
    .Y(_11602_));
 AOI21x1_ASAP7_75t_R _19823_ (.A1(net6260),
    .A2(net6259),
    .B(_11540_),
    .Y(_11603_));
 OA21x2_ASAP7_75t_R _19824_ (.A1(_11467_),
    .A2(net4950),
    .B(net6252),
    .Y(_11604_));
 NOR2x1_ASAP7_75t_R _19825_ (.A(net6248),
    .B(_11576_),
    .Y(_11605_));
 INVx1_ASAP7_75t_R _19826_ (.A(net5302),
    .Y(_11606_));
 OAI21x1_ASAP7_75t_R _19828_ (.A1(net5204),
    .A2(net5885),
    .B(net6244),
    .Y(_11608_));
 NAND2x1_ASAP7_75t_R _19829_ (.A(_11605_),
    .B(_11608_),
    .Y(_11609_));
 OAI22x1_ASAP7_75t_R _19830_ (.A1(_11599_),
    .A2(_11602_),
    .B1(_11604_),
    .B2(_11609_),
    .Y(_11610_));
 NOR2x1_ASAP7_75t_R _19831_ (.A(_11593_),
    .B(_11610_),
    .Y(_11611_));
 AOI21x1_ASAP7_75t_R _19834_ (.A1(_11583_),
    .A2(_11611_),
    .B(net6257),
    .Y(_11614_));
 AOI21x1_ASAP7_75t_R _19837_ (.A1(net5881),
    .A2(net6258),
    .B(net5258),
    .Y(_11617_));
 AOI21x1_ASAP7_75t_R _19838_ (.A1(_11443_),
    .A2(net5889),
    .B(net5009),
    .Y(_11618_));
 AO21x1_ASAP7_75t_R _19839_ (.A1(net6259),
    .A2(net6260),
    .B(_11594_),
    .Y(_11619_));
 INVx1_ASAP7_75t_R _19840_ (.A(_11619_),
    .Y(_11620_));
 NAND2x1_ASAP7_75t_R _19841_ (.A(net6244),
    .B(_11620_),
    .Y(_11621_));
 OAI21x1_ASAP7_75t_R _19842_ (.A1(net6244),
    .A2(_11618_),
    .B(_11621_),
    .Y(_11622_));
 OAI21x1_ASAP7_75t_R _19843_ (.A1(net6247),
    .A2(_11622_),
    .B(net5875),
    .Y(_11623_));
 INVx1_ASAP7_75t_R _19844_ (.A(_11541_),
    .Y(_11624_));
 AO21x1_ASAP7_75t_R _19845_ (.A1(net4951),
    .A2(_11624_),
    .B(net6244),
    .Y(_11625_));
 INVx1_ASAP7_75t_R _19847_ (.A(_11603_),
    .Y(_11627_));
 INVx1_ASAP7_75t_R _19848_ (.A(_11617_),
    .Y(_11628_));
 AO21x1_ASAP7_75t_R _19849_ (.A1(_11627_),
    .A2(net4771),
    .B(net6255),
    .Y(_11629_));
 AND3x1_ASAP7_75t_R _19850_ (.A(_11625_),
    .B(net6247),
    .C(_11629_),
    .Y(_11630_));
 OAI21x1_ASAP7_75t_R _19851_ (.A1(_11623_),
    .A2(_11630_),
    .B(net6257),
    .Y(_11631_));
 NAND2x1_ASAP7_75t_R _19853_ (.A(net5882),
    .B(net5877),
    .Y(_11633_));
 NOR2x1_ASAP7_75t_R _19854_ (.A(net6244),
    .B(_11586_),
    .Y(_11634_));
 NAND2x1_ASAP7_75t_R _19855_ (.A(_11633_),
    .B(_11634_),
    .Y(_11635_));
 NAND2x1_ASAP7_75t_R _19856_ (.A(net5887),
    .B(_11443_),
    .Y(_11636_));
 AOI21x1_ASAP7_75t_R _19857_ (.A1(net5882),
    .A2(net5891),
    .B(net6252),
    .Y(_11637_));
 NAND2x1_ASAP7_75t_R _19858_ (.A(_11636_),
    .B(_11637_),
    .Y(_11638_));
 AND2x2_ASAP7_75t_R _19859_ (.A(_11635_),
    .B(_11638_),
    .Y(_11639_));
 INVx1_ASAP7_75t_R _19860_ (.A(net6262),
    .Y(_11640_));
 INVx1_ASAP7_75t_R _19861_ (.A(net6261),
    .Y(_11641_));
 OAI21x1_ASAP7_75t_R _19862_ (.A1(_11640_),
    .A2(_11641_),
    .B(net5887),
    .Y(_11642_));
 NOR2x1_ASAP7_75t_R _19864_ (.A(net4775),
    .B(net6244),
    .Y(_11644_));
 OA21x2_ASAP7_75t_R _19865_ (.A1(_11642_),
    .A2(net5524),
    .B(_11644_),
    .Y(_11645_));
 AO21x1_ASAP7_75t_R _19867_ (.A1(net6258),
    .A2(net5881),
    .B(_11587_),
    .Y(_11647_));
 AO21x1_ASAP7_75t_R _19868_ (.A1(_11647_),
    .A2(_11627_),
    .B(net6255),
    .Y(_11648_));
 NAND2x1_ASAP7_75t_R _19869_ (.A(net6247),
    .B(_11648_),
    .Y(_11649_));
 OAI21x1_ASAP7_75t_R _19870_ (.A1(_11645_),
    .A2(_11649_),
    .B(net5879),
    .Y(_11650_));
 AOI21x1_ASAP7_75t_R _19871_ (.A1(net6249),
    .A2(_11639_),
    .B(_11650_),
    .Y(_11651_));
 NOR2x1_ASAP7_75t_R _19872_ (.A(_11631_),
    .B(_11651_),
    .Y(_11652_));
 INVx1_ASAP7_75t_R _19873_ (.A(_01093_),
    .Y(_11653_));
 AO21x1_ASAP7_75t_R _19874_ (.A1(net6258),
    .A2(net5881),
    .B(_11653_),
    .Y(_11654_));
 INVx1_ASAP7_75t_R _19876_ (.A(_11654_),
    .Y(_11656_));
 OAI21x1_ASAP7_75t_R _19877_ (.A1(_11656_),
    .A2(_11578_),
    .B(net6249),
    .Y(_11657_));
 NAND2x1_ASAP7_75t_R _19878_ (.A(net6251),
    .B(net5877),
    .Y(_11658_));
 OAI21x1_ASAP7_75t_R _19879_ (.A1(net5887),
    .A2(net5523),
    .B(net6252),
    .Y(_11659_));
 NOR2x1_ASAP7_75t_R _19880_ (.A(net5883),
    .B(net5891),
    .Y(_11660_));
 AOI21x1_ASAP7_75t_R _19881_ (.A1(_11658_),
    .A2(_11659_),
    .B(_11660_),
    .Y(_11661_));
 OAI21x1_ASAP7_75t_R _19883_ (.A1(_11657_),
    .A2(_11661_),
    .B(net5875),
    .Y(_11663_));
 AOI21x1_ASAP7_75t_R _19884_ (.A1(net6243),
    .A2(net6242),
    .B(_11452_),
    .Y(_11664_));
 OAI21x1_ASAP7_75t_R _19885_ (.A1(_11467_),
    .A2(_11664_),
    .B(net6256),
    .Y(_11665_));
 INVx1_ASAP7_75t_R _19886_ (.A(_11665_),
    .Y(_11666_));
 AOI211x1_ASAP7_75t_R _19887_ (.A1(net6261),
    .A2(net6262),
    .B(_11443_),
    .C(net5882),
    .Y(_11667_));
 OAI21x1_ASAP7_75t_R _19888_ (.A1(_11578_),
    .A2(_11667_),
    .B(net6247),
    .Y(_11668_));
 NOR2x1_ASAP7_75t_R _19889_ (.A(_11666_),
    .B(_11668_),
    .Y(_11669_));
 NOR2x1_ASAP7_75t_R _19890_ (.A(_11663_),
    .B(_11669_),
    .Y(_11670_));
 NAND2x1_ASAP7_75t_R _19891_ (.A(net6248),
    .B(_11659_),
    .Y(_11671_));
 NOR2x1_ASAP7_75t_R _19892_ (.A(net5523),
    .B(net5877),
    .Y(_11672_));
 AOI21x1_ASAP7_75t_R _19893_ (.A1(net5882),
    .A2(_11672_),
    .B(_11608_),
    .Y(_11673_));
 OAI21x1_ASAP7_75t_R _19894_ (.A1(_11671_),
    .A2(_11673_),
    .B(net5879),
    .Y(_11674_));
 AO21x1_ASAP7_75t_R _19895_ (.A1(net6259),
    .A2(net6260),
    .B(_11653_),
    .Y(_11675_));
 NAND2x1_ASAP7_75t_R _19896_ (.A(net6244),
    .B(_11675_),
    .Y(_11676_));
 OAI21x1_ASAP7_75t_R _19897_ (.A1(net4773),
    .A2(_11676_),
    .B(net6249),
    .Y(_11677_));
 NAND2x1_ASAP7_75t_R _19898_ (.A(net5523),
    .B(net5882),
    .Y(_11678_));
 INVx1_ASAP7_75t_R _19899_ (.A(_11678_),
    .Y(_11679_));
 NAND2x1_ASAP7_75t_R _19900_ (.A(net5882),
    .B(net5883),
    .Y(_11680_));
 OAI21x1_ASAP7_75t_R _19901_ (.A1(net5877),
    .A2(_11680_),
    .B(net6252),
    .Y(_11681_));
 NOR2x1_ASAP7_75t_R _19902_ (.A(_11679_),
    .B(_11681_),
    .Y(_11682_));
 NOR2x1_ASAP7_75t_R _19903_ (.A(_11677_),
    .B(_11682_),
    .Y(_11683_));
 OAI21x1_ASAP7_75t_R _19904_ (.A1(_11674_),
    .A2(_11683_),
    .B(net5880),
    .Y(_11684_));
 OAI21x1_ASAP7_75t_R _19905_ (.A1(_11670_),
    .A2(_11684_),
    .B(_11571_),
    .Y(_11685_));
 OAI22x1_ASAP7_75t_R _19906_ (.A1(_11573_),
    .A2(_11614_),
    .B1(_11652_),
    .B2(_11685_),
    .Y(_00040_));
 INVx1_ASAP7_75t_R _19907_ (.A(_11598_),
    .Y(_11686_));
 OAI21x1_ASAP7_75t_R _19908_ (.A1(net6252),
    .A2(_11672_),
    .B(net5206),
    .Y(_11687_));
 OAI21x1_ASAP7_75t_R _19909_ (.A1(_11686_),
    .A2(_11687_),
    .B(net5876),
    .Y(_11688_));
 AO21x1_ASAP7_75t_R _19910_ (.A1(net6258),
    .A2(net5881),
    .B(net5299),
    .Y(_11689_));
 INVx1_ASAP7_75t_R _19911_ (.A(_11689_),
    .Y(_11690_));
 OAI21x1_ASAP7_75t_R _19912_ (.A1(net5011),
    .A2(_11690_),
    .B(net6245),
    .Y(_11691_));
 NAND2x1_ASAP7_75t_R _19913_ (.A(net6248),
    .B(_11691_),
    .Y(_11692_));
 NOR2x1_ASAP7_75t_R _19914_ (.A(_11556_),
    .B(_11692_),
    .Y(_11693_));
 OAI21x1_ASAP7_75t_R _19915_ (.A1(_11688_),
    .A2(_11693_),
    .B(net6257),
    .Y(_11694_));
 AOI21x1_ASAP7_75t_R _19916_ (.A1(net5881),
    .A2(net6258),
    .B(_11606_),
    .Y(_11695_));
 NOR2x1_ASAP7_75t_R _19917_ (.A(_11695_),
    .B(net6244),
    .Y(_11696_));
 NOR2x1_ASAP7_75t_R _19918_ (.A(net4775),
    .B(net6256),
    .Y(_11697_));
 AOI221x1_ASAP7_75t_R _19919_ (.A1(net5521),
    .A2(net4702),
    .B1(_11680_),
    .B2(net4588),
    .C(net6248),
    .Y(_11698_));
 NAND2x1_ASAP7_75t_R _19920_ (.A(net5886),
    .B(net6245),
    .Y(_11699_));
 OAI21x1_ASAP7_75t_R _19921_ (.A1(_11640_),
    .A2(_11641_),
    .B(net5882),
    .Y(_11700_));
 INVx1_ASAP7_75t_R _19922_ (.A(_11700_),
    .Y(_11701_));
 NOR2x1_ASAP7_75t_R _19923_ (.A(_11699_),
    .B(_11701_),
    .Y(_11702_));
 NOR2x1_ASAP7_75t_R _19924_ (.A(net5887),
    .B(net5891),
    .Y(_11703_));
 OAI21x1_ASAP7_75t_R _19925_ (.A1(_11703_),
    .A2(_11584_),
    .B(net6248),
    .Y(_11704_));
 OAI21x1_ASAP7_75t_R _19926_ (.A1(_11702_),
    .A2(_11704_),
    .B(net5879),
    .Y(_11705_));
 NOR2x1_ASAP7_75t_R _19927_ (.A(_11698_),
    .B(_11705_),
    .Y(_11706_));
 OAI21x1_ASAP7_75t_R _19928_ (.A1(net5524),
    .A2(_11642_),
    .B(net6244),
    .Y(_11707_));
 INVx1_ASAP7_75t_R _19929_ (.A(_11707_),
    .Y(_11708_));
 NOR2x1_ASAP7_75t_R _19930_ (.A(net5302),
    .B(net5884),
    .Y(_11709_));
 AO21x1_ASAP7_75t_R _19931_ (.A1(_11709_),
    .A2(net6255),
    .B(net6249),
    .Y(_11710_));
 AOI21x1_ASAP7_75t_R _19932_ (.A1(net4771),
    .A2(_11708_),
    .B(_11710_),
    .Y(_11711_));
 OAI21x1_ASAP7_75t_R _19933_ (.A1(_11660_),
    .A2(_11676_),
    .B(net6249),
    .Y(_11712_));
 AOI21x1_ASAP7_75t_R _19934_ (.A1(net5888),
    .A2(net5889),
    .B(net5886),
    .Y(_11713_));
 INVx1_ASAP7_75t_R _19935_ (.A(_11713_),
    .Y(_11714_));
 NOR2x1_ASAP7_75t_R _19936_ (.A(net6244),
    .B(_11714_),
    .Y(_11715_));
 OAI21x1_ASAP7_75t_R _19937_ (.A1(_11712_),
    .A2(_11715_),
    .B(net5879),
    .Y(_11716_));
 NOR2x1_ASAP7_75t_R _19938_ (.A(_11711_),
    .B(_11716_),
    .Y(_11717_));
 OAI21x1_ASAP7_75t_R _19939_ (.A1(net4774),
    .A2(net5207),
    .B(net6245),
    .Y(_11718_));
 OAI21x1_ASAP7_75t_R _19940_ (.A1(net6245),
    .A2(_11542_),
    .B(_11718_),
    .Y(_11719_));
 OAI21x1_ASAP7_75t_R _19941_ (.A1(net6248),
    .A2(_11719_),
    .B(net5875),
    .Y(_11720_));
 AOI21x1_ASAP7_75t_R _19942_ (.A1(_11678_),
    .A2(net5520),
    .B(net6253),
    .Y(_11721_));
 NOR2x1_ASAP7_75t_R _19943_ (.A(net5011),
    .B(net6246),
    .Y(_11722_));
 AO21x1_ASAP7_75t_R _19944_ (.A1(_11722_),
    .A2(_11678_),
    .B(net6249),
    .Y(_11723_));
 NOR2x1_ASAP7_75t_R _19945_ (.A(_11721_),
    .B(_11723_),
    .Y(_11724_));
 OAI21x1_ASAP7_75t_R _19946_ (.A1(_11720_),
    .A2(_11724_),
    .B(net5880),
    .Y(_11725_));
 OAI22x1_ASAP7_75t_R _19947_ (.A1(_11694_),
    .A2(_11706_),
    .B1(_11717_),
    .B2(_11725_),
    .Y(_11726_));
 INVx1_ASAP7_75t_R _19948_ (.A(_11664_),
    .Y(_11727_));
 NOR2x1_ASAP7_75t_R _19949_ (.A(_11695_),
    .B(net6256),
    .Y(_11728_));
 AO21x1_ASAP7_75t_R _19950_ (.A1(_11727_),
    .A2(_11728_),
    .B(net6247),
    .Y(_11729_));
 AO21x1_ASAP7_75t_R _19951_ (.A1(net6262),
    .A2(net6261),
    .B(net5523),
    .Y(_11730_));
 AO21x1_ASAP7_75t_R _19952_ (.A1(_11634_),
    .A2(_11730_),
    .B(net5879),
    .Y(_11731_));
 NOR2x1_ASAP7_75t_R _19953_ (.A(_11729_),
    .B(_11731_),
    .Y(_11732_));
 AO21x1_ASAP7_75t_R _19954_ (.A1(net6259),
    .A2(net6260),
    .B(_01084_),
    .Y(_11733_));
 INVx1_ASAP7_75t_R _19955_ (.A(_11733_),
    .Y(_11734_));
 NAND2x1_ASAP7_75t_R _19956_ (.A(net6251),
    .B(_11678_),
    .Y(_11735_));
 NOR2x1_ASAP7_75t_R _19957_ (.A(_11734_),
    .B(_11735_),
    .Y(_11736_));
 NOR2x1_ASAP7_75t_R _19958_ (.A(net5883),
    .B(net6251),
    .Y(_11737_));
 NAND2x1_ASAP7_75t_R _19959_ (.A(_11642_),
    .B(_11737_),
    .Y(_11738_));
 NOR2x1_ASAP7_75t_R _19960_ (.A(net5523),
    .B(net6252),
    .Y(_11739_));
 NAND2x1_ASAP7_75t_R _19961_ (.A(net6249),
    .B(net5879),
    .Y(_11740_));
 AOI21x1_ASAP7_75t_R _19962_ (.A1(_11739_),
    .A2(net5519),
    .B(_11740_),
    .Y(_11741_));
 NAND2x1_ASAP7_75t_R _19963_ (.A(_11738_),
    .B(_11741_),
    .Y(_11742_));
 INVx1_ASAP7_75t_R _19964_ (.A(_01100_),
    .Y(_11743_));
 AOI21x1_ASAP7_75t_R _19965_ (.A1(_11574_),
    .A2(_11575_),
    .B(_11743_),
    .Y(_11744_));
 AOI21x1_ASAP7_75t_R _19966_ (.A1(net6244),
    .A2(_11744_),
    .B(net6249),
    .Y(_11745_));
 OAI21x1_ASAP7_75t_R _19967_ (.A1(net5883),
    .A2(_11642_),
    .B(_11530_),
    .Y(_11746_));
 AOI21x1_ASAP7_75t_R _19968_ (.A1(_11745_),
    .A2(_11746_),
    .B(_11465_),
    .Y(_11747_));
 OAI21x1_ASAP7_75t_R _19969_ (.A1(_11736_),
    .A2(_11742_),
    .B(_11747_),
    .Y(_11748_));
 OAI21x1_ASAP7_75t_R _19970_ (.A1(_11732_),
    .A2(_11748_),
    .B(_11571_),
    .Y(_11749_));
 INVx1_ASAP7_75t_R _19971_ (.A(_11543_),
    .Y(_11750_));
 NAND2x1_ASAP7_75t_R _19972_ (.A(_11750_),
    .B(_11689_),
    .Y(_11751_));
 AOI21x1_ASAP7_75t_R _19973_ (.A1(net6256),
    .A2(_11751_),
    .B(net6247),
    .Y(_11752_));
 OAI21x1_ASAP7_75t_R _19974_ (.A1(net5009),
    .A2(_11707_),
    .B(_11752_),
    .Y(_11753_));
 NOR2x1_ASAP7_75t_R _19975_ (.A(net6249),
    .B(_11697_),
    .Y(_11754_));
 NAND2x1_ASAP7_75t_R _19976_ (.A(net5523),
    .B(net5891),
    .Y(_11755_));
 AOI21x1_ASAP7_75t_R _19977_ (.A1(net5882),
    .A2(net5884),
    .B(net6244),
    .Y(_11756_));
 OAI21x1_ASAP7_75t_R _19978_ (.A1(net5882),
    .A2(net5201),
    .B(_11756_),
    .Y(_11757_));
 AOI21x1_ASAP7_75t_R _19979_ (.A1(_11754_),
    .A2(_11757_),
    .B(net5879),
    .Y(_11758_));
 NAND2x1_ASAP7_75t_R _19980_ (.A(_11753_),
    .B(_11758_),
    .Y(_11759_));
 NOR2x1_ASAP7_75t_R _19981_ (.A(net5523),
    .B(net5882),
    .Y(_11760_));
 OAI21x1_ASAP7_75t_R _19982_ (.A1(_11467_),
    .A2(_11760_),
    .B(net6256),
    .Y(_11761_));
 INVx1_ASAP7_75t_R _19983_ (.A(net5011),
    .Y(_11762_));
 AO21x1_ASAP7_75t_R _19984_ (.A1(_11762_),
    .A2(_11624_),
    .B(net6255),
    .Y(_11763_));
 AOI21x1_ASAP7_75t_R _19985_ (.A1(_11761_),
    .A2(_11763_),
    .B(net6247),
    .Y(_11764_));
 NAND2x1_ASAP7_75t_R _19986_ (.A(_11728_),
    .B(_11727_),
    .Y(_11765_));
 OAI21x1_ASAP7_75t_R _19987_ (.A1(net4950),
    .A2(_11679_),
    .B(net6256),
    .Y(_11766_));
 AOI21x1_ASAP7_75t_R _19988_ (.A1(_11765_),
    .A2(_11766_),
    .B(net6249),
    .Y(_11767_));
 OAI21x1_ASAP7_75t_R _19989_ (.A1(_11764_),
    .A2(_11767_),
    .B(net5879),
    .Y(_11768_));
 AOI21x1_ASAP7_75t_R _19990_ (.A1(_11759_),
    .A2(_11768_),
    .B(net6257),
    .Y(_11769_));
 NOR2x1_ASAP7_75t_R _19991_ (.A(_11749_),
    .B(_11769_),
    .Y(_11770_));
 AOI21x1_ASAP7_75t_R _19992_ (.A1(_11572_),
    .A2(_11726_),
    .B(_11770_),
    .Y(_00041_));
 NAND2x1_ASAP7_75t_R _19993_ (.A(net4949),
    .B(_11708_),
    .Y(_11771_));
 AND2x2_ASAP7_75t_R _19994_ (.A(_11681_),
    .B(_11591_),
    .Y(_11772_));
 NAND2x1_ASAP7_75t_R _19995_ (.A(net6256),
    .B(_11628_),
    .Y(_11773_));
 AO21x1_ASAP7_75t_R _19996_ (.A1(net5877),
    .A2(net5883),
    .B(_11773_),
    .Y(_11774_));
 OR3x1_ASAP7_75t_R _19997_ (.A(net5522),
    .B(net6253),
    .C(net5208),
    .Y(_11775_));
 AOI21x1_ASAP7_75t_R _19998_ (.A1(_11774_),
    .A2(_11775_),
    .B(_11740_),
    .Y(_11776_));
 AOI21x1_ASAP7_75t_R _19999_ (.A1(_11771_),
    .A2(_11772_),
    .B(_11776_),
    .Y(_11777_));
 NAND2x1_ASAP7_75t_R _20000_ (.A(net4948),
    .B(_11696_),
    .Y(_11778_));
 NAND2x1_ASAP7_75t_R _20001_ (.A(_11755_),
    .B(_11637_),
    .Y(_11779_));
 NAND2x1_ASAP7_75t_R _20002_ (.A(_11778_),
    .B(_11779_),
    .Y(_11780_));
 AOI21x1_ASAP7_75t_R _20003_ (.A1(net6249),
    .A2(_11780_),
    .B(net5879),
    .Y(_11781_));
 INVx1_ASAP7_75t_R _20004_ (.A(_11585_),
    .Y(_11782_));
 AND2x2_ASAP7_75t_R _20005_ (.A(net5206),
    .B(_11550_),
    .Y(_11783_));
 AOI21x1_ASAP7_75t_R _20006_ (.A1(net6244),
    .A2(_11783_),
    .B(net6250),
    .Y(_11784_));
 NAND2x1_ASAP7_75t_R _20007_ (.A(_11782_),
    .B(_11784_),
    .Y(_11785_));
 NAND2x1_ASAP7_75t_R _20008_ (.A(_11781_),
    .B(_11785_),
    .Y(_11786_));
 AOI21x1_ASAP7_75t_R _20009_ (.A1(_11777_),
    .A2(_11786_),
    .B(_11465_),
    .Y(_11787_));
 NOR2x1_ASAP7_75t_R _20010_ (.A(_11497_),
    .B(net6246),
    .Y(_11788_));
 NAND2x1_ASAP7_75t_R _20011_ (.A(_11678_),
    .B(_11788_),
    .Y(_11789_));
 NAND2x1_ASAP7_75t_R _20012_ (.A(_11762_),
    .B(_11697_),
    .Y(_11790_));
 AOI21x1_ASAP7_75t_R _20013_ (.A1(_11789_),
    .A2(_11790_),
    .B(net6249),
    .Y(_11791_));
 AO21x1_ASAP7_75t_R _20014_ (.A1(net6258),
    .A2(net5881),
    .B(_01091_),
    .Y(_11792_));
 NAND2x1_ASAP7_75t_R _20015_ (.A(net6246),
    .B(_11792_),
    .Y(_11793_));
 NOR2x1_ASAP7_75t_R _20016_ (.A(_11664_),
    .B(_11793_),
    .Y(_11794_));
 AO21x1_ASAP7_75t_R _20017_ (.A1(net6259),
    .A2(net6260),
    .B(net5299),
    .Y(_11795_));
 NAND2x1_ASAP7_75t_R _20018_ (.A(net6254),
    .B(_11795_),
    .Y(_11796_));
 OAI21x1_ASAP7_75t_R _20019_ (.A1(net5522),
    .A2(_11796_),
    .B(net6249),
    .Y(_11797_));
 NOR2x1_ASAP7_75t_R _20020_ (.A(_11794_),
    .B(_11797_),
    .Y(_11798_));
 OAI21x1_ASAP7_75t_R _20021_ (.A1(_11791_),
    .A2(_11798_),
    .B(net5879),
    .Y(_11799_));
 OAI21x1_ASAP7_75t_R _20022_ (.A1(net5207),
    .A2(net5522),
    .B(net6246),
    .Y(_11800_));
 AO21x1_ASAP7_75t_R _20023_ (.A1(_11795_),
    .A2(net5200),
    .B(net6246),
    .Y(_11801_));
 AOI21x1_ASAP7_75t_R _20024_ (.A1(_11800_),
    .A2(_11801_),
    .B(net6247),
    .Y(_11802_));
 INVx1_ASAP7_75t_R _20025_ (.A(_11549_),
    .Y(_11803_));
 AO21x1_ASAP7_75t_R _20026_ (.A1(net5200),
    .A2(_11803_),
    .B(net6246),
    .Y(_11804_));
 AOI21x1_ASAP7_75t_R _20027_ (.A1(net5302),
    .A2(net5884),
    .B(net6256),
    .Y(_11805_));
 NAND2x1_ASAP7_75t_R _20028_ (.A(net5205),
    .B(_11805_),
    .Y(_11806_));
 AOI21x1_ASAP7_75t_R _20029_ (.A1(_11804_),
    .A2(_11806_),
    .B(net6249),
    .Y(_11807_));
 OAI21x1_ASAP7_75t_R _20030_ (.A1(_11802_),
    .A2(_11807_),
    .B(net5875),
    .Y(_11808_));
 NAND2x1_ASAP7_75t_R _20031_ (.A(_11799_),
    .B(_11808_),
    .Y(_11809_));
 OAI21x1_ASAP7_75t_R _20032_ (.A1(net6257),
    .A2(_11809_),
    .B(_11571_),
    .Y(_11810_));
 AND3x1_ASAP7_75t_R _20033_ (.A(_11647_),
    .B(_11762_),
    .C(net6244),
    .Y(_11811_));
 NOR2x1_ASAP7_75t_R _20034_ (.A(net4950),
    .B(_11584_),
    .Y(_11812_));
 OAI21x1_ASAP7_75t_R _20035_ (.A1(_11811_),
    .A2(_11812_),
    .B(net6249),
    .Y(_11813_));
 AOI21x1_ASAP7_75t_R _20036_ (.A1(net5523),
    .A2(net5891),
    .B(net6251),
    .Y(_11814_));
 NOR2x1_ASAP7_75t_R _20037_ (.A(_11743_),
    .B(net6244),
    .Y(_11815_));
 AOI21x1_ASAP7_75t_R _20038_ (.A1(_11633_),
    .A2(_11814_),
    .B(_11815_),
    .Y(_11816_));
 AOI21x1_ASAP7_75t_R _20039_ (.A1(net6248),
    .A2(_11816_),
    .B(net5879),
    .Y(_11817_));
 NAND2x1_ASAP7_75t_R _20040_ (.A(_11813_),
    .B(_11817_),
    .Y(_11818_));
 NAND2x1_ASAP7_75t_R _20041_ (.A(net5888),
    .B(net6245),
    .Y(_11819_));
 AO21x1_ASAP7_75t_R _20042_ (.A1(_11819_),
    .A2(_11699_),
    .B(_11664_),
    .Y(_11820_));
 AOI21x1_ASAP7_75t_R _20043_ (.A1(net5524),
    .A2(net5889),
    .B(net5011),
    .Y(_11821_));
 AOI21x1_ASAP7_75t_R _20044_ (.A1(net6254),
    .A2(_11821_),
    .B(net6247),
    .Y(_11822_));
 NAND2x1_ASAP7_75t_R _20045_ (.A(_11820_),
    .B(_11822_),
    .Y(_11823_));
 OA21x2_ASAP7_75t_R _20046_ (.A1(net6245),
    .A2(_01098_),
    .B(net6247),
    .Y(_11824_));
 AOI21x1_ASAP7_75t_R _20047_ (.A1(net5258),
    .A2(net5884),
    .B(net6256),
    .Y(_11825_));
 OAI21x1_ASAP7_75t_R _20048_ (.A1(net5886),
    .A2(_11700_),
    .B(_11825_),
    .Y(_11826_));
 AOI21x1_ASAP7_75t_R _20049_ (.A1(_11824_),
    .A2(_11826_),
    .B(net5875),
    .Y(_11827_));
 AOI21x1_ASAP7_75t_R _20050_ (.A1(_11823_),
    .A2(_11827_),
    .B(net6257),
    .Y(_11828_));
 NAND2x1_ASAP7_75t_R _20051_ (.A(_11818_),
    .B(_11828_),
    .Y(_11829_));
 NAND2x1_ASAP7_75t_R _20052_ (.A(_01097_),
    .B(net6244),
    .Y(_11830_));
 NOR2x1_ASAP7_75t_R _20053_ (.A(_11490_),
    .B(_11519_),
    .Y(_11831_));
 INVx1_ASAP7_75t_R _20054_ (.A(_11831_),
    .Y(_11832_));
 AOI21x1_ASAP7_75t_R _20055_ (.A1(_11830_),
    .A2(_11681_),
    .B(_11832_),
    .Y(_11833_));
 NOR2x1_ASAP7_75t_R _20056_ (.A(net6244),
    .B(_11624_),
    .Y(_11834_));
 OA21x2_ASAP7_75t_R _20057_ (.A1(_11549_),
    .A2(net5009),
    .B(net6244),
    .Y(_11835_));
 OAI21x1_ASAP7_75t_R _20058_ (.A1(_11834_),
    .A2(_11835_),
    .B(_11591_),
    .Y(_11836_));
 NAND2x1_ASAP7_75t_R _20059_ (.A(net6257),
    .B(_11836_),
    .Y(_11837_));
 NOR2x1_ASAP7_75t_R _20060_ (.A(_11833_),
    .B(_11837_),
    .Y(_11838_));
 AND2x2_ASAP7_75t_R _20061_ (.A(_01086_),
    .B(net5302),
    .Y(_11839_));
 NAND2x1_ASAP7_75t_R _20062_ (.A(_11839_),
    .B(net5524),
    .Y(_11840_));
 NAND2x1_ASAP7_75t_R _20063_ (.A(net6244),
    .B(_11840_),
    .Y(_11841_));
 NOR2x1_ASAP7_75t_R _20064_ (.A(net5523),
    .B(_11642_),
    .Y(_11842_));
 NOR2x1_ASAP7_75t_R _20065_ (.A(net4701),
    .B(_11842_),
    .Y(_11843_));
 NAND2x1_ASAP7_75t_R _20066_ (.A(net5879),
    .B(_11746_),
    .Y(_11844_));
 OA21x2_ASAP7_75t_R _20067_ (.A1(net6244),
    .A2(_01102_),
    .B(net5875),
    .Y(_11845_));
 AOI21x1_ASAP7_75t_R _20068_ (.A1(_11845_),
    .A2(_11779_),
    .B(net6248),
    .Y(_11846_));
 OAI21x1_ASAP7_75t_R _20069_ (.A1(_11843_),
    .A2(_11844_),
    .B(_11846_),
    .Y(_11847_));
 AOI21x1_ASAP7_75t_R _20070_ (.A1(_11838_),
    .A2(_11847_),
    .B(_11571_),
    .Y(_11848_));
 NAND2x1_ASAP7_75t_R _20071_ (.A(_11829_),
    .B(_11848_),
    .Y(_11849_));
 OAI21x1_ASAP7_75t_R _20072_ (.A1(_11787_),
    .A2(_11810_),
    .B(_11849_),
    .Y(_00042_));
 NAND2x1_ASAP7_75t_R _20073_ (.A(net4590),
    .B(_11756_),
    .Y(_11850_));
 AO21x1_ASAP7_75t_R _20074_ (.A1(net6258),
    .A2(net5881),
    .B(_11839_),
    .Y(_11851_));
 AO21x1_ASAP7_75t_R _20075_ (.A1(net5199),
    .A2(_11851_),
    .B(net6254),
    .Y(_11852_));
 AO21x1_ASAP7_75t_R _20076_ (.A1(_11850_),
    .A2(_11852_),
    .B(_11832_),
    .Y(_11853_));
 NAND2x1_ASAP7_75t_R _20077_ (.A(net6246),
    .B(_11600_),
    .Y(_11854_));
 NAND2x1_ASAP7_75t_R _20078_ (.A(_11854_),
    .B(_11789_),
    .Y(_11855_));
 AOI21x1_ASAP7_75t_R _20079_ (.A1(_11591_),
    .A2(_11855_),
    .B(net5880),
    .Y(_11856_));
 NAND2x1_ASAP7_75t_R _20080_ (.A(_11853_),
    .B(_11856_),
    .Y(_11857_));
 NAND2x1p5_ASAP7_75t_R _20081_ (.A(net4775),
    .B(net6253),
    .Y(_11858_));
 OA21x2_ASAP7_75t_R _20082_ (.A1(net5875),
    .A2(_11858_),
    .B(_11535_),
    .Y(_11859_));
 NAND2x1_ASAP7_75t_R _20083_ (.A(_11530_),
    .B(net5201),
    .Y(_11860_));
 AO21x1_ASAP7_75t_R _20084_ (.A1(_11860_),
    .A2(_11621_),
    .B(net5879),
    .Y(_11861_));
 AOI21x1_ASAP7_75t_R _20085_ (.A1(_11859_),
    .A2(_11861_),
    .B(net6247),
    .Y(_11862_));
 OAI21x1_ASAP7_75t_R _20086_ (.A1(_11857_),
    .A2(_11862_),
    .B(_11571_),
    .Y(_11863_));
 AOI211x1_ASAP7_75t_R _20087_ (.A1(net5524),
    .A2(_11839_),
    .B(net4953),
    .C(net6254),
    .Y(_11864_));
 AOI21x1_ASAP7_75t_R _20088_ (.A1(_11530_),
    .A2(_11580_),
    .B(_11864_),
    .Y(_11865_));
 AND2x2_ASAP7_75t_R _20089_ (.A(_11797_),
    .B(net5875),
    .Y(_11866_));
 OAI21x1_ASAP7_75t_R _20090_ (.A1(net6249),
    .A2(_11865_),
    .B(_11866_),
    .Y(_11867_));
 NAND2x1_ASAP7_75t_R _20091_ (.A(_11858_),
    .B(_11793_),
    .Y(_11868_));
 INVx1_ASAP7_75t_R _20092_ (.A(_11868_),
    .Y(_11869_));
 OAI21x1_ASAP7_75t_R _20093_ (.A1(net5888),
    .A2(_11699_),
    .B(net6250),
    .Y(_11870_));
 AOI21x1_ASAP7_75t_R _20094_ (.A1(net4948),
    .A2(_11869_),
    .B(_11870_),
    .Y(_11871_));
 NOR2x1_ASAP7_75t_R _20095_ (.A(net6252),
    .B(_11542_),
    .Y(_11872_));
 NOR2x1_ASAP7_75t_R _20096_ (.A(_11872_),
    .B(_11704_),
    .Y(_11873_));
 OAI21x1_ASAP7_75t_R _20097_ (.A1(_11871_),
    .A2(_11873_),
    .B(net5879),
    .Y(_11874_));
 AOI21x1_ASAP7_75t_R _20098_ (.A1(_11867_),
    .A2(_11874_),
    .B(net6257),
    .Y(_11875_));
 NAND2x1_ASAP7_75t_R _20099_ (.A(_11647_),
    .B(_11636_),
    .Y(_11876_));
 OAI21x1_ASAP7_75t_R _20100_ (.A1(net5524),
    .A2(net5891),
    .B(net6245),
    .Y(_11877_));
 NOR2x1_ASAP7_75t_R _20101_ (.A(_11876_),
    .B(_11877_),
    .Y(_11878_));
 AO21x1_ASAP7_75t_R _20102_ (.A1(_11714_),
    .A2(_11722_),
    .B(net6249),
    .Y(_11879_));
 AOI21x1_ASAP7_75t_R _20103_ (.A1(net4951),
    .A2(net4589),
    .B(net6247),
    .Y(_11880_));
 AOI21x1_ASAP7_75t_R _20104_ (.A1(_11880_),
    .A2(_11638_),
    .B(net6257),
    .Y(_11881_));
 OAI21x1_ASAP7_75t_R _20105_ (.A1(_11878_),
    .A2(_11879_),
    .B(_11881_),
    .Y(_11882_));
 OAI21x1_ASAP7_75t_R _20106_ (.A1(_11664_),
    .A2(_11773_),
    .B(net6247),
    .Y(_11883_));
 AOI21x1_ASAP7_75t_R _20107_ (.A1(net4949),
    .A2(_11805_),
    .B(_11883_),
    .Y(_11884_));
 AOI21x1_ASAP7_75t_R _20108_ (.A1(_11624_),
    .A2(net4772),
    .B(net6255),
    .Y(_11885_));
 AOI211x1_ASAP7_75t_R _20109_ (.A1(_11876_),
    .A2(net6255),
    .B(_11885_),
    .C(net6247),
    .Y(_11886_));
 OAI21x1_ASAP7_75t_R _20110_ (.A1(_11884_),
    .A2(_11886_),
    .B(net6257),
    .Y(_11887_));
 AOI21x1_ASAP7_75t_R _20111_ (.A1(_11882_),
    .A2(_11887_),
    .B(net5875),
    .Y(_11888_));
 NOR2x1_ASAP7_75t_R _20112_ (.A(net4953),
    .B(_11773_),
    .Y(_11889_));
 NOR2x1_ASAP7_75t_R _20113_ (.A(_11889_),
    .B(_11712_),
    .Y(_11890_));
 OAI21x1_ASAP7_75t_R _20114_ (.A1(net5882),
    .A2(net5523),
    .B(net6247),
    .Y(_11891_));
 NOR2x1_ASAP7_75t_R _20115_ (.A(_11891_),
    .B(_11703_),
    .Y(_11892_));
 INVx1_ASAP7_75t_R _20116_ (.A(_11737_),
    .Y(_11893_));
 AO21x1_ASAP7_75t_R _20117_ (.A1(_11892_),
    .A2(_11893_),
    .B(net6257),
    .Y(_11894_));
 NOR2x1_ASAP7_75t_R _20118_ (.A(_11890_),
    .B(_11894_),
    .Y(_11895_));
 OAI21x1_ASAP7_75t_R _20119_ (.A1(net4481),
    .A2(net5203),
    .B(net6247),
    .Y(_11896_));
 AOI21x1_ASAP7_75t_R _20120_ (.A1(net5519),
    .A2(_11634_),
    .B(_11896_),
    .Y(_11897_));
 AO21x1_ASAP7_75t_R _20121_ (.A1(net4772),
    .A2(net6244),
    .B(net6247),
    .Y(_11898_));
 NOR2x1_ASAP7_75t_R _20122_ (.A(_11664_),
    .B(_11735_),
    .Y(_11899_));
 OAI21x1_ASAP7_75t_R _20123_ (.A1(_11898_),
    .A2(_11899_),
    .B(net6257),
    .Y(_11900_));
 OAI21x1_ASAP7_75t_R _20124_ (.A1(_11900_),
    .A2(_11897_),
    .B(net5875),
    .Y(_11901_));
 OAI21x1_ASAP7_75t_R _20125_ (.A1(_11901_),
    .A2(_11895_),
    .B(_11572_),
    .Y(_11902_));
 OAI22x1_ASAP7_75t_R _20126_ (.A1(_11863_),
    .A2(_11875_),
    .B1(_11902_),
    .B2(_11888_),
    .Y(_00043_));
 AOI21x1_ASAP7_75t_R _20127_ (.A1(net5303),
    .A2(net5884),
    .B(net6245),
    .Y(_11903_));
 NOR2x1_ASAP7_75t_R _20128_ (.A(net6247),
    .B(_11903_),
    .Y(_11904_));
 AO21x1_ASAP7_75t_R _20129_ (.A1(_11904_),
    .A2(_11707_),
    .B(net5875),
    .Y(_11905_));
 AOI21x1_ASAP7_75t_R _20130_ (.A1(net4770),
    .A2(net4702),
    .B(_11668_),
    .Y(_11906_));
 NOR2x1_ASAP7_75t_R _20131_ (.A(_11905_),
    .B(_11906_),
    .Y(_11907_));
 AO21x1_ASAP7_75t_R _20132_ (.A1(_11678_),
    .A2(net5199),
    .B(net6246),
    .Y(_11908_));
 NOR2x1_ASAP7_75t_R _20133_ (.A(net6249),
    .B(_11739_),
    .Y(_11909_));
 AO21x1_ASAP7_75t_R _20134_ (.A1(_11908_),
    .A2(_11909_),
    .B(net5879),
    .Y(_11910_));
 NOR2x1_ASAP7_75t_R _20135_ (.A(net6247),
    .B(_11834_),
    .Y(_11911_));
 NAND2x1_ASAP7_75t_R _20136_ (.A(net6256),
    .B(net5203),
    .Y(_11912_));
 AND3x1_ASAP7_75t_R _20137_ (.A(_11911_),
    .B(_11765_),
    .C(_11912_),
    .Y(_11913_));
 OAI21x1_ASAP7_75t_R _20138_ (.A1(_11910_),
    .A2(_11913_),
    .B(net5880),
    .Y(_11914_));
 NOR2x1_ASAP7_75t_R _20139_ (.A(_11907_),
    .B(_11914_),
    .Y(_11915_));
 NOR2x1_ASAP7_75t_R _20140_ (.A(net5522),
    .B(_11499_),
    .Y(_11916_));
 AOI21x1_ASAP7_75t_R _20141_ (.A1(_11642_),
    .A2(net5206),
    .B(net6244),
    .Y(_11917_));
 NOR2x1_ASAP7_75t_R _20142_ (.A(_11523_),
    .B(_11519_),
    .Y(_11918_));
 OAI21x1_ASAP7_75t_R _20143_ (.A1(_11916_),
    .A2(_11917_),
    .B(_11918_),
    .Y(_11919_));
 NAND2x1_ASAP7_75t_R _20144_ (.A(net5011),
    .B(net6245),
    .Y(_11920_));
 OA21x2_ASAP7_75t_R _20145_ (.A1(_01092_),
    .A2(net6244),
    .B(_11591_),
    .Y(_11921_));
 AOI21x1_ASAP7_75t_R _20146_ (.A1(net4769),
    .A2(_11921_),
    .B(_11465_),
    .Y(_11922_));
 NAND2x1_ASAP7_75t_R _20147_ (.A(_11919_),
    .B(_11922_),
    .Y(_11923_));
 AOI21x1_ASAP7_75t_R _20148_ (.A1(net5521),
    .A2(_11637_),
    .B(_11604_),
    .Y(_11924_));
 NAND2x1_ASAP7_75t_R _20149_ (.A(net5524),
    .B(net5887),
    .Y(_11925_));
 AOI21x1_ASAP7_75t_R _20150_ (.A1(_11925_),
    .A2(net5206),
    .B(net6244),
    .Y(_11926_));
 NAND2x1_ASAP7_75t_R _20151_ (.A(_11498_),
    .B(net5206),
    .Y(_11927_));
 INVx1_ASAP7_75t_R _20152_ (.A(_11927_),
    .Y(_11928_));
 OAI21x1_ASAP7_75t_R _20153_ (.A1(_11926_),
    .A2(_11928_),
    .B(_11605_),
    .Y(_11929_));
 OAI21x1_ASAP7_75t_R _20154_ (.A1(_11832_),
    .A2(_11924_),
    .B(_11929_),
    .Y(_11930_));
 OAI21x1_ASAP7_75t_R _20155_ (.A1(_11923_),
    .A2(_11930_),
    .B(_11571_),
    .Y(_11931_));
 NOR2x1_ASAP7_75t_R _20156_ (.A(net6247),
    .B(_11467_),
    .Y(_11932_));
 AO21x1_ASAP7_75t_R _20157_ (.A1(_11932_),
    .A2(_11499_),
    .B(net5875),
    .Y(_11933_));
 AOI21x1_ASAP7_75t_R _20158_ (.A1(net5883),
    .A2(net5891),
    .B(net6251),
    .Y(_11934_));
 OAI21x1_ASAP7_75t_R _20159_ (.A1(_11734_),
    .A2(_11735_),
    .B(net6247),
    .Y(_11935_));
 AOI21x1_ASAP7_75t_R _20160_ (.A1(net5202),
    .A2(_11934_),
    .B(_11935_),
    .Y(_11936_));
 OAI21x1_ASAP7_75t_R _20161_ (.A1(_11933_),
    .A2(_11936_),
    .B(net5880),
    .Y(_11937_));
 AOI21x1_ASAP7_75t_R _20162_ (.A1(net5519),
    .A2(_11727_),
    .B(net6244),
    .Y(_11938_));
 AOI21x1_ASAP7_75t_R _20163_ (.A1(_11627_),
    .A2(net5201),
    .B(net6255),
    .Y(_11939_));
 OAI21x1_ASAP7_75t_R _20164_ (.A1(_11938_),
    .A2(_11939_),
    .B(net6249),
    .Y(_11940_));
 NAND2x1_ASAP7_75t_R _20165_ (.A(_11730_),
    .B(_11634_),
    .Y(_11941_));
 NAND2x1_ASAP7_75t_R _20166_ (.A(_11633_),
    .B(_11814_),
    .Y(_11942_));
 AO21x1_ASAP7_75t_R _20167_ (.A1(_11941_),
    .A2(_11942_),
    .B(net6249),
    .Y(_11943_));
 AOI21x1_ASAP7_75t_R _20168_ (.A1(_11940_),
    .A2(_11943_),
    .B(net5879),
    .Y(_11944_));
 NOR2x1_ASAP7_75t_R _20169_ (.A(_11937_),
    .B(_11944_),
    .Y(_11945_));
 NAND2x1_ASAP7_75t_R _20170_ (.A(net5200),
    .B(net4769),
    .Y(_11946_));
 OAI21x1_ASAP7_75t_R _20171_ (.A1(_11686_),
    .A2(_11946_),
    .B(net5879),
    .Y(_11947_));
 NAND2x1_ASAP7_75t_R _20172_ (.A(net6251),
    .B(_11654_),
    .Y(_11948_));
 OAI21x1_ASAP7_75t_R _20173_ (.A1(_11620_),
    .A2(_11948_),
    .B(net6247),
    .Y(_11949_));
 NOR2x1_ASAP7_75t_R _20174_ (.A(_11949_),
    .B(_11502_),
    .Y(_11950_));
 OAI21x1_ASAP7_75t_R _20175_ (.A1(_11947_),
    .A2(_11950_),
    .B(net6257),
    .Y(_11951_));
 NOR2x1_ASAP7_75t_R _20176_ (.A(_11877_),
    .B(_11501_),
    .Y(_11952_));
 AO21x1_ASAP7_75t_R _20177_ (.A1(net4702),
    .A2(net4948),
    .B(net6248),
    .Y(_11953_));
 NOR2x1_ASAP7_75t_R _20178_ (.A(_11952_),
    .B(_11953_),
    .Y(_11954_));
 AOI21x1_ASAP7_75t_R _20179_ (.A1(net5885),
    .A2(net5891),
    .B(net4952),
    .Y(_11955_));
 OAI21x1_ASAP7_75t_R _20180_ (.A1(net6252),
    .A2(_11955_),
    .B(net6248),
    .Y(_11956_));
 OAI21x1_ASAP7_75t_R _20181_ (.A1(_11556_),
    .A2(_11956_),
    .B(net5876),
    .Y(_11957_));
 NOR2x1_ASAP7_75t_R _20182_ (.A(_11954_),
    .B(_11957_),
    .Y(_11958_));
 OAI21x1_ASAP7_75t_R _20183_ (.A1(_11951_),
    .A2(_11958_),
    .B(_11572_),
    .Y(_11959_));
 OAI22x1_ASAP7_75t_R _20184_ (.A1(_11915_),
    .A2(_11931_),
    .B1(_11945_),
    .B2(_11959_),
    .Y(_00044_));
 AO21x1_ASAP7_75t_R _20185_ (.A1(_11658_),
    .A2(_11659_),
    .B(_11667_),
    .Y(_11960_));
 AND2x2_ASAP7_75t_R _20186_ (.A(_11841_),
    .B(net6247),
    .Y(_11961_));
 AO21x1_ASAP7_75t_R _20187_ (.A1(_11598_),
    .A2(_11676_),
    .B(net5875),
    .Y(_11962_));
 AO21x1_ASAP7_75t_R _20188_ (.A1(_11960_),
    .A2(_11961_),
    .B(_11962_),
    .Y(_11963_));
 NAND2x1_ASAP7_75t_R _20189_ (.A(net5301),
    .B(net6246),
    .Y(_11964_));
 NAND2x1_ASAP7_75t_R _20190_ (.A(net6256),
    .B(_11580_),
    .Y(_11965_));
 AOI21x1_ASAP7_75t_R _20191_ (.A1(_11964_),
    .A2(_11965_),
    .B(_11832_),
    .Y(_11966_));
 AOI21x1_ASAP7_75t_R _20192_ (.A1(net4591),
    .A2(_11795_),
    .B(net6246),
    .Y(_11967_));
 NOR2x1_ASAP7_75t_R _20193_ (.A(_11527_),
    .B(_11597_),
    .Y(_11968_));
 OAI21x1_ASAP7_75t_R _20194_ (.A1(_11967_),
    .A2(_11968_),
    .B(_11918_),
    .Y(_11969_));
 NAND2x1_ASAP7_75t_R _20195_ (.A(net6257),
    .B(_11969_),
    .Y(_11970_));
 NOR2x1_ASAP7_75t_R _20196_ (.A(_11966_),
    .B(_11970_),
    .Y(_11971_));
 NAND2x1_ASAP7_75t_R _20197_ (.A(_11963_),
    .B(_11971_),
    .Y(_11972_));
 NOR2x1_ASAP7_75t_R _20198_ (.A(net5524),
    .B(_11700_),
    .Y(_11973_));
 AOI21x1_ASAP7_75t_R _20199_ (.A1(_11788_),
    .A2(net5205),
    .B(net6247),
    .Y(_11974_));
 OAI21x1_ASAP7_75t_R _20200_ (.A1(net4481),
    .A2(_11973_),
    .B(_11974_),
    .Y(_11975_));
 AND2x2_ASAP7_75t_R _20201_ (.A(_11819_),
    .B(net6247),
    .Y(_11976_));
 AOI21x1_ASAP7_75t_R _20202_ (.A1(_11976_),
    .A2(_11635_),
    .B(net5875),
    .Y(_11977_));
 AOI21x1_ASAP7_75t_R _20203_ (.A1(_11975_),
    .A2(_11977_),
    .B(net6257),
    .Y(_11978_));
 OA21x2_ASAP7_75t_R _20204_ (.A1(net4951),
    .A2(net6256),
    .B(net6249),
    .Y(_11979_));
 NOR2x1_ASAP7_75t_R _20205_ (.A(net5299),
    .B(net5524),
    .Y(_11980_));
 OAI21x1_ASAP7_75t_R _20206_ (.A1(_11980_),
    .A2(_11713_),
    .B(net6256),
    .Y(_11981_));
 AOI21x1_ASAP7_75t_R _20207_ (.A1(_11979_),
    .A2(_11981_),
    .B(net5879),
    .Y(_11982_));
 NAND2x1_ASAP7_75t_R _20208_ (.A(net6256),
    .B(net5522),
    .Y(_11983_));
 NAND2x1_ASAP7_75t_R _20209_ (.A(_11983_),
    .B(_11582_),
    .Y(_11984_));
 NAND2x1_ASAP7_75t_R _20210_ (.A(_11982_),
    .B(_11984_),
    .Y(_11985_));
 AOI21x1_ASAP7_75t_R _20211_ (.A1(_11978_),
    .A2(_11985_),
    .B(_11572_),
    .Y(_11986_));
 NAND2x1_ASAP7_75t_R _20212_ (.A(_11972_),
    .B(_11986_),
    .Y(_11987_));
 AO21x1_ASAP7_75t_R _20213_ (.A1(net5877),
    .A2(net6244),
    .B(net6250),
    .Y(_11988_));
 OAI21x1_ASAP7_75t_R _20214_ (.A1(_11988_),
    .A2(_11917_),
    .B(net5879),
    .Y(_11989_));
 NOR2x1_ASAP7_75t_R _20215_ (.A(_11589_),
    .B(_11713_),
    .Y(_11990_));
 INVx1_ASAP7_75t_R _20216_ (.A(_11642_),
    .Y(_11991_));
 OAI21x1_ASAP7_75t_R _20217_ (.A1(_11659_),
    .A2(_11991_),
    .B(net6250),
    .Y(_11992_));
 AOI21x1_ASAP7_75t_R _20218_ (.A1(net6244),
    .A2(_11990_),
    .B(_11992_),
    .Y(_11993_));
 NOR2x1_ASAP7_75t_R _20219_ (.A(_11989_),
    .B(_11993_),
    .Y(_11994_));
 NAND2x1_ASAP7_75t_R _20220_ (.A(_11755_),
    .B(_11903_),
    .Y(_11995_));
 AND2x2_ASAP7_75t_R _20221_ (.A(_11918_),
    .B(_11920_),
    .Y(_11996_));
 NAND2x1_ASAP7_75t_R _20222_ (.A(_11995_),
    .B(_11996_),
    .Y(_11997_));
 NAND2x1_ASAP7_75t_R _20223_ (.A(net6254),
    .B(_11980_),
    .Y(_11998_));
 OAI21x1_ASAP7_75t_R _20224_ (.A1(net4775),
    .A2(net4950),
    .B(net6245),
    .Y(_11999_));
 NAND3x1_ASAP7_75t_R _20225_ (.A(_11998_),
    .B(_11831_),
    .C(_11999_),
    .Y(_12000_));
 NAND3x1_ASAP7_75t_R _20226_ (.A(_11997_),
    .B(net6257),
    .C(_12000_),
    .Y(_12001_));
 NOR2x1_ASAP7_75t_R _20227_ (.A(_11994_),
    .B(_12001_),
    .Y(_12002_));
 AO21x1_ASAP7_75t_R _20228_ (.A1(_11739_),
    .A2(net5519),
    .B(net4702),
    .Y(_12003_));
 AOI21x1_ASAP7_75t_R _20229_ (.A1(net5882),
    .A2(_11739_),
    .B(net6249),
    .Y(_12004_));
 AOI21x1_ASAP7_75t_R _20230_ (.A1(_11868_),
    .A2(_12004_),
    .B(net5879),
    .Y(_12005_));
 OAI21x1_ASAP7_75t_R _20231_ (.A1(net6248),
    .A2(_12003_),
    .B(_12005_),
    .Y(_12006_));
 NAND2x1_ASAP7_75t_R _20232_ (.A(net4948),
    .B(_11728_),
    .Y(_12007_));
 AOI21x1_ASAP7_75t_R _20233_ (.A1(_12007_),
    .A2(_11665_),
    .B(net6249),
    .Y(_12008_));
 AO21x1_ASAP7_75t_R _20234_ (.A1(_11851_),
    .A2(_11803_),
    .B(net6254),
    .Y(_12009_));
 OAI21x1_ASAP7_75t_R _20235_ (.A1(net5886),
    .A2(_11700_),
    .B(_11788_),
    .Y(_12010_));
 AOI21x1_ASAP7_75t_R _20236_ (.A1(_12009_),
    .A2(_12010_),
    .B(net6247),
    .Y(_12011_));
 OAI21x1_ASAP7_75t_R _20237_ (.A1(_12008_),
    .A2(_12011_),
    .B(net5879),
    .Y(_12012_));
 AOI21x1_ASAP7_75t_R _20238_ (.A1(_12006_),
    .A2(_12012_),
    .B(net6257),
    .Y(_12013_));
 OAI21x1_ASAP7_75t_R _20239_ (.A1(_12002_),
    .A2(_12013_),
    .B(_11572_),
    .Y(_12014_));
 NAND2x1_ASAP7_75t_R _20240_ (.A(_11987_),
    .B(_12014_),
    .Y(_00045_));
 NAND2x1_ASAP7_75t_R _20241_ (.A(_11773_),
    .B(_11793_),
    .Y(_12015_));
 AOI21x1_ASAP7_75t_R _20242_ (.A1(_12015_),
    .A2(_12004_),
    .B(net5879),
    .Y(_12016_));
 NOR2x1_ASAP7_75t_R _20243_ (.A(net6248),
    .B(_11934_),
    .Y(_12017_));
 OAI21x1_ASAP7_75t_R _20244_ (.A1(_11679_),
    .A2(_11681_),
    .B(_12017_),
    .Y(_12018_));
 NAND2x1_ASAP7_75t_R _20245_ (.A(_12016_),
    .B(_12018_),
    .Y(_12019_));
 AO21x1_ASAP7_75t_R _20246_ (.A1(net5877),
    .A2(net5882),
    .B(net6251),
    .Y(_12020_));
 AOI21x1_ASAP7_75t_R _20247_ (.A1(_11948_),
    .A2(_12020_),
    .B(_11760_),
    .Y(_12021_));
 AOI21x1_ASAP7_75t_R _20248_ (.A1(_11658_),
    .A2(_11892_),
    .B(net5875),
    .Y(_12022_));
 OAI21x1_ASAP7_75t_R _20249_ (.A1(net6248),
    .A2(_12021_),
    .B(_12022_),
    .Y(_12023_));
 AOI21x1_ASAP7_75t_R _20250_ (.A1(_12019_),
    .A2(_12023_),
    .B(net6257),
    .Y(_12024_));
 AO21x1_ASAP7_75t_R _20251_ (.A1(net4591),
    .A2(_11795_),
    .B(net6254),
    .Y(_12025_));
 OA21x2_ASAP7_75t_R _20252_ (.A1(_11636_),
    .A2(net6245),
    .B(net6250),
    .Y(_12026_));
 NAND2x1_ASAP7_75t_R _20253_ (.A(_12026_),
    .B(_12025_),
    .Y(_12027_));
 AOI21x1_ASAP7_75t_R _20254_ (.A1(_01096_),
    .A2(net6245),
    .B(net6250),
    .Y(_12028_));
 NAND2x1_ASAP7_75t_R _20255_ (.A(_11788_),
    .B(net5206),
    .Y(_12029_));
 AOI21x1_ASAP7_75t_R _20256_ (.A1(_12028_),
    .A2(_12029_),
    .B(net5876),
    .Y(_12030_));
 INVx1_ASAP7_75t_R _20257_ (.A(_11918_),
    .Y(_12031_));
 AOI21x1_ASAP7_75t_R _20258_ (.A1(_11531_),
    .A2(_11927_),
    .B(_12031_),
    .Y(_12032_));
 AOI21x1_ASAP7_75t_R _20259_ (.A1(_12030_),
    .A2(_12027_),
    .B(_12032_),
    .Y(_12033_));
 NAND2x1_ASAP7_75t_R _20260_ (.A(net5876),
    .B(_11784_),
    .Y(_12034_));
 AOI21x1_ASAP7_75t_R _20261_ (.A1(_12033_),
    .A2(_12034_),
    .B(_11465_),
    .Y(_12035_));
 OAI21x1_ASAP7_75t_R _20262_ (.A1(_12024_),
    .A2(_12035_),
    .B(_11571_),
    .Y(_12036_));
 AO21x1_ASAP7_75t_R _20263_ (.A1(net5877),
    .A2(net5524),
    .B(net6253),
    .Y(_12037_));
 AO21x1_ASAP7_75t_R _20264_ (.A1(_11750_),
    .A2(net4591),
    .B(net6245),
    .Y(_12038_));
 OAI21x1_ASAP7_75t_R _20265_ (.A1(_11973_),
    .A2(_12037_),
    .B(_12038_),
    .Y(_12039_));
 NAND2x1_ASAP7_75t_R _20266_ (.A(_11858_),
    .B(_11605_),
    .Y(_12040_));
 AOI21x1_ASAP7_75t_R _20267_ (.A1(_11681_),
    .A2(_11830_),
    .B(_12040_),
    .Y(_12041_));
 AOI21x1_ASAP7_75t_R _20268_ (.A1(_11591_),
    .A2(_12039_),
    .B(_12041_),
    .Y(_12042_));
 AND2x2_ASAP7_75t_R _20269_ (.A(_11722_),
    .B(_11840_),
    .Y(_12043_));
 NAND2x1_ASAP7_75t_R _20270_ (.A(_12004_),
    .B(_11638_),
    .Y(_12044_));
 OR3x1_ASAP7_75t_R _20271_ (.A(_11588_),
    .B(net5879),
    .C(net6245),
    .Y(_12045_));
 NOR2x1_ASAP7_75t_R _20272_ (.A(net6254),
    .B(_11519_),
    .Y(_12046_));
 NAND2x1_ASAP7_75t_R _20273_ (.A(net5891),
    .B(_11925_),
    .Y(_12047_));
 AOI21x1_ASAP7_75t_R _20274_ (.A1(_12046_),
    .A2(_12047_),
    .B(_11831_),
    .Y(_12048_));
 NAND2x1_ASAP7_75t_R _20275_ (.A(_12045_),
    .B(_12048_),
    .Y(_12049_));
 OAI21x1_ASAP7_75t_R _20276_ (.A1(_12043_),
    .A2(_12044_),
    .B(_12049_),
    .Y(_12050_));
 AOI21x1_ASAP7_75t_R _20277_ (.A1(_12042_),
    .A2(_12050_),
    .B(_11465_),
    .Y(_12051_));
 AO21x1_ASAP7_75t_R _20278_ (.A1(net5200),
    .A2(_11750_),
    .B(net6253),
    .Y(_12052_));
 NAND2x1_ASAP7_75t_R _20279_ (.A(_12052_),
    .B(_11911_),
    .Y(_12053_));
 AND2x2_ASAP7_75t_R _20280_ (.A(_01095_),
    .B(_01101_),
    .Y(_12054_));
 OA21x2_ASAP7_75t_R _20281_ (.A1(net6245),
    .A2(_12054_),
    .B(net6248),
    .Y(_12055_));
 OAI21x1_ASAP7_75t_R _20282_ (.A1(_11701_),
    .A2(_11877_),
    .B(_12055_),
    .Y(_12056_));
 NAND3x1_ASAP7_75t_R _20283_ (.A(_12053_),
    .B(_12056_),
    .C(net5879),
    .Y(_12057_));
 NOR2x1_ASAP7_75t_R _20284_ (.A(_11839_),
    .B(net5524),
    .Y(_12058_));
 NOR2x1_ASAP7_75t_R _20285_ (.A(_12058_),
    .B(_11793_),
    .Y(_12059_));
 AOI21x1_ASAP7_75t_R _20286_ (.A1(net6254),
    .A2(net5522),
    .B(net5879),
    .Y(_12060_));
 NAND2x1_ASAP7_75t_R _20287_ (.A(_11558_),
    .B(_12060_),
    .Y(_12061_));
 NOR2x1_ASAP7_75t_R _20288_ (.A(_12059_),
    .B(_12061_),
    .Y(_12062_));
 NAND2x1_ASAP7_75t_R _20289_ (.A(_11654_),
    .B(_11788_),
    .Y(_12063_));
 AOI21x1_ASAP7_75t_R _20290_ (.A1(net5520),
    .A2(_11739_),
    .B(_11534_),
    .Y(_12064_));
 AOI21x1_ASAP7_75t_R _20291_ (.A1(_12063_),
    .A2(_12064_),
    .B(_11832_),
    .Y(_12065_));
 NOR2x1_ASAP7_75t_R _20292_ (.A(_12062_),
    .B(_12065_),
    .Y(_12066_));
 AOI21x1_ASAP7_75t_R _20293_ (.A1(_12057_),
    .A2(_12066_),
    .B(net6257),
    .Y(_12067_));
 OAI21x1_ASAP7_75t_R _20294_ (.A1(_12051_),
    .A2(_12067_),
    .B(_11572_),
    .Y(_12068_));
 NAND2x1_ASAP7_75t_R _20295_ (.A(_12068_),
    .B(_12036_),
    .Y(_00046_));
 AO21x1_ASAP7_75t_R _20296_ (.A1(net6251),
    .A2(net4773),
    .B(net6249),
    .Y(_12069_));
 INVx1_ASAP7_75t_R _20297_ (.A(_11738_),
    .Y(_12070_));
 OAI21x1_ASAP7_75t_R _20298_ (.A1(_12069_),
    .A2(_12070_),
    .B(net5875),
    .Y(_12071_));
 NOR2x1_ASAP7_75t_R _20299_ (.A(_11773_),
    .B(_11842_),
    .Y(_12072_));
 OAI21x1_ASAP7_75t_R _20300_ (.A1(net6251),
    .A2(_11501_),
    .B(net6249),
    .Y(_12073_));
 NOR2x1_ASAP7_75t_R _20301_ (.A(_12072_),
    .B(_12073_),
    .Y(_12074_));
 OAI21x1_ASAP7_75t_R _20302_ (.A1(_12071_),
    .A2(_12074_),
    .B(net6257),
    .Y(_12075_));
 NOR2x1_ASAP7_75t_R _20303_ (.A(net5887),
    .B(net6244),
    .Y(_12076_));
 AOI21x1_ASAP7_75t_R _20304_ (.A1(net5202),
    .A2(_11934_),
    .B(_12076_),
    .Y(_12077_));
 OAI21x1_ASAP7_75t_R _20305_ (.A1(net6248),
    .A2(_12077_),
    .B(net5879),
    .Y(_12078_));
 AO21x1_ASAP7_75t_R _20306_ (.A1(net5877),
    .A2(net5523),
    .B(net6244),
    .Y(_12079_));
 NOR2x1_ASAP7_75t_R _20307_ (.A(_11842_),
    .B(_12079_),
    .Y(_12080_));
 AO21x1_ASAP7_75t_R _20308_ (.A1(_11814_),
    .A2(_11633_),
    .B(net6249),
    .Y(_12081_));
 NOR2x1_ASAP7_75t_R _20309_ (.A(_12080_),
    .B(_12081_),
    .Y(_12082_));
 NOR2x1_ASAP7_75t_R _20310_ (.A(_12078_),
    .B(_12082_),
    .Y(_12083_));
 OAI21x1_ASAP7_75t_R _20311_ (.A1(_12075_),
    .A2(_12083_),
    .B(_11571_),
    .Y(_12084_));
 AO21x1_ASAP7_75t_R _20312_ (.A1(_11701_),
    .A2(net5524),
    .B(_11659_),
    .Y(_12085_));
 NOR2x1_ASAP7_75t_R _20313_ (.A(net4952),
    .B(_11664_),
    .Y(_12086_));
 NOR2x1_ASAP7_75t_R _20314_ (.A(net6253),
    .B(_12086_),
    .Y(_12087_));
 NOR2x1_ASAP7_75t_R _20315_ (.A(_11870_),
    .B(_12087_),
    .Y(_12088_));
 AO21x1_ASAP7_75t_R _20316_ (.A1(_11654_),
    .A2(net6252),
    .B(net6250),
    .Y(_12089_));
 OAI21x1_ASAP7_75t_R _20317_ (.A1(_12089_),
    .A2(_11928_),
    .B(net5879),
    .Y(_12090_));
 AOI21x1_ASAP7_75t_R _20318_ (.A1(_12085_),
    .A2(_12088_),
    .B(_12090_),
    .Y(_12091_));
 OAI21x1_ASAP7_75t_R _20319_ (.A1(net4774),
    .A2(_11659_),
    .B(_11691_),
    .Y(_12092_));
 AOI21x1_ASAP7_75t_R _20320_ (.A1(_11918_),
    .A2(_12092_),
    .B(net6257),
    .Y(_12093_));
 AO21x1_ASAP7_75t_R _20321_ (.A1(_11820_),
    .A2(_12063_),
    .B(_11832_),
    .Y(_12094_));
 NAND2x1_ASAP7_75t_R _20322_ (.A(_12093_),
    .B(_12094_),
    .Y(_12095_));
 NOR2x1_ASAP7_75t_R _20323_ (.A(_12091_),
    .B(_12095_),
    .Y(_12096_));
 INVx1_ASAP7_75t_R _20324_ (.A(_11546_),
    .Y(_12097_));
 AOI211x1_ASAP7_75t_R _20325_ (.A1(net6244),
    .A2(net5203),
    .B(_12097_),
    .C(net4952),
    .Y(_12098_));
 AO21x1_ASAP7_75t_R _20326_ (.A1(net6252),
    .A2(net5204),
    .B(net6248),
    .Y(_12099_));
 NOR2x1_ASAP7_75t_R _20327_ (.A(_11701_),
    .B(_11877_),
    .Y(_12100_));
 OAI21x1_ASAP7_75t_R _20328_ (.A1(_12099_),
    .A2(_12100_),
    .B(net5876),
    .Y(_12101_));
 OAI21x1_ASAP7_75t_R _20329_ (.A1(_12098_),
    .A2(_12101_),
    .B(_11465_),
    .Y(_12102_));
 AOI21x1_ASAP7_75t_R _20330_ (.A1(_11756_),
    .A2(_12086_),
    .B(net5875),
    .Y(_12103_));
 OAI21x1_ASAP7_75t_R _20331_ (.A1(net4481),
    .A2(net4703),
    .B(_12103_),
    .Y(_12104_));
 AO21x1_ASAP7_75t_R _20332_ (.A1(net5877),
    .A2(net6252),
    .B(net6248),
    .Y(_12105_));
 AOI211x1_ASAP7_75t_R _20333_ (.A1(net5883),
    .A2(_12076_),
    .B(_12105_),
    .C(_11864_),
    .Y(_12106_));
 AOI21x1_ASAP7_75t_R _20334_ (.A1(_11740_),
    .A2(_12104_),
    .B(_12106_),
    .Y(_12107_));
 NOR2x1_ASAP7_75t_R _20335_ (.A(_12102_),
    .B(_12107_),
    .Y(_12108_));
 AND2x2_ASAP7_75t_R _20336_ (.A(_12047_),
    .B(net6252),
    .Y(_12109_));
 NAND2x1_ASAP7_75t_R _20337_ (.A(_01092_),
    .B(net6244),
    .Y(_12110_));
 AOI21x1_ASAP7_75t_R _20338_ (.A1(_12110_),
    .A2(_11546_),
    .B(net5876),
    .Y(_12111_));
 OA21x2_ASAP7_75t_R _20339_ (.A1(_11729_),
    .A2(_12109_),
    .B(_12111_),
    .Y(_12112_));
 AO21x1_ASAP7_75t_R _20340_ (.A1(net4772),
    .A2(net5200),
    .B(net6245),
    .Y(_12113_));
 OA21x2_ASAP7_75t_R _20341_ (.A1(_01101_),
    .A2(net6253),
    .B(_12113_),
    .Y(_12114_));
 OAI21x1_ASAP7_75t_R _20342_ (.A1(net4774),
    .A2(net5010),
    .B(net6244),
    .Y(_12115_));
 OAI21x1_ASAP7_75t_R _20343_ (.A1(_11659_),
    .A2(_11660_),
    .B(_12115_),
    .Y(_12116_));
 AOI21x1_ASAP7_75t_R _20344_ (.A1(_11918_),
    .A2(_12116_),
    .B(_11465_),
    .Y(_12117_));
 OAI21x1_ASAP7_75t_R _20345_ (.A1(_11832_),
    .A2(_12114_),
    .B(_12117_),
    .Y(_12118_));
 OAI21x1_ASAP7_75t_R _20346_ (.A1(_12112_),
    .A2(_12118_),
    .B(_11572_),
    .Y(_12119_));
 OAI22x1_ASAP7_75t_R _20347_ (.A1(_12084_),
    .A2(_12096_),
    .B1(_12108_),
    .B2(_12119_),
    .Y(_00047_));
 NOR2x1_ASAP7_75t_R _20348_ (.A(net6657),
    .B(_00450_),
    .Y(_12120_));
 XOR2x2_ASAP7_75t_R _20349_ (.A(net6613),
    .B(_00630_),
    .Y(_12121_));
 XOR2x2_ASAP7_75t_R _20350_ (.A(net6439),
    .B(net6552),
    .Y(_12122_));
 XOR2x2_ASAP7_75t_R _20351_ (.A(_00598_),
    .B(_00591_),
    .Y(_12123_));
 XOR2x2_ASAP7_75t_R _20352_ (.A(net6584),
    .B(net6611),
    .Y(_12124_));
 XOR2x2_ASAP7_75t_R _20353_ (.A(_12124_),
    .B(_12123_),
    .Y(_12125_));
 NAND2x1p5_ASAP7_75t_R _20354_ (.A(_12122_),
    .B(_12125_),
    .Y(_12126_));
 INVx1_ASAP7_75t_R _20355_ (.A(net6552),
    .Y(_12127_));
 XOR2x2_ASAP7_75t_R _20356_ (.A(net6439),
    .B(_12127_),
    .Y(_12128_));
 XNOR2x2_ASAP7_75t_R _20357_ (.A(net6639),
    .B(_00598_),
    .Y(_12129_));
 XOR2x2_ASAP7_75t_R _20358_ (.A(_12129_),
    .B(_12124_),
    .Y(_12130_));
 NAND2x1_ASAP7_75t_R _20359_ (.A(_12128_),
    .B(_12130_),
    .Y(_12131_));
 AOI21x1_ASAP7_75t_R _20360_ (.A1(_12126_),
    .A2(_12131_),
    .B(net6454),
    .Y(_12132_));
 OAI21x1_ASAP7_75t_R _20361_ (.A1(_12120_),
    .A2(_12132_),
    .B(net6483),
    .Y(_12133_));
 AND2x2_ASAP7_75t_R _20362_ (.A(net6454),
    .B(_00450_),
    .Y(_12134_));
 NAND2x1p5_ASAP7_75t_R _20363_ (.A(_12128_),
    .B(_12125_),
    .Y(_12135_));
 NAND2x1_ASAP7_75t_R _20364_ (.A(_12122_),
    .B(_12130_),
    .Y(_12136_));
 AOI21x1_ASAP7_75t_R _20365_ (.A1(_12135_),
    .A2(_12136_),
    .B(net6454),
    .Y(_12137_));
 OAI21x1_ASAP7_75t_R _20366_ (.A1(_12134_),
    .A2(_12137_),
    .B(_08881_),
    .Y(_12138_));
 NAND2x2_ASAP7_75t_R _20367_ (.A(_12138_),
    .B(_12133_),
    .Y(_12139_));
 INVx1_ASAP7_75t_R _20369_ (.A(net6553),
    .Y(_12140_));
 XOR2x2_ASAP7_75t_R _20370_ (.A(net6631),
    .B(net6606),
    .Y(_12141_));
 NAND2x1_ASAP7_75t_R _20371_ (.A(net6434),
    .B(_12141_),
    .Y(_12142_));
 XNOR2x2_ASAP7_75t_R _20372_ (.A(net6631),
    .B(net6606),
    .Y(_12143_));
 NAND2x1_ASAP7_75t_R _20373_ (.A(net6553),
    .B(_12143_),
    .Y(_12144_));
 XOR2x2_ASAP7_75t_R _20374_ (.A(net6585),
    .B(net6612),
    .Y(_12145_));
 INVx2_ASAP7_75t_R _20375_ (.A(_12145_),
    .Y(_12146_));
 AOI21x1_ASAP7_75t_R _20376_ (.A1(_12142_),
    .A2(_12144_),
    .B(_12146_),
    .Y(_12147_));
 NAND2x1_ASAP7_75t_R _20377_ (.A(net6553),
    .B(_12141_),
    .Y(_12148_));
 NAND2x1_ASAP7_75t_R _20378_ (.A(net6434),
    .B(_12143_),
    .Y(_12149_));
 AOI21x1_ASAP7_75t_R _20379_ (.A1(_12148_),
    .A2(_12149_),
    .B(_12145_),
    .Y(_12150_));
 OAI21x1_ASAP7_75t_R _20381_ (.A1(_12147_),
    .A2(_12150_),
    .B(net6657),
    .Y(_12152_));
 OR2x2_ASAP7_75t_R _20383_ (.A(net6657),
    .B(_00451_),
    .Y(_12154_));
 NAND3x1_ASAP7_75t_R _20384_ (.A(net6361),
    .B(_08875_),
    .C(net6432),
    .Y(_12155_));
 AO21x1_ASAP7_75t_R _20385_ (.A1(net6361),
    .A2(net6432),
    .B(_08875_),
    .Y(_12156_));
 NAND2x2_ASAP7_75t_R _20386_ (.A(_12155_),
    .B(_12156_),
    .Y(_01110_));
 NOR2x1_ASAP7_75t_R _20387_ (.A(net6656),
    .B(_00452_),
    .Y(_12157_));
 INVx1_ASAP7_75t_R _20388_ (.A(_12157_),
    .Y(_12158_));
 INVx1_ASAP7_75t_R _20389_ (.A(net6610),
    .Y(_12159_));
 XOR2x2_ASAP7_75t_R _20390_ (.A(_00592_),
    .B(net6611),
    .Y(_12160_));
 NAND2x1_ASAP7_75t_R _20391_ (.A(_12159_),
    .B(net6431),
    .Y(_12161_));
 XNOR2x2_ASAP7_75t_R _20392_ (.A(net6611),
    .B(_00592_),
    .Y(_12162_));
 NAND2x1_ASAP7_75t_R _20393_ (.A(net6610),
    .B(net6429),
    .Y(_12163_));
 XNOR2x2_ASAP7_75t_R _20394_ (.A(_00657_),
    .B(_00689_),
    .Y(_12164_));
 AOI21x1_ASAP7_75t_R _20395_ (.A1(_12161_),
    .A2(_12163_),
    .B(_12164_),
    .Y(_12165_));
 NAND2x1_ASAP7_75t_R _20396_ (.A(net6610),
    .B(net6431),
    .Y(_12166_));
 NAND2x1_ASAP7_75t_R _20397_ (.A(_12159_),
    .B(net6429),
    .Y(_12167_));
 XOR2x2_ASAP7_75t_R _20398_ (.A(_00657_),
    .B(_00689_),
    .Y(_12168_));
 AOI21x1_ASAP7_75t_R _20399_ (.A1(_12166_),
    .A2(_12167_),
    .B(_12168_),
    .Y(_12169_));
 OAI21x1_ASAP7_75t_R _20400_ (.A1(_12165_),
    .A2(_12169_),
    .B(net6657),
    .Y(_12170_));
 AOI21x1_ASAP7_75t_R _20401_ (.A1(_12158_),
    .A2(_12170_),
    .B(net6482),
    .Y(_12171_));
 INVx1_ASAP7_75t_R _20402_ (.A(_12171_),
    .Y(_12172_));
 NAND3x1_ASAP7_75t_R _20403_ (.A(_12170_),
    .B(net6482),
    .C(_12158_),
    .Y(_12173_));
 NAND2x1_ASAP7_75t_R _20404_ (.A(_12172_),
    .B(_12173_),
    .Y(_12174_));
 NAND3x1_ASAP7_75t_R _20407_ (.A(_12152_),
    .B(net6484),
    .C(_12154_),
    .Y(_12176_));
 AO21x1_ASAP7_75t_R _20408_ (.A1(_12152_),
    .A2(_12154_),
    .B(net6484),
    .Y(_12177_));
 NAND2x1p5_ASAP7_75t_R _20409_ (.A(_12176_),
    .B(_12177_),
    .Y(_12178_));
 INVx1_ASAP7_75t_R _20411_ (.A(net6482),
    .Y(_12179_));
 NAND3x1_ASAP7_75t_R _20412_ (.A(_12170_),
    .B(_12179_),
    .C(_12158_),
    .Y(_12180_));
 AO21x1_ASAP7_75t_R _20413_ (.A1(_12170_),
    .A2(_12158_),
    .B(_12179_),
    .Y(_12181_));
 NAND2x1_ASAP7_75t_R _20414_ (.A(_12180_),
    .B(_12181_),
    .Y(_12182_));
 AO21x1_ASAP7_75t_R _20418_ (.A1(net6239),
    .A2(net6240),
    .B(net4991),
    .Y(_12185_));
 INVx1_ASAP7_75t_R _20420_ (.A(_01105_),
    .Y(_12187_));
 AO21x1_ASAP7_75t_R _20421_ (.A1(net6241),
    .A2(net5871),
    .B(_12187_),
    .Y(_12188_));
 XOR2x2_ASAP7_75t_R _20422_ (.A(_00593_),
    .B(net6629),
    .Y(_12189_));
 XNOR2x2_ASAP7_75t_R _20423_ (.A(net6609),
    .B(_12189_),
    .Y(_12190_));
 XNOR2x2_ASAP7_75t_R _20424_ (.A(_00658_),
    .B(_00690_),
    .Y(_12191_));
 XOR2x2_ASAP7_75t_R _20425_ (.A(net6610),
    .B(net6605),
    .Y(_12192_));
 XOR2x2_ASAP7_75t_R _20426_ (.A(_12191_),
    .B(net6428),
    .Y(_12193_));
 NOR2x1_ASAP7_75t_R _20427_ (.A(_12190_),
    .B(_12193_),
    .Y(_12194_));
 XOR2x2_ASAP7_75t_R _20428_ (.A(_12189_),
    .B(net6609),
    .Y(_12195_));
 XOR2x2_ASAP7_75t_R _20429_ (.A(_00658_),
    .B(_00690_),
    .Y(_12196_));
 XOR2x2_ASAP7_75t_R _20430_ (.A(net6428),
    .B(_12196_),
    .Y(_12197_));
 OAI21x1_ASAP7_75t_R _20431_ (.A1(_12195_),
    .A2(_12197_),
    .B(net6657),
    .Y(_12198_));
 NAND2x1_ASAP7_75t_R _20432_ (.A(_00517_),
    .B(net6454),
    .Y(_12199_));
 OAI21x1_ASAP7_75t_R _20433_ (.A1(_12194_),
    .A2(_12198_),
    .B(_12199_),
    .Y(_12200_));
 XOR2x2_ASAP7_75t_R _20434_ (.A(_12200_),
    .B(_08892_),
    .Y(_12201_));
 AO21x1_ASAP7_75t_R _20437_ (.A1(_12185_),
    .A2(_12188_),
    .B(net6238),
    .Y(_12204_));
 AO21x1_ASAP7_75t_R _20438_ (.A1(net6239),
    .A2(net6240),
    .B(_12187_),
    .Y(_12205_));
 INVx1_ASAP7_75t_R _20439_ (.A(_01111_),
    .Y(_12206_));
 AO21x1_ASAP7_75t_R _20440_ (.A1(net6241),
    .A2(net5871),
    .B(_12206_),
    .Y(_12207_));
 XOR2x2_ASAP7_75t_R _20441_ (.A(_12200_),
    .B(net6481),
    .Y(_12208_));
 AO21x1_ASAP7_75t_R _20444_ (.A1(net4700),
    .A2(_12207_),
    .B(net6232),
    .Y(_12211_));
 XNOR2x2_ASAP7_75t_R _20445_ (.A(net6609),
    .B(net6604),
    .Y(_12212_));
 XOR2x2_ASAP7_75t_R _20446_ (.A(_00659_),
    .B(_00691_),
    .Y(_12213_));
 XOR2x2_ASAP7_75t_R _20447_ (.A(_12212_),
    .B(_12213_),
    .Y(_12214_));
 XOR2x2_ASAP7_75t_R _20448_ (.A(net6633),
    .B(net6630),
    .Y(_12215_));
 XOR2x2_ASAP7_75t_R _20449_ (.A(_12215_),
    .B(net6608),
    .Y(_12216_));
 XOR2x2_ASAP7_75t_R _20450_ (.A(_12214_),
    .B(_12216_),
    .Y(_12217_));
 NOR2x1_ASAP7_75t_R _20451_ (.A(net6656),
    .B(_00515_),
    .Y(_12218_));
 AOI21x1_ASAP7_75t_R _20452_ (.A1(net6656),
    .A2(_12217_),
    .B(_12218_),
    .Y(_12219_));
 XOR2x2_ASAP7_75t_R _20453_ (.A(_12219_),
    .B(_00922_),
    .Y(_12220_));
 AO21x1_ASAP7_75t_R _20456_ (.A1(_12204_),
    .A2(_12211_),
    .B(net6228),
    .Y(_12223_));
 NOR2x1_ASAP7_75t_R _20457_ (.A(net5868),
    .B(net5874),
    .Y(_12224_));
 INVx1_ASAP7_75t_R _20458_ (.A(net4991),
    .Y(_12225_));
 AOI21x1_ASAP7_75t_R _20459_ (.A1(net6240),
    .A2(net6239),
    .B(_12225_),
    .Y(_12226_));
 OA21x2_ASAP7_75t_R _20461_ (.A1(net5517),
    .A2(net4587),
    .B(net6236),
    .Y(_12228_));
 AOI21x1_ASAP7_75t_R _20462_ (.A1(net5871),
    .A2(net6241),
    .B(_12225_),
    .Y(_12229_));
 INVx1_ASAP7_75t_R _20463_ (.A(_12229_),
    .Y(_12230_));
 XOR2x2_ASAP7_75t_R _20465_ (.A(_12219_),
    .B(_08895_),
    .Y(_12232_));
 AO21x1_ASAP7_75t_R _20467_ (.A1(_12230_),
    .A2(net6231),
    .B(net6225),
    .Y(_12234_));
 XOR2x2_ASAP7_75t_R _20468_ (.A(_00595_),
    .B(_00627_),
    .Y(_12235_));
 INVx1_ASAP7_75t_R _20469_ (.A(_00692_),
    .Y(_12236_));
 XOR2x2_ASAP7_75t_R _20470_ (.A(_12235_),
    .B(_12236_),
    .Y(_12237_));
 XOR2x2_ASAP7_75t_R _20471_ (.A(_00628_),
    .B(_00660_),
    .Y(_12238_));
 XOR2x2_ASAP7_75t_R _20472_ (.A(_12237_),
    .B(_12238_),
    .Y(_12239_));
 NOR2x1_ASAP7_75t_R _20475_ (.A(net6656),
    .B(_00514_),
    .Y(_12242_));
 AO21x1_ASAP7_75t_R _20476_ (.A1(_12239_),
    .A2(net6656),
    .B(_12242_),
    .Y(_12243_));
 XOR2x2_ASAP7_75t_R _20477_ (.A(_12243_),
    .B(_08898_),
    .Y(_12244_));
 INVx1_ASAP7_75t_R _20478_ (.A(_12244_),
    .Y(_12245_));
 OA21x2_ASAP7_75t_R _20480_ (.A1(_12228_),
    .A2(_12234_),
    .B(net5867),
    .Y(_12247_));
 NAND2x1_ASAP7_75t_R _20481_ (.A(_12223_),
    .B(_12247_),
    .Y(_12248_));
 NAND2x1_ASAP7_75t_R _20483_ (.A(net5873),
    .B(net5874),
    .Y(_12250_));
 NOR2x1_ASAP7_75t_R _20484_ (.A(net5869),
    .B(_12250_),
    .Y(_12251_));
 NOR2x1_ASAP7_75t_R _20485_ (.A(net6231),
    .B(net4587),
    .Y(_12252_));
 INVx1_ASAP7_75t_R _20486_ (.A(_12252_),
    .Y(_12253_));
 AO21x1_ASAP7_75t_R _20488_ (.A1(net6239),
    .A2(net6240),
    .B(_12206_),
    .Y(_12255_));
 NAND2x1_ASAP7_75t_R _20489_ (.A(_12188_),
    .B(_12255_),
    .Y(_12256_));
 AOI21x1_ASAP7_75t_R _20491_ (.A1(net6231),
    .A2(_12256_),
    .B(net6227),
    .Y(_12258_));
 OA21x2_ASAP7_75t_R _20492_ (.A1(_12251_),
    .A2(_12253_),
    .B(_12258_),
    .Y(_12259_));
 NAND2x1_ASAP7_75t_R _20495_ (.A(_12174_),
    .B(net5873),
    .Y(_12262_));
 NAND2x1_ASAP7_75t_R _20496_ (.A(net5870),
    .B(net5874),
    .Y(_12263_));
 NAND2x1_ASAP7_75t_R _20497_ (.A(_12262_),
    .B(net5512),
    .Y(_12264_));
 OAI21x1_ASAP7_75t_R _20498_ (.A1(net6234),
    .A2(net4947),
    .B(net6227),
    .Y(_12265_));
 AOI21x1_ASAP7_75t_R _20499_ (.A1(net6234),
    .A2(net4947),
    .B(_12265_),
    .Y(_12266_));
 OAI21x1_ASAP7_75t_R _20502_ (.A1(_12259_),
    .A2(_12266_),
    .B(net6222),
    .Y(_12269_));
 XNOR2x2_ASAP7_75t_R _20503_ (.A(_00629_),
    .B(_00661_),
    .Y(_12270_));
 XOR2x2_ASAP7_75t_R _20504_ (.A(_12270_),
    .B(_00693_),
    .Y(_12271_));
 XOR2x2_ASAP7_75t_R _20505_ (.A(net6632),
    .B(_00628_),
    .Y(_12272_));
 XOR2x2_ASAP7_75t_R _20506_ (.A(_12271_),
    .B(_12272_),
    .Y(_12273_));
 NOR2x1_ASAP7_75t_R _20507_ (.A(net6656),
    .B(_00513_),
    .Y(_12274_));
 AO21x1_ASAP7_75t_R _20508_ (.A1(_12273_),
    .A2(net6656),
    .B(_12274_),
    .Y(_12275_));
 XOR2x2_ASAP7_75t_R _20509_ (.A(_12275_),
    .B(_00925_),
    .Y(_12276_));
 INVx1_ASAP7_75t_R _20510_ (.A(_12276_),
    .Y(_12277_));
 AOI21x1_ASAP7_75t_R _20512_ (.A1(_12248_),
    .A2(_12269_),
    .B(net5865),
    .Y(_12279_));
 AO21x1_ASAP7_75t_R _20514_ (.A1(net5870),
    .A2(net5518),
    .B(net6231),
    .Y(_12281_));
 NAND2x1_ASAP7_75t_R _20515_ (.A(net6224),
    .B(_12281_),
    .Y(_12282_));
 INVx1_ASAP7_75t_R _20518_ (.A(net5298),
    .Y(_12285_));
 AO21x1_ASAP7_75t_R _20519_ (.A1(net6239),
    .A2(net6240),
    .B(_12285_),
    .Y(_12286_));
 NAND2x1_ASAP7_75t_R _20520_ (.A(net6231),
    .B(_12286_),
    .Y(_12287_));
 NOR2x1_ASAP7_75t_R _20522_ (.A(net5869),
    .B(net5512),
    .Y(_12289_));
 NOR2x1_ASAP7_75t_R _20523_ (.A(net4698),
    .B(_12289_),
    .Y(_12290_));
 NOR2x1_ASAP7_75t_R _20524_ (.A(_12282_),
    .B(_12290_),
    .Y(_12291_));
 NOR2x2_ASAP7_75t_R _20525_ (.A(_12226_),
    .B(net6238),
    .Y(_12292_));
 INVx1_ASAP7_75t_R _20526_ (.A(_01114_),
    .Y(_12293_));
 AO21x1_ASAP7_75t_R _20527_ (.A1(net6241),
    .A2(net5871),
    .B(_12293_),
    .Y(_12294_));
 AO21x1_ASAP7_75t_R _20528_ (.A1(net4945),
    .A2(_12292_),
    .B(net6225),
    .Y(_12295_));
 AO21x1_ASAP7_75t_R _20529_ (.A1(net5870),
    .A2(net5869),
    .B(net6231),
    .Y(_12296_));
 NOR2x1_ASAP7_75t_R _20530_ (.A(_12296_),
    .B(_12289_),
    .Y(_12297_));
 OAI21x1_ASAP7_75t_R _20531_ (.A1(_12295_),
    .A2(_12297_),
    .B(net6223),
    .Y(_12298_));
 OAI21x1_ASAP7_75t_R _20532_ (.A1(_12291_),
    .A2(_12298_),
    .B(net5865),
    .Y(_12299_));
 AO21x1_ASAP7_75t_R _20533_ (.A1(net5874),
    .A2(net5873),
    .B(net5518),
    .Y(_12300_));
 AOI21x1_ASAP7_75t_R _20536_ (.A1(_12262_),
    .A2(_12300_),
    .B(net6235),
    .Y(_12303_));
 AOI21x1_ASAP7_75t_R _20537_ (.A1(net6240),
    .A2(net6239),
    .B(_01107_),
    .Y(_12304_));
 INVx1_ASAP7_75t_R _20538_ (.A(_12304_),
    .Y(_12305_));
 OAI21x1_ASAP7_75t_R _20539_ (.A1(net6231),
    .A2(_12305_),
    .B(net6225),
    .Y(_12306_));
 AO21x1_ASAP7_75t_R _20540_ (.A1(net6235),
    .A2(net5517),
    .B(_12306_),
    .Y(_12307_));
 OAI21x1_ASAP7_75t_R _20541_ (.A1(_12303_),
    .A2(_12307_),
    .B(net5866),
    .Y(_12308_));
 OA21x2_ASAP7_75t_R _20542_ (.A1(_12132_),
    .A2(_12120_),
    .B(net6467),
    .Y(_12309_));
 OA21x2_ASAP7_75t_R _20543_ (.A1(_12137_),
    .A2(_12134_),
    .B(net6483),
    .Y(_12310_));
 OAI21x1_ASAP7_75t_R _20544_ (.A1(_12309_),
    .A2(_12310_),
    .B(net5869),
    .Y(_12311_));
 NAND2x1_ASAP7_75t_R _20545_ (.A(net6234),
    .B(_12311_),
    .Y(_12312_));
 NAND2x1_ASAP7_75t_R _20546_ (.A(net5518),
    .B(net5870),
    .Y(_12313_));
 AOI21x1_ASAP7_75t_R _20547_ (.A1(net5296),
    .A2(net5868),
    .B(net6238),
    .Y(_12314_));
 NAND2x1_ASAP7_75t_R _20548_ (.A(_12313_),
    .B(_12314_),
    .Y(_12315_));
 OA211x2_ASAP7_75t_R _20549_ (.A1(_12289_),
    .A2(_12312_),
    .B(_12315_),
    .C(net6227),
    .Y(_12316_));
 NOR2x1_ASAP7_75t_R _20550_ (.A(_12308_),
    .B(_12316_),
    .Y(_12317_));
 XNOR2x2_ASAP7_75t_R _20551_ (.A(_00597_),
    .B(net6607),
    .Y(_12318_));
 INVx1_ASAP7_75t_R _20552_ (.A(net6549),
    .Y(_12319_));
 XOR2x2_ASAP7_75t_R _20553_ (.A(_12318_),
    .B(net6427),
    .Y(_12320_));
 XNOR2x2_ASAP7_75t_R _20554_ (.A(net6604),
    .B(net6580),
    .Y(_12321_));
 XOR2x2_ASAP7_75t_R _20555_ (.A(_12320_),
    .B(_12321_),
    .Y(_12322_));
 NOR2x1_ASAP7_75t_R _20557_ (.A(net6656),
    .B(_00512_),
    .Y(_12324_));
 AO21x1_ASAP7_75t_R _20558_ (.A1(_12322_),
    .A2(net6656),
    .B(_12324_),
    .Y(_12325_));
 XOR2x2_ASAP7_75t_R _20559_ (.A(_12325_),
    .B(_00926_),
    .Y(_12326_));
 OAI21x1_ASAP7_75t_R _20561_ (.A1(_12299_),
    .A2(_12317_),
    .B(net6220),
    .Y(_12328_));
 AOI21x1_ASAP7_75t_R _20562_ (.A1(net5871),
    .A2(net6241),
    .B(net5298),
    .Y(_12329_));
 AOI21x1_ASAP7_75t_R _20563_ (.A1(net6240),
    .A2(net6239),
    .B(_01112_),
    .Y(_12330_));
 OAI21x1_ASAP7_75t_R _20564_ (.A1(net5195),
    .A2(net4943),
    .B(net6236),
    .Y(_12331_));
 OA21x2_ASAP7_75t_R _20565_ (.A1(net6236),
    .A2(net4586),
    .B(_12331_),
    .Y(_12332_));
 AOI21x1_ASAP7_75t_R _20567_ (.A1(net6229),
    .A2(_12332_),
    .B(net6223),
    .Y(_12334_));
 INVx1_ASAP7_75t_R _20568_ (.A(_12262_),
    .Y(_12335_));
 NAND2x1_ASAP7_75t_R _20569_ (.A(net5870),
    .B(net5869),
    .Y(_12336_));
 NAND2x1_ASAP7_75t_R _20570_ (.A(_12336_),
    .B(_12311_),
    .Y(_12337_));
 NOR2x1_ASAP7_75t_R _20571_ (.A(_12335_),
    .B(_12337_),
    .Y(_12338_));
 INVx1_ASAP7_75t_R _20573_ (.A(_12329_),
    .Y(_12340_));
 NOR2x1_ASAP7_75t_R _20574_ (.A(_12208_),
    .B(_12340_),
    .Y(_12341_));
 NOR2x1_ASAP7_75t_R _20575_ (.A(net6229),
    .B(_12341_),
    .Y(_12342_));
 OAI21x1_ASAP7_75t_R _20576_ (.A1(net6236),
    .A2(_12338_),
    .B(_12342_),
    .Y(_12343_));
 AND2x2_ASAP7_75t_R _20577_ (.A(_12334_),
    .B(_12343_),
    .Y(_12344_));
 AO21x1_ASAP7_75t_R _20578_ (.A1(_12188_),
    .A2(net4697),
    .B(net6231),
    .Y(_12345_));
 OA21x2_ASAP7_75t_R _20579_ (.A1(net5518),
    .A2(net5197),
    .B(net6232),
    .Y(_12346_));
 NOR2x1_ASAP7_75t_R _20580_ (.A(net6224),
    .B(_12346_),
    .Y(_12347_));
 AOI21x1_ASAP7_75t_R _20581_ (.A1(_12345_),
    .A2(_12347_),
    .B(net5866),
    .Y(_12348_));
 AOI21x1_ASAP7_75t_R _20582_ (.A1(net5871),
    .A2(net6241),
    .B(net4991),
    .Y(_12349_));
 INVx2_ASAP7_75t_R _20583_ (.A(_12349_),
    .Y(_12350_));
 AOI21x1_ASAP7_75t_R _20584_ (.A1(net5868),
    .A2(net5874),
    .B(net6232),
    .Y(_12351_));
 AOI21x1_ASAP7_75t_R _20585_ (.A1(net4584),
    .A2(_12351_),
    .B(net6228),
    .Y(_12352_));
 NAND2x1_ASAP7_75t_R _20586_ (.A(net5873),
    .B(net5869),
    .Y(_12353_));
 AO21x1_ASAP7_75t_R _20588_ (.A1(net5509),
    .A2(_12207_),
    .B(net6237),
    .Y(_12355_));
 NAND2x1_ASAP7_75t_R _20589_ (.A(_12352_),
    .B(_12355_),
    .Y(_12356_));
 AO21x1_ASAP7_75t_R _20590_ (.A1(_12348_),
    .A2(_12356_),
    .B(net6221),
    .Y(_12357_));
 NOR2x1_ASAP7_75t_R _20591_ (.A(net5518),
    .B(net5512),
    .Y(_12358_));
 AO21x1_ASAP7_75t_R _20592_ (.A1(net6241),
    .A2(net5871),
    .B(_01111_),
    .Y(_12359_));
 NAND2x1_ASAP7_75t_R _20593_ (.A(net6236),
    .B(_12359_),
    .Y(_12360_));
 NAND2x1_ASAP7_75t_R _20594_ (.A(net6233),
    .B(_12304_),
    .Y(_12361_));
 AND2x2_ASAP7_75t_R _20595_ (.A(_12361_),
    .B(net6229),
    .Y(_12362_));
 OAI21x1_ASAP7_75t_R _20596_ (.A1(_12358_),
    .A2(_12360_),
    .B(_12362_),
    .Y(_12363_));
 INVx1_ASAP7_75t_R _20597_ (.A(_12306_),
    .Y(_12364_));
 AOI21x1_ASAP7_75t_R _20598_ (.A1(net5070),
    .A2(net5518),
    .B(net6238),
    .Y(_12365_));
 OAI21x1_ASAP7_75t_R _20599_ (.A1(net5518),
    .A2(net5512),
    .B(net4940),
    .Y(_12366_));
 AOI21x1_ASAP7_75t_R _20601_ (.A1(_12364_),
    .A2(_12366_),
    .B(net5866),
    .Y(_12368_));
 AOI21x1_ASAP7_75t_R _20602_ (.A1(_12363_),
    .A2(_12368_),
    .B(net5865),
    .Y(_12369_));
 AOI21x1_ASAP7_75t_R _20603_ (.A1(net5868),
    .A2(net5514),
    .B(net5195),
    .Y(_12370_));
 NOR2x1_ASAP7_75t_R _20604_ (.A(net6230),
    .B(_12370_),
    .Y(_12371_));
 AO21x1_ASAP7_75t_R _20605_ (.A1(net6241),
    .A2(net5871),
    .B(_01107_),
    .Y(_12372_));
 OA21x2_ASAP7_75t_R _20607_ (.A1(_12372_),
    .A2(net6233),
    .B(net6226),
    .Y(_12374_));
 AO21x1_ASAP7_75t_R _20608_ (.A1(net5198),
    .A2(net4700),
    .B(net6236),
    .Y(_12375_));
 NAND2x1_ASAP7_75t_R _20609_ (.A(_12374_),
    .B(_12375_),
    .Y(_12376_));
 AO21x1_ASAP7_75t_R _20610_ (.A1(net6236),
    .A2(net4767),
    .B(net6226),
    .Y(_12377_));
 NOR2x1_ASAP7_75t_R _20611_ (.A(_01119_),
    .B(net6236),
    .Y(_12378_));
 OA21x2_ASAP7_75t_R _20612_ (.A1(_12377_),
    .A2(_12378_),
    .B(net5867),
    .Y(_12379_));
 OAI21x1_ASAP7_75t_R _20613_ (.A1(_12371_),
    .A2(_12376_),
    .B(_12379_),
    .Y(_12380_));
 AOI21x1_ASAP7_75t_R _20614_ (.A1(_12369_),
    .A2(_12380_),
    .B(net6220),
    .Y(_12381_));
 OAI21x1_ASAP7_75t_R _20615_ (.A1(_12344_),
    .A2(_12357_),
    .B(_12381_),
    .Y(_12382_));
 OAI21x1_ASAP7_75t_R _20616_ (.A1(_12279_),
    .A2(_12328_),
    .B(_12382_),
    .Y(_00048_));
 AND3x1_ASAP7_75t_R _20618_ (.A(net5867),
    .B(_01121_),
    .C(net6232),
    .Y(_12384_));
 NOR2x1_ASAP7_75t_R _20619_ (.A(net5518),
    .B(_12250_),
    .Y(_12385_));
 NOR2x1_ASAP7_75t_R _20620_ (.A(_12360_),
    .B(_12385_),
    .Y(_12386_));
 OR3x1_ASAP7_75t_R _20621_ (.A(_12384_),
    .B(_12386_),
    .C(net5865),
    .Y(_12387_));
 NOR2x1_ASAP7_75t_R _20622_ (.A(net6223),
    .B(_12292_),
    .Y(_12388_));
 OA21x2_ASAP7_75t_R _20623_ (.A1(_12385_),
    .A2(_12281_),
    .B(_12388_),
    .Y(_12389_));
 AO21x1_ASAP7_75t_R _20624_ (.A1(net5510),
    .A2(_12188_),
    .B(net6231),
    .Y(_12390_));
 INVx4_ASAP7_75t_R _20625_ (.A(_12139_),
    .Y(_01104_));
 NAND2x1_ASAP7_75t_R _20626_ (.A(net5518),
    .B(net5507),
    .Y(_12391_));
 NAND2x1_ASAP7_75t_R _20627_ (.A(_12391_),
    .B(_12346_),
    .Y(_12392_));
 AND3x1_ASAP7_75t_R _20629_ (.A(_12390_),
    .B(_12392_),
    .C(net6223),
    .Y(_12394_));
 OAI21x1_ASAP7_75t_R _20630_ (.A1(_12389_),
    .A2(_12394_),
    .B(net5865),
    .Y(_12395_));
 AOI21x1_ASAP7_75t_R _20632_ (.A1(_12387_),
    .A2(_12395_),
    .B(net6227),
    .Y(_12397_));
 AO21x1_ASAP7_75t_R _20634_ (.A1(net5873),
    .A2(net5869),
    .B(net6231),
    .Y(_12399_));
 NAND2x1_ASAP7_75t_R _20635_ (.A(net5518),
    .B(net5874),
    .Y(_12400_));
 INVx1_ASAP7_75t_R _20636_ (.A(_12400_),
    .Y(_12401_));
 OA21x2_ASAP7_75t_R _20637_ (.A1(_12399_),
    .A2(_12401_),
    .B(_12392_),
    .Y(_12402_));
 NOR2x1_ASAP7_75t_R _20638_ (.A(net5072),
    .B(net5869),
    .Y(_12403_));
 OAI21x1_ASAP7_75t_R _20639_ (.A1(_12403_),
    .A2(_12296_),
    .B(net6223),
    .Y(_12404_));
 AOI21x1_ASAP7_75t_R _20640_ (.A1(net5870),
    .A2(net5874),
    .B(net5868),
    .Y(_12405_));
 INVx1_ASAP7_75t_R _20641_ (.A(_12405_),
    .Y(_12406_));
 AOI21x1_ASAP7_75t_R _20642_ (.A1(_12406_),
    .A2(_12300_),
    .B(net6237),
    .Y(_12407_));
 OAI21x1_ASAP7_75t_R _20643_ (.A1(_12404_),
    .A2(_12407_),
    .B(net6221),
    .Y(_12408_));
 AOI21x1_ASAP7_75t_R _20644_ (.A1(net5866),
    .A2(_12402_),
    .B(_12408_),
    .Y(_12409_));
 AOI21x1_ASAP7_75t_R _20645_ (.A1(net5872),
    .A2(net5874),
    .B(net5868),
    .Y(_12410_));
 OA21x2_ASAP7_75t_R _20646_ (.A1(_12410_),
    .A2(net4587),
    .B(net6231),
    .Y(_12411_));
 AO21x1_ASAP7_75t_R _20647_ (.A1(net6239),
    .A2(net6240),
    .B(net5296),
    .Y(_12412_));
 AO21x1_ASAP7_75t_R _20648_ (.A1(_12412_),
    .A2(_12372_),
    .B(net6233),
    .Y(_12413_));
 NAND2x1_ASAP7_75t_R _20649_ (.A(net5867),
    .B(_12413_),
    .Y(_12414_));
 OAI21x1_ASAP7_75t_R _20650_ (.A1(_12411_),
    .A2(_12414_),
    .B(net5865),
    .Y(_12415_));
 NOR2x1p5_ASAP7_75t_R _20651_ (.A(net6238),
    .B(_12350_),
    .Y(_12416_));
 AOI21x1_ASAP7_75t_R _20652_ (.A1(net6234),
    .A2(net4942),
    .B(net4479),
    .Y(_12417_));
 INVx1_ASAP7_75t_R _20653_ (.A(_12205_),
    .Y(_12418_));
 NAND2x1_ASAP7_75t_R _20654_ (.A(net6231),
    .B(_12418_),
    .Y(_12419_));
 OA21x2_ASAP7_75t_R _20655_ (.A1(net6231),
    .A2(net4697),
    .B(net6223),
    .Y(_12420_));
 AND3x1_ASAP7_75t_R _20656_ (.A(_12417_),
    .B(_12419_),
    .C(_12420_),
    .Y(_12421_));
 OAI21x1_ASAP7_75t_R _20657_ (.A1(_12415_),
    .A2(_12421_),
    .B(net6227),
    .Y(_12422_));
 OAI21x1_ASAP7_75t_R _20658_ (.A1(_12409_),
    .A2(_12422_),
    .B(net6220),
    .Y(_12423_));
 NOR2x1_ASAP7_75t_R _20659_ (.A(net5518),
    .B(net5874),
    .Y(_12424_));
 NAND2x1_ASAP7_75t_R _20660_ (.A(net6233),
    .B(_12294_),
    .Y(_12425_));
 OAI21x1_ASAP7_75t_R _20661_ (.A1(_12424_),
    .A2(_12425_),
    .B(net6227),
    .Y(_12426_));
 AOI21x1_ASAP7_75t_R _20662_ (.A1(net6234),
    .A2(_12337_),
    .B(_12426_),
    .Y(_12427_));
 AO21x1_ASAP7_75t_R _20663_ (.A1(net6239),
    .A2(net6240),
    .B(net5298),
    .Y(_12428_));
 INVx1_ASAP7_75t_R _20664_ (.A(net5194),
    .Y(_12429_));
 AO21x1_ASAP7_75t_R _20665_ (.A1(_12429_),
    .A2(net6234),
    .B(net6227),
    .Y(_12430_));
 OAI21x1_ASAP7_75t_R _20666_ (.A1(_12430_),
    .A2(_12411_),
    .B(net6223),
    .Y(_12431_));
 NOR2x1_ASAP7_75t_R _20667_ (.A(_12427_),
    .B(_12431_),
    .Y(_12432_));
 AND2x2_ASAP7_75t_R _20668_ (.A(_12340_),
    .B(_12292_),
    .Y(_12433_));
 NAND2x1_ASAP7_75t_R _20669_ (.A(net4700),
    .B(net5198),
    .Y(_12434_));
 NOR2x1_ASAP7_75t_R _20670_ (.A(net6233),
    .B(_12434_),
    .Y(_12435_));
 OAI21x1_ASAP7_75t_R _20671_ (.A1(_12433_),
    .A2(_12435_),
    .B(net6228),
    .Y(_12436_));
 NOR2x1_ASAP7_75t_R _20672_ (.A(net6232),
    .B(net4767),
    .Y(_12437_));
 AOI21x1_ASAP7_75t_R _20674_ (.A1(net5510),
    .A2(_12437_),
    .B(net6227),
    .Y(_12439_));
 AO21x1_ASAP7_75t_R _20675_ (.A1(net5516),
    .A2(net5510),
    .B(net6234),
    .Y(_12440_));
 AOI21x1_ASAP7_75t_R _20676_ (.A1(_12439_),
    .A2(_12440_),
    .B(net6223),
    .Y(_12441_));
 AO21x1_ASAP7_75t_R _20677_ (.A1(_12436_),
    .A2(_12441_),
    .B(net6221),
    .Y(_12442_));
 AO21x1_ASAP7_75t_R _20679_ (.A1(net6239),
    .A2(net6240),
    .B(_12293_),
    .Y(_12444_));
 NOR2x1_ASAP7_75t_R _20680_ (.A(net6238),
    .B(_12229_),
    .Y(_12445_));
 AOI21x1_ASAP7_75t_R _20681_ (.A1(net4939),
    .A2(_12445_),
    .B(net6229),
    .Y(_12446_));
 OAI21x1_ASAP7_75t_R _20682_ (.A1(net6230),
    .A2(_12370_),
    .B(_12446_),
    .Y(_12447_));
 AOI21x1_ASAP7_75t_R _20683_ (.A1(net6230),
    .A2(_12400_),
    .B(_12424_),
    .Y(_12448_));
 NOR2x1_ASAP7_75t_R _20684_ (.A(net6226),
    .B(_12341_),
    .Y(_12449_));
 AOI21x1_ASAP7_75t_R _20685_ (.A1(_12448_),
    .A2(_12449_),
    .B(net6223),
    .Y(_12450_));
 AOI21x1_ASAP7_75t_R _20686_ (.A1(_12447_),
    .A2(_12450_),
    .B(net5865),
    .Y(_12451_));
 AND3x1_ASAP7_75t_R _20687_ (.A(net5198),
    .B(net6236),
    .C(net4946),
    .Y(_12452_));
 AO21x1_ASAP7_75t_R _20689_ (.A1(_12292_),
    .A2(net5196),
    .B(net6224),
    .Y(_12454_));
 NOR2x1_ASAP7_75t_R _20690_ (.A(net5869),
    .B(_12201_),
    .Y(_12455_));
 NAND2x1_ASAP7_75t_R _20691_ (.A(_12455_),
    .B(net5512),
    .Y(_12456_));
 NAND2x1_ASAP7_75t_R _20692_ (.A(net5870),
    .B(net5507),
    .Y(_12457_));
 AOI21x1_ASAP7_75t_R _20693_ (.A1(_12351_),
    .A2(_12457_),
    .B(net6228),
    .Y(_12458_));
 AOI21x1_ASAP7_75t_R _20694_ (.A1(_12456_),
    .A2(_12458_),
    .B(net5867),
    .Y(_12459_));
 OAI21x1_ASAP7_75t_R _20695_ (.A1(_12452_),
    .A2(_12454_),
    .B(_12459_),
    .Y(_12460_));
 AOI21x1_ASAP7_75t_R _20696_ (.A1(_12451_),
    .A2(_12460_),
    .B(net6220),
    .Y(_12461_));
 OAI21x1_ASAP7_75t_R _20697_ (.A1(_12432_),
    .A2(_12442_),
    .B(_12461_),
    .Y(_12462_));
 OAI21x1_ASAP7_75t_R _20698_ (.A1(_12397_),
    .A2(_12423_),
    .B(_12462_),
    .Y(_00049_));
 INVx1_ASAP7_75t_R _20699_ (.A(_12326_),
    .Y(_12463_));
 NAND2x1_ASAP7_75t_R _20700_ (.A(net4584),
    .B(_12351_),
    .Y(_12464_));
 AOI21x1_ASAP7_75t_R _20701_ (.A1(net6230),
    .A2(_12370_),
    .B(net6229),
    .Y(_12465_));
 NAND2x1_ASAP7_75t_R _20702_ (.A(_12464_),
    .B(_12465_),
    .Y(_12466_));
 OAI21x1_ASAP7_75t_R _20703_ (.A1(net5870),
    .A2(net5868),
    .B(net5874),
    .Y(_12467_));
 NAND2x1_ASAP7_75t_R _20704_ (.A(net6232),
    .B(_12467_),
    .Y(_12468_));
 AOI21x1_ASAP7_75t_R _20705_ (.A1(net5871),
    .A2(net6241),
    .B(net5296),
    .Y(_12469_));
 INVx1_ASAP7_75t_R _20706_ (.A(_12469_),
    .Y(_12470_));
 AO21x1_ASAP7_75t_R _20707_ (.A1(_12428_),
    .A2(_12470_),
    .B(net6233),
    .Y(_12471_));
 NAND2x1_ASAP7_75t_R _20708_ (.A(_12468_),
    .B(_12471_),
    .Y(_12472_));
 AOI21x1_ASAP7_75t_R _20709_ (.A1(net6228),
    .A2(_12472_),
    .B(net6222),
    .Y(_12473_));
 NAND2x1_ASAP7_75t_R _20710_ (.A(_12466_),
    .B(_12473_),
    .Y(_12474_));
 NOR2x1_ASAP7_75t_R _20711_ (.A(net5518),
    .B(net5870),
    .Y(_12475_));
 INVx1_ASAP7_75t_R _20712_ (.A(_12372_),
    .Y(_12476_));
 OAI21x1_ASAP7_75t_R _20713_ (.A1(net5192),
    .A2(_12476_),
    .B(net6233),
    .Y(_12477_));
 INVx1_ASAP7_75t_R _20714_ (.A(_12185_),
    .Y(_12478_));
 OAI21x1_ASAP7_75t_R _20715_ (.A1(_12478_),
    .A2(net5517),
    .B(net6238),
    .Y(_12479_));
 AOI21x1_ASAP7_75t_R _20716_ (.A1(_12477_),
    .A2(_12479_),
    .B(net6224),
    .Y(_12480_));
 OAI21x1_ASAP7_75t_R _20717_ (.A1(net5507),
    .A2(_12313_),
    .B(net6238),
    .Y(_12481_));
 OAI21x1_ASAP7_75t_R _20718_ (.A1(net5868),
    .A2(net5515),
    .B(_12314_),
    .Y(_12482_));
 AOI21x1_ASAP7_75t_R _20719_ (.A1(_12481_),
    .A2(_12482_),
    .B(net6228),
    .Y(_12483_));
 NOR2x1_ASAP7_75t_R _20720_ (.A(_12480_),
    .B(_12483_),
    .Y(_12484_));
 AOI21x1_ASAP7_75t_R _20721_ (.A1(net6222),
    .A2(_12484_),
    .B(net5865),
    .Y(_12485_));
 OAI21x1_ASAP7_75t_R _20722_ (.A1(net5193),
    .A2(net4943),
    .B(net6236),
    .Y(_12486_));
 OAI21x1_ASAP7_75t_R _20723_ (.A1(net5195),
    .A2(_12475_),
    .B(net6233),
    .Y(_12487_));
 AOI21x1_ASAP7_75t_R _20724_ (.A1(_12486_),
    .A2(_12487_),
    .B(net6226),
    .Y(_12488_));
 AOI21x1_ASAP7_75t_R _20725_ (.A1(net5297),
    .A2(net5518),
    .B(net6236),
    .Y(_12489_));
 NAND2x1_ASAP7_75t_R _20726_ (.A(net5511),
    .B(_12489_),
    .Y(_12490_));
 AOI21x1_ASAP7_75t_R _20727_ (.A1(_12331_),
    .A2(_12490_),
    .B(net6229),
    .Y(_12491_));
 OAI21x1_ASAP7_75t_R _20728_ (.A1(_12488_),
    .A2(_12491_),
    .B(net5867),
    .Y(_12492_));
 OAI21x1_ASAP7_75t_R _20729_ (.A1(net5296),
    .A2(net5868),
    .B(net6238),
    .Y(_12493_));
 OAI21x1_ASAP7_75t_R _20730_ (.A1(net5192),
    .A2(_12493_),
    .B(net6228),
    .Y(_12494_));
 INVx1_ASAP7_75t_R _20731_ (.A(_12330_),
    .Y(_12495_));
 NAND2x1_ASAP7_75t_R _20732_ (.A(net6232),
    .B(_12495_),
    .Y(_12496_));
 NOR2x1_ASAP7_75t_R _20733_ (.A(net5517),
    .B(_12496_),
    .Y(_12497_));
 NOR2x1_ASAP7_75t_R _20734_ (.A(_12494_),
    .B(_12497_),
    .Y(_12498_));
 NAND2x1p5_ASAP7_75t_R _20735_ (.A(net4584),
    .B(_12292_),
    .Y(_12499_));
 NOR2x1_ASAP7_75t_R _20736_ (.A(net5070),
    .B(net5868),
    .Y(_12500_));
 OAI21x1_ASAP7_75t_R _20737_ (.A1(_12500_),
    .A2(net5192),
    .B(net6238),
    .Y(_12501_));
 AOI21x1_ASAP7_75t_R _20738_ (.A1(_12499_),
    .A2(_12501_),
    .B(net6228),
    .Y(_12502_));
 OAI21x1_ASAP7_75t_R _20739_ (.A1(_12498_),
    .A2(_12502_),
    .B(net6222),
    .Y(_12503_));
 AOI21x1_ASAP7_75t_R _20741_ (.A1(_12492_),
    .A2(_12503_),
    .B(net6221),
    .Y(_12505_));
 AOI21x1_ASAP7_75t_R _20742_ (.A1(_12474_),
    .A2(_12485_),
    .B(_12505_),
    .Y(_12506_));
 NAND2x1_ASAP7_75t_R _20743_ (.A(net5868),
    .B(net5874),
    .Y(_12507_));
 AO21x1_ASAP7_75t_R _20744_ (.A1(net5506),
    .A2(_12188_),
    .B(net6232),
    .Y(_12508_));
 AO21x1_ASAP7_75t_R _20745_ (.A1(_12255_),
    .A2(net4584),
    .B(net6238),
    .Y(_12509_));
 AND3x1_ASAP7_75t_R _20746_ (.A(_12508_),
    .B(net6228),
    .C(_12509_),
    .Y(_12510_));
 AOI21x1_ASAP7_75t_R _20747_ (.A1(net5870),
    .A2(net5507),
    .B(net6238),
    .Y(_12511_));
 AND2x2_ASAP7_75t_R _20748_ (.A(net6238),
    .B(_01121_),
    .Y(_12512_));
 AOI21x1_ASAP7_75t_R _20749_ (.A1(net5506),
    .A2(_12511_),
    .B(_12512_),
    .Y(_12513_));
 AO21x1_ASAP7_75t_R _20750_ (.A1(_12513_),
    .A2(net6224),
    .B(net6222),
    .Y(_12514_));
 OR2x2_ASAP7_75t_R _20751_ (.A(_01119_),
    .B(net6232),
    .Y(_12515_));
 OAI21x1_ASAP7_75t_R _20752_ (.A1(net5518),
    .A2(net5513),
    .B(_12445_),
    .Y(_12516_));
 AOI21x1_ASAP7_75t_R _20753_ (.A1(_12515_),
    .A2(_12516_),
    .B(net6228),
    .Y(_12517_));
 NOR2x1_ASAP7_75t_R _20754_ (.A(net5870),
    .B(net6238),
    .Y(_12518_));
 OAI21x1_ASAP7_75t_R _20755_ (.A1(_12455_),
    .A2(_12518_),
    .B(_12391_),
    .Y(_12519_));
 AOI21x1_ASAP7_75t_R _20756_ (.A1(_12464_),
    .A2(_12519_),
    .B(net6224),
    .Y(_12520_));
 OAI21x1_ASAP7_75t_R _20757_ (.A1(_12517_),
    .A2(_12520_),
    .B(net6222),
    .Y(_12521_));
 OAI21x1_ASAP7_75t_R _20758_ (.A1(_12510_),
    .A2(_12514_),
    .B(_12521_),
    .Y(_12522_));
 OA21x2_ASAP7_75t_R _20759_ (.A1(_01123_),
    .A2(net6232),
    .B(net6228),
    .Y(_12523_));
 AOI21x1_ASAP7_75t_R _20760_ (.A1(_12523_),
    .A2(_12468_),
    .B(net6222),
    .Y(_12524_));
 NAND2x1_ASAP7_75t_R _20761_ (.A(_01118_),
    .B(net6232),
    .Y(_12525_));
 NAND3x1_ASAP7_75t_R _20762_ (.A(_12481_),
    .B(net6224),
    .C(_12525_),
    .Y(_12526_));
 AOI21x1_ASAP7_75t_R _20763_ (.A1(_12524_),
    .A2(_12526_),
    .B(net5865),
    .Y(_12527_));
 AND2x2_ASAP7_75t_R _20764_ (.A(_01107_),
    .B(net5297),
    .Y(_12528_));
 NOR2x1_ASAP7_75t_R _20765_ (.A(_12528_),
    .B(net5518),
    .Y(_12529_));
 OA21x2_ASAP7_75t_R _20766_ (.A1(_12410_),
    .A2(_12529_),
    .B(net6233),
    .Y(_12530_));
 OAI21x1_ASAP7_75t_R _20767_ (.A1(_12360_),
    .A2(_12385_),
    .B(net6229),
    .Y(_12531_));
 AO21x1_ASAP7_75t_R _20768_ (.A1(net4768),
    .A2(_12340_),
    .B(net6236),
    .Y(_12532_));
 NOR2x1_ASAP7_75t_R _20769_ (.A(net6233),
    .B(net4700),
    .Y(_12533_));
 NOR2x1_ASAP7_75t_R _20770_ (.A(net6229),
    .B(_12533_),
    .Y(_12534_));
 AOI21x1_ASAP7_75t_R _20771_ (.A1(_12532_),
    .A2(_12534_),
    .B(net5867),
    .Y(_12535_));
 OAI21x1_ASAP7_75t_R _20772_ (.A1(_12530_),
    .A2(_12531_),
    .B(_12535_),
    .Y(_12536_));
 AOI21x1_ASAP7_75t_R _20773_ (.A1(_12527_),
    .A2(_12536_),
    .B(net6220),
    .Y(_12537_));
 OAI21x1_ASAP7_75t_R _20774_ (.A1(net6221),
    .A2(_12522_),
    .B(_12537_),
    .Y(_12538_));
 OAI21x1_ASAP7_75t_R _20775_ (.A1(_12463_),
    .A2(_12506_),
    .B(_12538_),
    .Y(_00050_));
 NOR2x1_ASAP7_75t_R _20777_ (.A(net6222),
    .B(_12445_),
    .Y(_12540_));
 AO21x1_ASAP7_75t_R _20778_ (.A1(net5506),
    .A2(net4941),
    .B(net6232),
    .Y(_12541_));
 NAND2x1_ASAP7_75t_R _20779_ (.A(net6238),
    .B(_12226_),
    .Y(_12542_));
 OAI21x1_ASAP7_75t_R _20780_ (.A1(net4478),
    .A2(net5867),
    .B(net4696),
    .Y(_12543_));
 AOI21x1_ASAP7_75t_R _20781_ (.A1(_12540_),
    .A2(_12541_),
    .B(_12543_),
    .Y(_12544_));
 OAI21x1_ASAP7_75t_R _20782_ (.A1(net6224),
    .A2(_12544_),
    .B(net6221),
    .Y(_12545_));
 OAI21x1_ASAP7_75t_R _20783_ (.A1(net5193),
    .A2(net4695),
    .B(net6233),
    .Y(_12546_));
 NOR2x1_ASAP7_75t_R _20784_ (.A(net4587),
    .B(_12281_),
    .Y(_12547_));
 NOR2x1_ASAP7_75t_R _20785_ (.A(net6223),
    .B(_12547_),
    .Y(_12548_));
 OA21x2_ASAP7_75t_R _20786_ (.A1(net6238),
    .A2(_12495_),
    .B(net6222),
    .Y(_12549_));
 AO21x1_ASAP7_75t_R _20787_ (.A1(_12549_),
    .A2(_12501_),
    .B(net6228),
    .Y(_12550_));
 AOI21x1_ASAP7_75t_R _20788_ (.A1(_12546_),
    .A2(_12548_),
    .B(_12550_),
    .Y(_12551_));
 OAI21x1_ASAP7_75t_R _20789_ (.A1(_12545_),
    .A2(_12551_),
    .B(net6220),
    .Y(_12552_));
 NAND2x1_ASAP7_75t_R _20790_ (.A(_12528_),
    .B(net5868),
    .Y(_12553_));
 NAND2x1_ASAP7_75t_R _20791_ (.A(_12553_),
    .B(net4940),
    .Y(_12554_));
 OA21x2_ASAP7_75t_R _20792_ (.A1(_12385_),
    .A2(_12360_),
    .B(_12554_),
    .Y(_12555_));
 AND2x2_ASAP7_75t_R _20793_ (.A(_12494_),
    .B(net5867),
    .Y(_12556_));
 OAI21x1_ASAP7_75t_R _20794_ (.A1(net6229),
    .A2(_12555_),
    .B(_12556_),
    .Y(_12557_));
 AND2x2_ASAP7_75t_R _20795_ (.A(_12458_),
    .B(_12375_),
    .Y(_12558_));
 NAND2x1_ASAP7_75t_R _20796_ (.A(_12495_),
    .B(net5196),
    .Y(_12559_));
 AOI21x1_ASAP7_75t_R _20797_ (.A1(net4938),
    .A2(net4768),
    .B(net6233),
    .Y(_12560_));
 AOI211x1_ASAP7_75t_R _20798_ (.A1(_12559_),
    .A2(net6233),
    .B(_12560_),
    .C(net6226),
    .Y(_12561_));
 OAI21x1_ASAP7_75t_R _20799_ (.A1(_12558_),
    .A2(_12561_),
    .B(net6223),
    .Y(_12562_));
 AOI21x1_ASAP7_75t_R _20800_ (.A1(_12557_),
    .A2(_12562_),
    .B(net6221),
    .Y(_12563_));
 OA21x2_ASAP7_75t_R _20801_ (.A1(_12500_),
    .A2(net4586),
    .B(net6238),
    .Y(_12564_));
 NOR2x1_ASAP7_75t_R _20802_ (.A(_12564_),
    .B(_12426_),
    .Y(_12565_));
 OAI21x1_ASAP7_75t_R _20803_ (.A1(net5874),
    .A2(net5873),
    .B(net6224),
    .Y(_12566_));
 NOR2x1_ASAP7_75t_R _20804_ (.A(_12335_),
    .B(_12566_),
    .Y(_12567_));
 NAND2x1_ASAP7_75t_R _20805_ (.A(net5869),
    .B(net6231),
    .Y(_12568_));
 AO21x1_ASAP7_75t_R _20806_ (.A1(_12567_),
    .A2(_12568_),
    .B(net6223),
    .Y(_12569_));
 OAI21x1_ASAP7_75t_R _20807_ (.A1(_12565_),
    .A2(_12569_),
    .B(net5865),
    .Y(_12570_));
 NAND2x1_ASAP7_75t_R _20808_ (.A(_12255_),
    .B(_12406_),
    .Y(_12571_));
 AOI21x1_ASAP7_75t_R _20809_ (.A1(_12437_),
    .A2(_12300_),
    .B(net6227),
    .Y(_12572_));
 OAI21x1_ASAP7_75t_R _20810_ (.A1(net6237),
    .A2(_12571_),
    .B(_12572_),
    .Y(_12573_));
 AO21x1_ASAP7_75t_R _20811_ (.A1(_12252_),
    .A2(_12207_),
    .B(net6224),
    .Y(_12574_));
 NOR2x1_ASAP7_75t_R _20812_ (.A(net6235),
    .B(_12264_),
    .Y(_12575_));
 OR2x2_ASAP7_75t_R _20813_ (.A(_12574_),
    .B(_12575_),
    .Y(_12576_));
 AOI21x1_ASAP7_75t_R _20814_ (.A1(_12573_),
    .A2(_12576_),
    .B(net5866),
    .Y(_12577_));
 NOR2x1_ASAP7_75t_R _20815_ (.A(_12570_),
    .B(_12577_),
    .Y(_12578_));
 AND2x2_ASAP7_75t_R _20816_ (.A(_12489_),
    .B(net4939),
    .Y(_12579_));
 NAND2x1_ASAP7_75t_R _20817_ (.A(net6236),
    .B(_12185_),
    .Y(_12580_));
 NOR2x1_ASAP7_75t_R _20818_ (.A(net5517),
    .B(_12580_),
    .Y(_12581_));
 OAI21x1_ASAP7_75t_R _20819_ (.A1(_12579_),
    .A2(_12581_),
    .B(net6225),
    .Y(_12582_));
 AOI21x1_ASAP7_75t_R _20820_ (.A1(_12255_),
    .A2(net5198),
    .B(net6232),
    .Y(_12583_));
 OA21x2_ASAP7_75t_R _20821_ (.A1(_12418_),
    .A2(net4585),
    .B(net6231),
    .Y(_12584_));
 OAI21x1_ASAP7_75t_R _20822_ (.A1(_12583_),
    .A2(_12584_),
    .B(net6229),
    .Y(_12585_));
 AOI21x1_ASAP7_75t_R _20823_ (.A1(_12582_),
    .A2(_12585_),
    .B(net5867),
    .Y(_12586_));
 NOR2x1_ASAP7_75t_R _20824_ (.A(net5517),
    .B(_12296_),
    .Y(_12587_));
 OAI21x1_ASAP7_75t_R _20825_ (.A1(_12234_),
    .A2(_12587_),
    .B(net5866),
    .Y(_12588_));
 INVx1_ASAP7_75t_R _20826_ (.A(net5512),
    .Y(_12589_));
 NOR2x1_ASAP7_75t_R _20827_ (.A(_12589_),
    .B(_12399_),
    .Y(_12590_));
 AO21x1_ASAP7_75t_R _20828_ (.A1(_12292_),
    .A2(_12391_),
    .B(net6227),
    .Y(_12591_));
 NOR2x1_ASAP7_75t_R _20829_ (.A(_12590_),
    .B(_12591_),
    .Y(_12592_));
 OAI21x1_ASAP7_75t_R _20830_ (.A1(_12588_),
    .A2(_12592_),
    .B(net6221),
    .Y(_12593_));
 OAI21x1_ASAP7_75t_R _20831_ (.A1(_12586_),
    .A2(_12593_),
    .B(_12463_),
    .Y(_12594_));
 OAI22x1_ASAP7_75t_R _20832_ (.A1(_12552_),
    .A2(_12563_),
    .B1(_12594_),
    .B2(_12578_),
    .Y(_00051_));
 OAI21x1_ASAP7_75t_R _20833_ (.A1(_12403_),
    .A2(_12296_),
    .B(net6224),
    .Y(_12595_));
 AND3x1_ASAP7_75t_R _20834_ (.A(_12400_),
    .B(net6231),
    .C(net5510),
    .Y(_12596_));
 NAND2x1_ASAP7_75t_R _20835_ (.A(net6227),
    .B(net4697),
    .Y(_12597_));
 OA21x2_ASAP7_75t_R _20836_ (.A1(_12597_),
    .A2(net4940),
    .B(net6223),
    .Y(_12598_));
 OAI21x1_ASAP7_75t_R _20837_ (.A1(_12595_),
    .A2(_12596_),
    .B(_12598_),
    .Y(_12599_));
 NAND2x1_ASAP7_75t_R _20838_ (.A(net5865),
    .B(_12599_),
    .Y(_12600_));
 AO21x1_ASAP7_75t_R _20839_ (.A1(net5506),
    .A2(_12188_),
    .B(_12201_),
    .Y(_12601_));
 INVx1_ASAP7_75t_R _20840_ (.A(net5515),
    .Y(_12602_));
 NOR2x1_ASAP7_75t_R _20841_ (.A(_12602_),
    .B(_12312_),
    .Y(_12603_));
 NOR2x1_ASAP7_75t_R _20842_ (.A(net6224),
    .B(_12603_),
    .Y(_12604_));
 OAI21x1_ASAP7_75t_R _20843_ (.A1(_12401_),
    .A2(_12399_),
    .B(net6224),
    .Y(_12605_));
 INVx1_ASAP7_75t_R _20844_ (.A(_12507_),
    .Y(_12606_));
 INVx1_ASAP7_75t_R _20845_ (.A(_12511_),
    .Y(_12607_));
 NOR2x1_ASAP7_75t_R _20846_ (.A(_12606_),
    .B(_12607_),
    .Y(_12608_));
 OAI21x1_ASAP7_75t_R _20847_ (.A1(_12605_),
    .A2(_12608_),
    .B(net5866),
    .Y(_12609_));
 AOI21x1_ASAP7_75t_R _20848_ (.A1(_12601_),
    .A2(_12604_),
    .B(_12609_),
    .Y(_12610_));
 OAI21x1_ASAP7_75t_R _20849_ (.A1(_12600_),
    .A2(_12610_),
    .B(_12463_),
    .Y(_12611_));
 NOR2x1_ASAP7_75t_R _20850_ (.A(net4943),
    .B(_12416_),
    .Y(_12612_));
 AO21x1_ASAP7_75t_R _20851_ (.A1(_12612_),
    .A2(_12449_),
    .B(net5866),
    .Y(_12613_));
 NAND2x1_ASAP7_75t_R _20852_ (.A(net6236),
    .B(_12444_),
    .Y(_12614_));
 NOR2x1_ASAP7_75t_R _20853_ (.A(net4585),
    .B(_12614_),
    .Y(_12615_));
 NAND2x1_ASAP7_75t_R _20854_ (.A(net6225),
    .B(_12366_),
    .Y(_12616_));
 NOR2x1_ASAP7_75t_R _20855_ (.A(_12615_),
    .B(_12616_),
    .Y(_12617_));
 OAI21x1_ASAP7_75t_R _20856_ (.A1(_12617_),
    .A2(_12613_),
    .B(net6221),
    .Y(_12618_));
 NOR2x1_ASAP7_75t_R _20857_ (.A(net6234),
    .B(_12358_),
    .Y(_12619_));
 NAND2x1_ASAP7_75t_R _20858_ (.A(net6229),
    .B(_12471_),
    .Y(_12620_));
 AOI21x1_ASAP7_75t_R _20859_ (.A1(_12391_),
    .A2(_12619_),
    .B(_12620_),
    .Y(_12621_));
 AOI21x1_ASAP7_75t_R _20860_ (.A1(net6230),
    .A2(_12418_),
    .B(net6227),
    .Y(_12622_));
 OAI21x1_ASAP7_75t_R _20861_ (.A1(net6234),
    .A2(_12400_),
    .B(_12622_),
    .Y(_12623_));
 OAI21x1_ASAP7_75t_R _20862_ (.A1(_12371_),
    .A2(_12623_),
    .B(net5866),
    .Y(_12624_));
 NOR2x1_ASAP7_75t_R _20863_ (.A(_12621_),
    .B(_12624_),
    .Y(_12625_));
 NOR2x1_ASAP7_75t_R _20864_ (.A(_12625_),
    .B(_12618_),
    .Y(_12626_));
 AOI21x1_ASAP7_75t_R _20865_ (.A1(net5071),
    .A2(net5518),
    .B(net6232),
    .Y(_12627_));
 NOR2x1_ASAP7_75t_R _20866_ (.A(net6235),
    .B(_12251_),
    .Y(_12628_));
 OAI21x1_ASAP7_75t_R _20867_ (.A1(_12627_),
    .A2(_12628_),
    .B(net6227),
    .Y(_12629_));
 AOI21x1_ASAP7_75t_R _20868_ (.A1(_12230_),
    .A2(_12428_),
    .B(net6231),
    .Y(_12630_));
 OAI21x1_ASAP7_75t_R _20869_ (.A1(net4435),
    .A2(_12303_),
    .B(net6224),
    .Y(_12631_));
 AOI21x1_ASAP7_75t_R _20870_ (.A1(_12629_),
    .A2(_12631_),
    .B(net5866),
    .Y(_12632_));
 AO21x1_ASAP7_75t_R _20871_ (.A1(net5510),
    .A2(net4938),
    .B(net6231),
    .Y(_12633_));
 NOR2x1_ASAP7_75t_R _20872_ (.A(net6227),
    .B(_12455_),
    .Y(_12634_));
 AO21x1_ASAP7_75t_R _20873_ (.A1(_12633_),
    .A2(_12634_),
    .B(net6223),
    .Y(_12635_));
 AO21x1_ASAP7_75t_R _20874_ (.A1(_12418_),
    .A2(net6236),
    .B(net6226),
    .Y(_12636_));
 NOR2x1_ASAP7_75t_R _20875_ (.A(net5517),
    .B(_12287_),
    .Y(_12637_));
 NOR2x1_ASAP7_75t_R _20876_ (.A(net6230),
    .B(_12391_),
    .Y(_12638_));
 NOR3x1_ASAP7_75t_R _20877_ (.A(_12636_),
    .B(_12637_),
    .C(_12638_),
    .Y(_12639_));
 OAI21x1_ASAP7_75t_R _20878_ (.A1(_12635_),
    .A2(_12639_),
    .B(net5865),
    .Y(_12640_));
 NOR2x1_ASAP7_75t_R _20879_ (.A(_12632_),
    .B(_12640_),
    .Y(_12641_));
 OA21x2_ASAP7_75t_R _20880_ (.A1(_12424_),
    .A2(net5192),
    .B(net6234),
    .Y(_12642_));
 AO21x1_ASAP7_75t_R _20881_ (.A1(net4940),
    .A2(net5511),
    .B(net6225),
    .Y(_12643_));
 NOR2x1_ASAP7_75t_R _20882_ (.A(_12642_),
    .B(_12643_),
    .Y(_12644_));
 INVx1_ASAP7_75t_R _20883_ (.A(_01113_),
    .Y(_12645_));
 AOI21x1_ASAP7_75t_R _20884_ (.A1(_12645_),
    .A2(net6234),
    .B(net4479),
    .Y(_12646_));
 OAI21x1_ASAP7_75t_R _20885_ (.A1(net6227),
    .A2(_12646_),
    .B(net6223),
    .Y(_12647_));
 OAI21x1_ASAP7_75t_R _20886_ (.A1(_12644_),
    .A2(_12647_),
    .B(net6221),
    .Y(_12648_));
 AOI21x1_ASAP7_75t_R _20887_ (.A1(net5516),
    .A2(net5511),
    .B(net6231),
    .Y(_12649_));
 AND2x2_ASAP7_75t_R _20888_ (.A(net4940),
    .B(net5509),
    .Y(_12650_));
 OAI21x1_ASAP7_75t_R _20889_ (.A1(_12649_),
    .A2(_12650_),
    .B(net6227),
    .Y(_12651_));
 INVx1_ASAP7_75t_R _20890_ (.A(_12345_),
    .Y(_12652_));
 OAI21x1_ASAP7_75t_R _20891_ (.A1(_12652_),
    .A2(net4694),
    .B(net6224),
    .Y(_12653_));
 AOI21x1_ASAP7_75t_R _20892_ (.A1(_12651_),
    .A2(_12653_),
    .B(net6223),
    .Y(_12654_));
 OAI21x1_ASAP7_75t_R _20893_ (.A1(_12648_),
    .A2(_12654_),
    .B(net6220),
    .Y(_12655_));
 OAI22x1_ASAP7_75t_R _20894_ (.A1(_12626_),
    .A2(_12611_),
    .B1(_12641_),
    .B2(_12655_),
    .Y(_00052_));
 AND3x1_ASAP7_75t_R _20895_ (.A(net4946),
    .B(net4945),
    .C(net6231),
    .Y(_12656_));
 NOR2x1_ASAP7_75t_R _20896_ (.A(_12656_),
    .B(_12307_),
    .Y(_12657_));
 INVx1_ASAP7_75t_R _20897_ (.A(net5070),
    .Y(_12658_));
 OA21x2_ASAP7_75t_R _20898_ (.A1(net5868),
    .A2(_12658_),
    .B(net6238),
    .Y(_12659_));
 OA21x2_ASAP7_75t_R _20899_ (.A1(net5518),
    .A2(net5512),
    .B(_12659_),
    .Y(_12660_));
 OAI21x1_ASAP7_75t_R _20900_ (.A1(net5297),
    .A2(net6236),
    .B(_12362_),
    .Y(_12661_));
 OAI21x1_ASAP7_75t_R _20901_ (.A1(_12660_),
    .A2(_12661_),
    .B(net6223),
    .Y(_12662_));
 NOR2x1_ASAP7_75t_R _20902_ (.A(_12657_),
    .B(_12662_),
    .Y(_12663_));
 AOI22x1_ASAP7_75t_R _20903_ (.A1(net5512),
    .A2(_12455_),
    .B1(net6236),
    .B2(net4946),
    .Y(_12664_));
 AO21x1_ASAP7_75t_R _20904_ (.A1(_12664_),
    .A2(net6227),
    .B(net6222),
    .Y(_12665_));
 AO21x1_ASAP7_75t_R _20905_ (.A1(_12313_),
    .A2(_12495_),
    .B(net6236),
    .Y(_12666_));
 AND3x1_ASAP7_75t_R _20906_ (.A(net4525),
    .B(net6224),
    .C(_12253_),
    .Y(_12667_));
 OAI21x1_ASAP7_75t_R _20907_ (.A1(_12665_),
    .A2(_12667_),
    .B(net5865),
    .Y(_12668_));
 OAI21x1_ASAP7_75t_R _20908_ (.A1(_12663_),
    .A2(_12668_),
    .B(_12463_),
    .Y(_12669_));
 AO21x1_ASAP7_75t_R _20909_ (.A1(_12627_),
    .A2(net5506),
    .B(net4480),
    .Y(_12670_));
 NAND2x1_ASAP7_75t_R _20910_ (.A(net6227),
    .B(_12670_),
    .Y(_12671_));
 AO221x1_ASAP7_75t_R _20911_ (.A1(net6237),
    .A2(net4938),
    .B1(_12292_),
    .B2(_12188_),
    .C(net6227),
    .Y(_12672_));
 AOI21x1_ASAP7_75t_R _20912_ (.A1(_12671_),
    .A2(_12672_),
    .B(net6222),
    .Y(_12673_));
 AO21x1_ASAP7_75t_R _20913_ (.A1(net5874),
    .A2(net6231),
    .B(net6227),
    .Y(_12674_));
 OAI21x1_ASAP7_75t_R _20914_ (.A1(_12674_),
    .A2(_12603_),
    .B(net6222),
    .Y(_12675_));
 NAND2x1_ASAP7_75t_R _20915_ (.A(net4699),
    .B(_12300_),
    .Y(_12676_));
 INVx1_ASAP7_75t_R _20916_ (.A(_12313_),
    .Y(_12677_));
 OA21x2_ASAP7_75t_R _20917_ (.A1(_12602_),
    .A2(_12677_),
    .B(net6234),
    .Y(_12678_));
 AOI211x1_ASAP7_75t_R _20918_ (.A1(_12676_),
    .A2(net6231),
    .B(_12678_),
    .C(net6224),
    .Y(_12679_));
 OAI21x1_ASAP7_75t_R _20919_ (.A1(_12675_),
    .A2(_12679_),
    .B(net6221),
    .Y(_12680_));
 NOR2x1_ASAP7_75t_R _20920_ (.A(_12680_),
    .B(_12673_),
    .Y(_12681_));
 NOR2x1_ASAP7_75t_R _20921_ (.A(net6228),
    .B(_12518_),
    .Y(_12682_));
 AO21x1_ASAP7_75t_R _20922_ (.A1(net5512),
    .A2(net5198),
    .B(net6232),
    .Y(_12683_));
 AOI21x1_ASAP7_75t_R _20923_ (.A1(_12682_),
    .A2(_12683_),
    .B(net5866),
    .Y(_12684_));
 OAI21x1_ASAP7_75t_R _20924_ (.A1(net5868),
    .A2(net5512),
    .B(_12292_),
    .Y(_12685_));
 AOI21x1_ASAP7_75t_R _20925_ (.A1(net5511),
    .A2(_12659_),
    .B(net6226),
    .Y(_12686_));
 NAND2x1_ASAP7_75t_R _20926_ (.A(_12685_),
    .B(_12686_),
    .Y(_12687_));
 AO21x1_ASAP7_75t_R _20927_ (.A1(_12684_),
    .A2(_12687_),
    .B(net6221),
    .Y(_12688_));
 OAI21x1_ASAP7_75t_R _20928_ (.A1(net6237),
    .A2(_12207_),
    .B(net6227),
    .Y(_12689_));
 NOR2x1_ASAP7_75t_R _20929_ (.A(net5872),
    .B(net6232),
    .Y(_12690_));
 OA21x2_ASAP7_75t_R _20930_ (.A1(_12351_),
    .A2(_12690_),
    .B(net4945),
    .Y(_12691_));
 OAI21x1_ASAP7_75t_R _20931_ (.A1(_12689_),
    .A2(_12691_),
    .B(net5866),
    .Y(_12692_));
 NAND2x1_ASAP7_75t_R _20932_ (.A(net6236),
    .B(_12475_),
    .Y(_12693_));
 INVx1_ASAP7_75t_R _20933_ (.A(_12693_),
    .Y(_12694_));
 NOR2x1_ASAP7_75t_R _20934_ (.A(_12694_),
    .B(_12343_),
    .Y(_12695_));
 NOR2x1_ASAP7_75t_R _20935_ (.A(_12692_),
    .B(_12695_),
    .Y(_12696_));
 AOI21x1_ASAP7_75t_R _20936_ (.A1(net6233),
    .A2(_12553_),
    .B(net6229),
    .Y(_12697_));
 OAI21x1_ASAP7_75t_R _20937_ (.A1(_12385_),
    .A2(_12481_),
    .B(_12697_),
    .Y(_12698_));
 AOI21x1_ASAP7_75t_R _20938_ (.A1(_12425_),
    .A2(_12449_),
    .B(net5867),
    .Y(_12699_));
 AOI21x1_ASAP7_75t_R _20939_ (.A1(_12698_),
    .A2(_12699_),
    .B(net5865),
    .Y(_12700_));
 OA21x2_ASAP7_75t_R _20940_ (.A1(_12206_),
    .A2(net6238),
    .B(net6224),
    .Y(_12701_));
 NOR2x1_ASAP7_75t_R _20941_ (.A(_12690_),
    .B(_12351_),
    .Y(_12702_));
 AOI21x1_ASAP7_75t_R _20942_ (.A1(_12701_),
    .A2(_12702_),
    .B(net6222),
    .Y(_12703_));
 OAI21x1_ASAP7_75t_R _20943_ (.A1(net5193),
    .A2(net4586),
    .B(net6238),
    .Y(_12704_));
 NAND2x1_ASAP7_75t_R _20944_ (.A(net6228),
    .B(_12704_),
    .Y(_12705_));
 AO21x1_ASAP7_75t_R _20945_ (.A1(_12292_),
    .A2(net4941),
    .B(_12705_),
    .Y(_12706_));
 NAND2x1_ASAP7_75t_R _20946_ (.A(_12703_),
    .B(_12706_),
    .Y(_12707_));
 AOI21x1_ASAP7_75t_R _20947_ (.A1(_12700_),
    .A2(_12707_),
    .B(_12463_),
    .Y(_12708_));
 OAI21x1_ASAP7_75t_R _20948_ (.A1(_12688_),
    .A2(_12696_),
    .B(_12708_),
    .Y(_12709_));
 OAI21x1_ASAP7_75t_R _20949_ (.A1(_12669_),
    .A2(_12681_),
    .B(_12709_),
    .Y(_00053_));
 NAND2x1_ASAP7_75t_R _20950_ (.A(net5511),
    .B(net4940),
    .Y(_12710_));
 AOI21x1_ASAP7_75t_R _20951_ (.A1(_12360_),
    .A2(_12710_),
    .B(net6226),
    .Y(_12711_));
 OAI21x1_ASAP7_75t_R _20952_ (.A1(_12711_),
    .A2(_12465_),
    .B(net5867),
    .Y(_12712_));
 AO21x1_ASAP7_75t_R _20953_ (.A1(_01117_),
    .A2(net6233),
    .B(net6229),
    .Y(_12713_));
 AO21x1_ASAP7_75t_R _20954_ (.A1(net5511),
    .A2(_12659_),
    .B(_12713_),
    .Y(_12714_));
 INVx1_ASAP7_75t_R _20955_ (.A(net4586),
    .Y(_12715_));
 AO21x1_ASAP7_75t_R _20956_ (.A1(_12470_),
    .A2(_12715_),
    .B(net6238),
    .Y(_12716_));
 OA21x2_ASAP7_75t_R _20957_ (.A1(net5198),
    .A2(net6233),
    .B(net6229),
    .Y(_12717_));
 AOI21x1_ASAP7_75t_R _20958_ (.A1(_12716_),
    .A2(_12717_),
    .B(net5867),
    .Y(_12718_));
 NAND2x1_ASAP7_75t_R _20959_ (.A(_12714_),
    .B(_12718_),
    .Y(_12719_));
 AOI21x1_ASAP7_75t_R _20960_ (.A1(_12712_),
    .A2(_12719_),
    .B(net5865),
    .Y(_12720_));
 AO21x1_ASAP7_75t_R _20961_ (.A1(_12400_),
    .A2(net6231),
    .B(net6224),
    .Y(_12721_));
 OA21x2_ASAP7_75t_R _20962_ (.A1(_12185_),
    .A2(net6231),
    .B(net6225),
    .Y(_12722_));
 AOI21x1_ASAP7_75t_R _20963_ (.A1(_12722_),
    .A2(_12666_),
    .B(net6223),
    .Y(_12723_));
 OAI21x1_ASAP7_75t_R _20964_ (.A1(_12297_),
    .A2(_12721_),
    .B(_12723_),
    .Y(_12724_));
 AOI21x1_ASAP7_75t_R _20965_ (.A1(_12614_),
    .A2(_12607_),
    .B(net4942),
    .Y(_12725_));
 NAND2x1_ASAP7_75t_R _20966_ (.A(net6238),
    .B(net5507),
    .Y(_12726_));
 AOI21x1_ASAP7_75t_R _20967_ (.A1(_12726_),
    .A2(_12567_),
    .B(net5867),
    .Y(_12727_));
 OAI21x1_ASAP7_75t_R _20968_ (.A1(net6224),
    .A2(_12725_),
    .B(_12727_),
    .Y(_12728_));
 AOI21x1_ASAP7_75t_R _20969_ (.A1(_12724_),
    .A2(_12728_),
    .B(net6221),
    .Y(_12729_));
 OAI21x1_ASAP7_75t_R _20970_ (.A1(_12720_),
    .A2(_12729_),
    .B(net6220),
    .Y(_12730_));
 NOR2x1_ASAP7_75t_R _20971_ (.A(net6236),
    .B(_12476_),
    .Y(_12731_));
 NOR2x1_ASAP7_75t_R _20972_ (.A(net5195),
    .B(net4943),
    .Y(_12732_));
 AOI211x1_ASAP7_75t_R _20973_ (.A1(_12731_),
    .A2(_12732_),
    .B(_12694_),
    .C(net4583),
    .Y(_12733_));
 OAI21x1_ASAP7_75t_R _20974_ (.A1(net4944),
    .A2(_12410_),
    .B(net6233),
    .Y(_12734_));
 NAND2x1_ASAP7_75t_R _20975_ (.A(_12444_),
    .B(_12659_),
    .Y(_12735_));
 AOI21x1_ASAP7_75t_R _20976_ (.A1(_12734_),
    .A2(_12735_),
    .B(net6229),
    .Y(_12736_));
 OA21x2_ASAP7_75t_R _20977_ (.A1(_12733_),
    .A2(_12736_),
    .B(net5867),
    .Y(_12737_));
 OA21x2_ASAP7_75t_R _20978_ (.A1(_12476_),
    .A2(net4943),
    .B(net6233),
    .Y(_12738_));
 OA21x2_ASAP7_75t_R _20979_ (.A1(_12738_),
    .A2(_12636_),
    .B(net6223),
    .Y(_12739_));
 AO21x1_ASAP7_75t_R _20980_ (.A1(net5507),
    .A2(net5518),
    .B(net6236),
    .Y(_12740_));
 AO21x1_ASAP7_75t_R _20981_ (.A1(_01116_),
    .A2(_01122_),
    .B(net6233),
    .Y(_12741_));
 AND2x2_ASAP7_75t_R _20982_ (.A(_12741_),
    .B(net6226),
    .Y(_12742_));
 OAI21x1_ASAP7_75t_R _20983_ (.A1(_12589_),
    .A2(_12740_),
    .B(_12742_),
    .Y(_12743_));
 AO21x1_ASAP7_75t_R _20984_ (.A1(_12739_),
    .A2(_12743_),
    .B(net6221),
    .Y(_12744_));
 OAI21x1_ASAP7_75t_R _20985_ (.A1(_12478_),
    .A2(_12405_),
    .B(net6238),
    .Y(_12745_));
 AOI21x1_ASAP7_75t_R _20986_ (.A1(_12525_),
    .A2(_12745_),
    .B(net6224),
    .Y(_12746_));
 AO21x1_ASAP7_75t_R _20987_ (.A1(_12372_),
    .A2(_12715_),
    .B(net6232),
    .Y(_12747_));
 OAI21x1_ASAP7_75t_R _20988_ (.A1(_12405_),
    .A2(_12606_),
    .B(net6232),
    .Y(_12748_));
 AOI21x1_ASAP7_75t_R _20989_ (.A1(_12747_),
    .A2(_12748_),
    .B(net6228),
    .Y(_12749_));
 OAI21x1_ASAP7_75t_R _20990_ (.A1(_12746_),
    .A2(_12749_),
    .B(net6222),
    .Y(_12750_));
 OA21x2_ASAP7_75t_R _20991_ (.A1(_12207_),
    .A2(net6231),
    .B(net6227),
    .Y(_12751_));
 AO21x1_ASAP7_75t_R _20992_ (.A1(_12353_),
    .A2(net5874),
    .B(net6235),
    .Y(_12752_));
 AOI21x1_ASAP7_75t_R _20993_ (.A1(_12751_),
    .A2(_12752_),
    .B(net6222),
    .Y(_12753_));
 AOI21x1_ASAP7_75t_R _20994_ (.A1(net5869),
    .A2(net5512),
    .B(_12677_),
    .Y(_12754_));
 NOR2x1_ASAP7_75t_R _20995_ (.A(_12306_),
    .B(_12630_),
    .Y(_12755_));
 OAI21x1_ASAP7_75t_R _20996_ (.A1(net6235),
    .A2(_12754_),
    .B(_12755_),
    .Y(_12756_));
 AOI21x1_ASAP7_75t_R _20997_ (.A1(_12753_),
    .A2(_12756_),
    .B(net5865),
    .Y(_12757_));
 AOI21x1_ASAP7_75t_R _20998_ (.A1(_12750_),
    .A2(_12757_),
    .B(net6220),
    .Y(_12758_));
 OAI21x1_ASAP7_75t_R _20999_ (.A1(_12737_),
    .A2(_12744_),
    .B(_12758_),
    .Y(_12759_));
 NAND2x1_ASAP7_75t_R _21000_ (.A(_12730_),
    .B(_12759_),
    .Y(_00054_));
 AND2x2_ASAP7_75t_R _21001_ (.A(_12735_),
    .B(_12519_),
    .Y(_12760_));
 AO21x1_ASAP7_75t_R _21002_ (.A1(_12445_),
    .A2(net4939),
    .B(net6226),
    .Y(_12761_));
 OAI21x1_ASAP7_75t_R _21003_ (.A1(_12547_),
    .A2(_12761_),
    .B(net5867),
    .Y(_12762_));
 AOI21x1_ASAP7_75t_R _21004_ (.A1(net6226),
    .A2(_12760_),
    .B(_12762_),
    .Y(_12763_));
 AO21x1_ASAP7_75t_R _21005_ (.A1(net4939),
    .A2(net6234),
    .B(net6227),
    .Y(_12764_));
 INVx1_ASAP7_75t_R _21006_ (.A(_12710_),
    .Y(_12765_));
 OAI21x1_ASAP7_75t_R _21007_ (.A1(_12764_),
    .A2(_12765_),
    .B(net6223),
    .Y(_12766_));
 OA21x2_ASAP7_75t_R _21008_ (.A1(_12410_),
    .A2(_12418_),
    .B(net6230),
    .Y(_12767_));
 OAI21x1_ASAP7_75t_R _21009_ (.A1(_12281_),
    .A2(_12358_),
    .B(net6227),
    .Y(_12768_));
 NOR2x1_ASAP7_75t_R _21010_ (.A(_12767_),
    .B(_12768_),
    .Y(_12769_));
 OAI21x1_ASAP7_75t_R _21011_ (.A1(_12766_),
    .A2(_12769_),
    .B(net5865),
    .Y(_12770_));
 OAI21x1_ASAP7_75t_R _21012_ (.A1(_12763_),
    .A2(_12770_),
    .B(net6220),
    .Y(_12771_));
 NOR2x1_ASAP7_75t_R _21013_ (.A(_12580_),
    .B(_12251_),
    .Y(_12772_));
 OAI21x1_ASAP7_75t_R _21014_ (.A1(net6234),
    .A2(_12358_),
    .B(net6227),
    .Y(_12773_));
 NOR2x1_ASAP7_75t_R _21015_ (.A(_12772_),
    .B(_12773_),
    .Y(_12774_));
 AO21x1_ASAP7_75t_R _21016_ (.A1(net5874),
    .A2(net5873),
    .B(_12568_),
    .Y(_12775_));
 AND2x2_ASAP7_75t_R _21017_ (.A(_12542_),
    .B(net6224),
    .Y(_12776_));
 AO21x1_ASAP7_75t_R _21018_ (.A1(_12775_),
    .A2(_12776_),
    .B(net6223),
    .Y(_12777_));
 OAI21x1_ASAP7_75t_R _21019_ (.A1(_12774_),
    .A2(_12777_),
    .B(net6221),
    .Y(_12778_));
 NAND2x1_ASAP7_75t_R _21020_ (.A(net5509),
    .B(_12391_),
    .Y(_12779_));
 AO21x1_ASAP7_75t_R _21021_ (.A1(net5870),
    .A2(net6234),
    .B(net6224),
    .Y(_12780_));
 AO21x1_ASAP7_75t_R _21022_ (.A1(_12779_),
    .A2(net6231),
    .B(_12780_),
    .Y(_12781_));
 NOR2x1_ASAP7_75t_R _21023_ (.A(_12312_),
    .B(_12251_),
    .Y(_12782_));
 OAI21x1_ASAP7_75t_R _21024_ (.A1(_12608_),
    .A2(_12782_),
    .B(net6224),
    .Y(_12783_));
 AOI21x1_ASAP7_75t_R _21025_ (.A1(_12781_),
    .A2(_12783_),
    .B(net5866),
    .Y(_12784_));
 NOR2x1_ASAP7_75t_R _21026_ (.A(_12778_),
    .B(_12784_),
    .Y(_12785_));
 OA21x2_ASAP7_75t_R _21027_ (.A1(net5874),
    .A2(net6230),
    .B(net6229),
    .Y(_12786_));
 OA21x2_ASAP7_75t_R _21028_ (.A1(net6230),
    .A2(net5196),
    .B(_12786_),
    .Y(_12787_));
 AOI21x1_ASAP7_75t_R _21029_ (.A1(net4526),
    .A2(_12787_),
    .B(net5867),
    .Y(_12788_));
 OA21x2_ASAP7_75t_R _21030_ (.A1(_12410_),
    .A2(_12418_),
    .B(net6236),
    .Y(_12789_));
 AND3x1_ASAP7_75t_R _21031_ (.A(net4768),
    .B(net4941),
    .C(net6233),
    .Y(_12790_));
 OR3x1_ASAP7_75t_R _21032_ (.A(_12789_),
    .B(net6229),
    .C(_12790_),
    .Y(_12791_));
 OA21x2_ASAP7_75t_R _21033_ (.A1(net5297),
    .A2(net6230),
    .B(net6229),
    .Y(_12792_));
 OA21x2_ASAP7_75t_R _21034_ (.A1(_12740_),
    .A2(_12589_),
    .B(_12792_),
    .Y(_12793_));
 INVx1_ASAP7_75t_R _21035_ (.A(_12374_),
    .Y(_12794_));
 AO21x1_ASAP7_75t_R _21036_ (.A1(net5517),
    .A2(net6230),
    .B(_12418_),
    .Y(_12795_));
 OAI21x1_ASAP7_75t_R _21037_ (.A1(_12794_),
    .A2(_12795_),
    .B(net5866),
    .Y(_12796_));
 OAI21x1_ASAP7_75t_R _21038_ (.A1(_12793_),
    .A2(_12796_),
    .B(net5865),
    .Y(_12797_));
 AOI21x1_ASAP7_75t_R _21039_ (.A1(_12788_),
    .A2(_12791_),
    .B(_12797_),
    .Y(_12798_));
 NOR2x1_ASAP7_75t_R _21040_ (.A(_12424_),
    .B(_12281_),
    .Y(_12799_));
 AO21x1_ASAP7_75t_R _21041_ (.A1(_12445_),
    .A2(net4768),
    .B(net6226),
    .Y(_12800_));
 OA21x2_ASAP7_75t_R _21042_ (.A1(_01122_),
    .A2(net6236),
    .B(net6226),
    .Y(_12801_));
 AO21x1_ASAP7_75t_R _21043_ (.A1(_12495_),
    .A2(_12230_),
    .B(net6231),
    .Y(_12802_));
 AOI21x1_ASAP7_75t_R _21044_ (.A1(_12801_),
    .A2(_12802_),
    .B(net6223),
    .Y(_12803_));
 OA21x2_ASAP7_75t_R _21045_ (.A1(_12799_),
    .A2(_12800_),
    .B(_12803_),
    .Y(_12804_));
 NAND2x1_ASAP7_75t_R _21046_ (.A(_12693_),
    .B(_12786_),
    .Y(_12805_));
 NOR2x1_ASAP7_75t_R _21047_ (.A(_12637_),
    .B(_12805_),
    .Y(_12806_));
 NAND2x1_ASAP7_75t_R _21048_ (.A(_01113_),
    .B(net6230),
    .Y(_12807_));
 AO21x1_ASAP7_75t_R _21049_ (.A1(_12374_),
    .A2(_12807_),
    .B(net5866),
    .Y(_12808_));
 OAI21x1_ASAP7_75t_R _21050_ (.A1(_12806_),
    .A2(_12808_),
    .B(net6221),
    .Y(_12809_));
 OAI21x1_ASAP7_75t_R _21051_ (.A1(_12804_),
    .A2(_12809_),
    .B(_12463_),
    .Y(_12810_));
 OAI22x1_ASAP7_75t_R _21052_ (.A1(_12771_),
    .A2(_12785_),
    .B1(_12798_),
    .B2(_12810_),
    .Y(_00055_));
 NOR2x1_ASAP7_75t_R _21053_ (.A(net6663),
    .B(_00453_),
    .Y(_12811_));
 XOR2x2_ASAP7_75t_R _21054_ (.A(_00631_),
    .B(_00638_),
    .Y(_12812_));
 XOR2x2_ASAP7_75t_R _21055_ (.A(net6546),
    .B(_12812_),
    .Y(_12813_));
 XOR2x2_ASAP7_75t_R _21056_ (.A(_00606_),
    .B(_00599_),
    .Y(_12814_));
 XOR2x2_ASAP7_75t_R _21057_ (.A(_00632_),
    .B(_00664_),
    .Y(_12815_));
 XOR2x2_ASAP7_75t_R _21058_ (.A(_12814_),
    .B(_12815_),
    .Y(_12816_));
 NAND2x1p5_ASAP7_75t_R _21059_ (.A(_12813_),
    .B(_12816_),
    .Y(_12817_));
 INVx1_ASAP7_75t_R _21060_ (.A(net6547),
    .Y(_12818_));
 XOR2x2_ASAP7_75t_R _21061_ (.A(_12812_),
    .B(_12818_),
    .Y(_12819_));
 XNOR2x2_ASAP7_75t_R _21062_ (.A(_00599_),
    .B(_00606_),
    .Y(_12820_));
 XOR2x2_ASAP7_75t_R _21063_ (.A(_12820_),
    .B(_12815_),
    .Y(_12821_));
 NAND2x1_ASAP7_75t_R _21064_ (.A(_12819_),
    .B(_12821_),
    .Y(_12822_));
 AOI21x1_ASAP7_75t_R _21065_ (.A1(_12817_),
    .A2(_12822_),
    .B(net6460),
    .Y(_12823_));
 OAI21x1_ASAP7_75t_R _21066_ (.A1(_12811_),
    .A2(_12823_),
    .B(_00951_),
    .Y(_12824_));
 AND2x2_ASAP7_75t_R _21068_ (.A(net6460),
    .B(_00453_),
    .Y(_12826_));
 NAND2x1_ASAP7_75t_R _21069_ (.A(_12819_),
    .B(_12816_),
    .Y(_12827_));
 NAND2x1_ASAP7_75t_R _21070_ (.A(_12813_),
    .B(_12821_),
    .Y(_12828_));
 AOI21x1_ASAP7_75t_R _21071_ (.A1(_12827_),
    .A2(_12828_),
    .B(net6460),
    .Y(_12829_));
 INVx1_ASAP7_75t_R _21072_ (.A(_00951_),
    .Y(_12830_));
 OAI21x1_ASAP7_75t_R _21073_ (.A1(_12826_),
    .A2(_12829_),
    .B(_12830_),
    .Y(_12831_));
 NAND2x2_ASAP7_75t_R _21074_ (.A(_12831_),
    .B(_12824_),
    .Y(_12832_));
 INVx1_ASAP7_75t_R _21076_ (.A(net6548),
    .Y(_12833_));
 XOR2x2_ASAP7_75t_R _21077_ (.A(net6624),
    .B(net6601),
    .Y(_12834_));
 NAND2x1_ASAP7_75t_R _21078_ (.A(_12833_),
    .B(_12834_),
    .Y(_12835_));
 XNOR2x2_ASAP7_75t_R _21079_ (.A(net6624),
    .B(net6601),
    .Y(_12836_));
 NAND2x1_ASAP7_75t_R _21080_ (.A(net6548),
    .B(_12836_),
    .Y(_12837_));
 XOR2x2_ASAP7_75t_R _21081_ (.A(_00631_),
    .B(net6577),
    .Y(_12838_));
 INVx1_ASAP7_75t_R _21082_ (.A(_12838_),
    .Y(_12839_));
 AOI21x1_ASAP7_75t_R _21083_ (.A1(_12835_),
    .A2(_12837_),
    .B(_12839_),
    .Y(_12840_));
 NAND2x1_ASAP7_75t_R _21084_ (.A(net6548),
    .B(_12834_),
    .Y(_12841_));
 NAND2x1_ASAP7_75t_R _21085_ (.A(_12833_),
    .B(_12836_),
    .Y(_12842_));
 AOI21x1_ASAP7_75t_R _21086_ (.A1(_12841_),
    .A2(_12842_),
    .B(net6423),
    .Y(_12843_));
 OAI21x1_ASAP7_75t_R _21087_ (.A1(_12840_),
    .A2(_12843_),
    .B(net6663),
    .Y(_12844_));
 INVx1_ASAP7_75t_R _21088_ (.A(_00950_),
    .Y(_12845_));
 OR2x2_ASAP7_75t_R _21089_ (.A(net6664),
    .B(_00454_),
    .Y(_12846_));
 NAND3x1_ASAP7_75t_R _21090_ (.A(net6360),
    .B(_12845_),
    .C(net6422),
    .Y(_12847_));
 AO21x1_ASAP7_75t_R _21091_ (.A1(net6360),
    .A2(net6422),
    .B(_12845_),
    .Y(_12848_));
 NAND2x1_ASAP7_75t_R _21092_ (.A(_12847_),
    .B(_12848_),
    .Y(_12849_));
 INVx1_ASAP7_75t_R _21094_ (.A(net6602),
    .Y(_12850_));
 XOR2x2_ASAP7_75t_R _21095_ (.A(_00600_),
    .B(_00632_),
    .Y(_12851_));
 NAND2x1_ASAP7_75t_R _21096_ (.A(_12850_),
    .B(net6421),
    .Y(_12852_));
 XNOR2x2_ASAP7_75t_R _21097_ (.A(_00632_),
    .B(_00600_),
    .Y(_12853_));
 NAND2x1_ASAP7_75t_R _21098_ (.A(net6602),
    .B(net6420),
    .Y(_12854_));
 XNOR2x2_ASAP7_75t_R _21099_ (.A(net6574),
    .B(net6544),
    .Y(_12855_));
 AOI21x1_ASAP7_75t_R _21100_ (.A1(_12852_),
    .A2(_12854_),
    .B(_12855_),
    .Y(_12856_));
 NAND2x1_ASAP7_75t_R _21101_ (.A(net6602),
    .B(net6421),
    .Y(_12857_));
 NAND2x1_ASAP7_75t_R _21102_ (.A(_12850_),
    .B(net6420),
    .Y(_12858_));
 XOR2x2_ASAP7_75t_R _21103_ (.A(net6574),
    .B(net6544),
    .Y(_12859_));
 AOI21x1_ASAP7_75t_R _21104_ (.A1(_12857_),
    .A2(_12858_),
    .B(_12859_),
    .Y(_12860_));
 OAI21x1_ASAP7_75t_R _21105_ (.A1(_12856_),
    .A2(_12860_),
    .B(net6661),
    .Y(_12861_));
 NOR2x1_ASAP7_75t_R _21106_ (.A(net6664),
    .B(_00455_),
    .Y(_12862_));
 INVx1_ASAP7_75t_R _21107_ (.A(_12862_),
    .Y(_12863_));
 NAND3x1_ASAP7_75t_R _21108_ (.A(_12861_),
    .B(_00952_),
    .C(_12863_),
    .Y(_12864_));
 AO21x1_ASAP7_75t_R _21109_ (.A1(_12861_),
    .A2(_12863_),
    .B(_00952_),
    .Y(_12865_));
 NAND2x1_ASAP7_75t_R _21110_ (.A(_12864_),
    .B(_12865_),
    .Y(_12866_));
 NAND3x1_ASAP7_75t_R _21113_ (.A(_12844_),
    .B(_00950_),
    .C(_12846_),
    .Y(_12868_));
 AO21x1_ASAP7_75t_R _21114_ (.A1(_12844_),
    .A2(_12846_),
    .B(_00950_),
    .Y(_12869_));
 NAND2x1_ASAP7_75t_R _21115_ (.A(_12868_),
    .B(_12869_),
    .Y(_12870_));
 INVx1_ASAP7_75t_R _21117_ (.A(_00952_),
    .Y(_12871_));
 NAND3x1_ASAP7_75t_R _21118_ (.A(_12861_),
    .B(_12871_),
    .C(_12863_),
    .Y(_12872_));
 AO21x1_ASAP7_75t_R _21119_ (.A1(_12861_),
    .A2(_12863_),
    .B(_12871_),
    .Y(_12873_));
 NAND2x2_ASAP7_75t_R _21120_ (.A(_12872_),
    .B(_12873_),
    .Y(_12874_));
 AND2x2_ASAP7_75t_R _21125_ (.A(_01128_),
    .B(_01130_),
    .Y(_12878_));
 AO21x1_ASAP7_75t_R _21126_ (.A1(net6217),
    .A2(net6218),
    .B(net4937),
    .Y(_12879_));
 AO21x1_ASAP7_75t_R _21128_ (.A1(net5864),
    .A2(net5859),
    .B(net5860),
    .Y(_12881_));
 XOR2x2_ASAP7_75t_R _21129_ (.A(_00601_),
    .B(net6624),
    .Y(_12882_));
 XNOR2x2_ASAP7_75t_R _21130_ (.A(_00634_),
    .B(_12882_),
    .Y(_12883_));
 XNOR2x2_ASAP7_75t_R _21131_ (.A(net6573),
    .B(_00698_),
    .Y(_12884_));
 XOR2x2_ASAP7_75t_R _21132_ (.A(_00633_),
    .B(net6600),
    .Y(_12885_));
 XOR2x2_ASAP7_75t_R _21133_ (.A(_12884_),
    .B(_12885_),
    .Y(_12886_));
 NOR2x1_ASAP7_75t_R _21134_ (.A(_12883_),
    .B(_12886_),
    .Y(_12887_));
 XOR2x2_ASAP7_75t_R _21135_ (.A(_12882_),
    .B(_00634_),
    .Y(_12888_));
 XOR2x2_ASAP7_75t_R _21136_ (.A(net6573),
    .B(_00698_),
    .Y(_12889_));
 XOR2x2_ASAP7_75t_R _21137_ (.A(_12885_),
    .B(_12889_),
    .Y(_12890_));
 OAI21x1_ASAP7_75t_R _21138_ (.A1(_12888_),
    .A2(_12890_),
    .B(net6662),
    .Y(_12891_));
 NAND2x1_ASAP7_75t_R _21139_ (.A(_00539_),
    .B(net6460),
    .Y(_12892_));
 OAI21x1_ASAP7_75t_R _21140_ (.A1(_12887_),
    .A2(_12891_),
    .B(_12892_),
    .Y(_12893_));
 XOR2x2_ASAP7_75t_R _21141_ (.A(_12893_),
    .B(_00953_),
    .Y(_12894_));
 AOI21x1_ASAP7_75t_R _21144_ (.A1(_12879_),
    .A2(_12881_),
    .B(net6209),
    .Y(_12897_));
 INVx1_ASAP7_75t_R _21150_ (.A(_01126_),
    .Y(_12903_));
 AOI21x1_ASAP7_75t_R _21151_ (.A1(net6216),
    .A2(net6215),
    .B(_12903_),
    .Y(_12904_));
 INVx1_ASAP7_75t_R _21152_ (.A(_12904_),
    .Y(_12905_));
 OAI21x1_ASAP7_75t_R _21153_ (.A1(net5859),
    .A2(net5857),
    .B(net4524),
    .Y(_12906_));
 XNOR2x2_ASAP7_75t_R _21154_ (.A(_00667_),
    .B(_00699_),
    .Y(_12907_));
 XOR2x2_ASAP7_75t_R _21155_ (.A(_00634_),
    .B(net6600),
    .Y(_12908_));
 XOR2x2_ASAP7_75t_R _21156_ (.A(_12907_),
    .B(_12908_),
    .Y(_12909_));
 XOR2x2_ASAP7_75t_R _21157_ (.A(_00602_),
    .B(net6624),
    .Y(_12910_));
 XOR2x2_ASAP7_75t_R _21158_ (.A(_12910_),
    .B(_00635_),
    .Y(_12911_));
 XOR2x2_ASAP7_75t_R _21159_ (.A(_12909_),
    .B(_12911_),
    .Y(_12912_));
 NOR2x1_ASAP7_75t_R _21160_ (.A(net6663),
    .B(_00538_),
    .Y(_12913_));
 AOI21x1_ASAP7_75t_R _21161_ (.A1(net6663),
    .A2(_12912_),
    .B(_12913_),
    .Y(_12914_));
 XNOR2x2_ASAP7_75t_R _21162_ (.A(_00954_),
    .B(_12914_),
    .Y(_12915_));
 INVx2_ASAP7_75t_R _21163_ (.A(_12915_),
    .Y(_12916_));
 AOI21x1_ASAP7_75t_R _21166_ (.A1(net6208),
    .A2(_12906_),
    .B(net5856),
    .Y(_12919_));
 INVx1_ASAP7_75t_R _21167_ (.A(_12919_),
    .Y(_12920_));
 XNOR2x2_ASAP7_75t_R _21168_ (.A(_00953_),
    .B(_12893_),
    .Y(_12921_));
 OR2x2_ASAP7_75t_R _21170_ (.A(_01140_),
    .B(net6206),
    .Y(_12923_));
 AOI21x1_ASAP7_75t_R _21171_ (.A1(net6218),
    .A2(net6217),
    .B(net4989),
    .Y(_12924_));
 INVx2_ASAP7_75t_R _21172_ (.A(_12924_),
    .Y(_12925_));
 OA21x2_ASAP7_75t_R _21174_ (.A1(_12925_),
    .A2(net6211),
    .B(net5853),
    .Y(_12927_));
 XOR2x2_ASAP7_75t_R _21175_ (.A(_00604_),
    .B(_00636_),
    .Y(_12928_));
 XOR2x2_ASAP7_75t_R _21176_ (.A(_00637_),
    .B(_00669_),
    .Y(_12929_));
 XOR2x2_ASAP7_75t_R _21177_ (.A(_12929_),
    .B(_00701_),
    .Y(_12930_));
 XNOR2x2_ASAP7_75t_R _21178_ (.A(_12928_),
    .B(_12930_),
    .Y(_12931_));
 NOR2x1_ASAP7_75t_R _21179_ (.A(net6658),
    .B(_00536_),
    .Y(_12932_));
 AO21x1_ASAP7_75t_R _21180_ (.A1(_12931_),
    .A2(net6658),
    .B(_12932_),
    .Y(_12933_));
 XOR2x2_ASAP7_75t_R _21181_ (.A(_12933_),
    .B(_00957_),
    .Y(_12934_));
 INVx1_ASAP7_75t_R _21182_ (.A(_12934_),
    .Y(_12935_));
 AOI21x1_ASAP7_75t_R _21183_ (.A1(_12923_),
    .A2(_12927_),
    .B(_12935_),
    .Y(_12936_));
 OAI21x1_ASAP7_75t_R _21184_ (.A1(_12897_),
    .A2(_12920_),
    .B(_12936_),
    .Y(_12937_));
 AO21x1_ASAP7_75t_R _21185_ (.A1(net6217),
    .A2(net6218),
    .B(net5295),
    .Y(_12938_));
 INVx1_ASAP7_75t_R _21186_ (.A(_12938_),
    .Y(_12939_));
 AO21x1_ASAP7_75t_R _21189_ (.A1(_12939_),
    .A2(net6201),
    .B(net5856),
    .Y(_12942_));
 NAND2x1_ASAP7_75t_R _21190_ (.A(net5863),
    .B(net5862),
    .Y(_12943_));
 AO21x1_ASAP7_75t_R _21191_ (.A1(net5864),
    .A2(net5863),
    .B(net5862),
    .Y(_12944_));
 AOI21x1_ASAP7_75t_R _21192_ (.A1(_12943_),
    .A2(_12944_),
    .B(net6205),
    .Y(_12945_));
 INVx1_ASAP7_75t_R _21194_ (.A(net4990),
    .Y(_12947_));
 AO21x1_ASAP7_75t_R _21195_ (.A1(net6215),
    .A2(net6216),
    .B(_12947_),
    .Y(_12948_));
 AOI21x1_ASAP7_75t_R _21197_ (.A1(net6211),
    .A2(_12948_),
    .B(net6207),
    .Y(_12950_));
 AOI21x1_ASAP7_75t_R _21198_ (.A1(net6216),
    .A2(net6215),
    .B(net5067),
    .Y(_12951_));
 OAI21x1_ASAP7_75t_R _21200_ (.A1(net4935),
    .A2(_12939_),
    .B(net6202),
    .Y(_12953_));
 AOI21x1_ASAP7_75t_R _21201_ (.A1(_12950_),
    .A2(_12953_),
    .B(net6200),
    .Y(_12954_));
 OAI21x1_ASAP7_75t_R _21202_ (.A1(_12942_),
    .A2(net5189),
    .B(_12954_),
    .Y(_12955_));
 XOR2x2_ASAP7_75t_R _21203_ (.A(_00603_),
    .B(_00635_),
    .Y(_12956_));
 INVx1_ASAP7_75t_R _21204_ (.A(_00700_),
    .Y(_12957_));
 XOR2x2_ASAP7_75t_R _21205_ (.A(_12956_),
    .B(_12957_),
    .Y(_12958_));
 XOR2x2_ASAP7_75t_R _21206_ (.A(_00636_),
    .B(_00668_),
    .Y(_12959_));
 XOR2x2_ASAP7_75t_R _21207_ (.A(_12958_),
    .B(_12959_),
    .Y(_12960_));
 NAND2x1_ASAP7_75t_R _21208_ (.A(net6663),
    .B(_12960_),
    .Y(_12961_));
 OR2x2_ASAP7_75t_R _21210_ (.A(net6663),
    .B(_00537_),
    .Y(_12963_));
 NAND3x1_ASAP7_75t_R _21211_ (.A(_12961_),
    .B(_00955_),
    .C(_12963_),
    .Y(_12964_));
 AO21x1_ASAP7_75t_R _21212_ (.A1(_12961_),
    .A2(_12963_),
    .B(_00955_),
    .Y(_12965_));
 NAND2x1_ASAP7_75t_R _21213_ (.A(_12964_),
    .B(_12965_),
    .Y(_12966_));
 NAND3x1_ASAP7_75t_R _21216_ (.A(_12937_),
    .B(_12955_),
    .C(net5848),
    .Y(_12969_));
 AO21x1_ASAP7_75t_R _21217_ (.A1(net5858),
    .A2(net5295),
    .B(net6204),
    .Y(_12970_));
 AO21x1_ASAP7_75t_R _21218_ (.A1(net6217),
    .A2(net6218),
    .B(_12903_),
    .Y(_12971_));
 AO21x1_ASAP7_75t_R _21220_ (.A1(net6215),
    .A2(net6216),
    .B(net5069),
    .Y(_12973_));
 AO21x1_ASAP7_75t_R _21221_ (.A1(_12971_),
    .A2(net4933),
    .B(net6214),
    .Y(_12974_));
 AOI21x1_ASAP7_75t_R _21223_ (.A1(net5188),
    .A2(_12974_),
    .B(net6207),
    .Y(_12976_));
 AOI21x1_ASAP7_75t_R _21224_ (.A1(net5858),
    .A2(net5864),
    .B(net6213),
    .Y(_12977_));
 NAND2x1_ASAP7_75t_R _21225_ (.A(_12925_),
    .B(_12977_),
    .Y(_12978_));
 NAND2x1_ASAP7_75t_R _21226_ (.A(net5863),
    .B(net5858),
    .Y(_12979_));
 INVx1_ASAP7_75t_R _21227_ (.A(_01132_),
    .Y(_12980_));
 AO21x1_ASAP7_75t_R _21228_ (.A1(net6217),
    .A2(net6218),
    .B(_12980_),
    .Y(_12981_));
 AO21x1_ASAP7_75t_R _21230_ (.A1(_12979_),
    .A2(_12981_),
    .B(net6204),
    .Y(_12983_));
 AOI21x1_ASAP7_75t_R _21232_ (.A1(_12978_),
    .A2(_12983_),
    .B(net5852),
    .Y(_12985_));
 OAI21x1_ASAP7_75t_R _21233_ (.A1(_12976_),
    .A2(_12985_),
    .B(net5850),
    .Y(_12986_));
 INVx1_ASAP7_75t_R _21234_ (.A(_01133_),
    .Y(_12987_));
 AO21x1_ASAP7_75t_R _21235_ (.A1(net6217),
    .A2(net6218),
    .B(_12987_),
    .Y(_12988_));
 NAND2x1_ASAP7_75t_R _21236_ (.A(net6212),
    .B(_12988_),
    .Y(_12989_));
 NAND2x1_ASAP7_75t_R _21237_ (.A(net5859),
    .B(net5864),
    .Y(_12990_));
 NOR2x1_ASAP7_75t_R _21238_ (.A(net5862),
    .B(net5503),
    .Y(_12991_));
 NOR2x1_ASAP7_75t_R _21239_ (.A(net5069),
    .B(net5862),
    .Y(_12992_));
 AOI21x1_ASAP7_75t_R _21240_ (.A1(net6202),
    .A2(_12992_),
    .B(_12916_),
    .Y(_12993_));
 OAI21x1_ASAP7_75t_R _21241_ (.A1(_12989_),
    .A2(_12991_),
    .B(net4691),
    .Y(_12994_));
 NOR2x1_ASAP7_75t_R _21243_ (.A(net6206),
    .B(_12973_),
    .Y(_12996_));
 NOR2x1_ASAP7_75t_R _21244_ (.A(net6207),
    .B(_12996_),
    .Y(_12997_));
 OA21x2_ASAP7_75t_R _21246_ (.A1(net5858),
    .A2(net5068),
    .B(net6205),
    .Y(_12999_));
 OAI21x1_ASAP7_75t_R _21247_ (.A1(net5862),
    .A2(net5503),
    .B(_12999_),
    .Y(_13000_));
 AOI21x1_ASAP7_75t_R _21248_ (.A1(_12997_),
    .A2(_13000_),
    .B(_12935_),
    .Y(_13001_));
 AOI21x1_ASAP7_75t_R _21250_ (.A1(_12994_),
    .A2(_13001_),
    .B(net5848),
    .Y(_13003_));
 XNOR2x2_ASAP7_75t_R _21251_ (.A(net6601),
    .B(net6570),
    .Y(_13004_));
 XOR2x2_ASAP7_75t_R _21252_ (.A(_13004_),
    .B(net6542),
    .Y(_13005_));
 XOR2x2_ASAP7_75t_R _21253_ (.A(_00605_),
    .B(_00637_),
    .Y(_13006_));
 XOR2x2_ASAP7_75t_R _21254_ (.A(_13005_),
    .B(_13006_),
    .Y(_13007_));
 NOR2x1_ASAP7_75t_R _21255_ (.A(net6661),
    .B(_00535_),
    .Y(_13008_));
 AO21x1_ASAP7_75t_R _21256_ (.A1(_13007_),
    .A2(net6662),
    .B(_13008_),
    .Y(_13009_));
 XOR2x2_ASAP7_75t_R _21257_ (.A(_13009_),
    .B(_00958_),
    .Y(_13010_));
 AOI21x1_ASAP7_75t_R _21258_ (.A1(_12986_),
    .A2(_13003_),
    .B(net6199),
    .Y(_13011_));
 NAND2x1_ASAP7_75t_R _21259_ (.A(_12969_),
    .B(_13011_),
    .Y(_13012_));
 NOR2x1_ASAP7_75t_R _21260_ (.A(net5859),
    .B(net5858),
    .Y(_13013_));
 AO21x1_ASAP7_75t_R _21261_ (.A1(net5864),
    .A2(net5859),
    .B(net6204),
    .Y(_13014_));
 NOR2x1_ASAP7_75t_R _21262_ (.A(_13013_),
    .B(_13014_),
    .Y(_13015_));
 INVx1_ASAP7_75t_R _21263_ (.A(_13015_),
    .Y(_13016_));
 AO21x1_ASAP7_75t_R _21265_ (.A1(net5503),
    .A2(_12943_),
    .B(net6212),
    .Y(_13018_));
 AND3x1_ASAP7_75t_R _21266_ (.A(_13016_),
    .B(net5853),
    .C(_13018_),
    .Y(_13019_));
 AO21x1_ASAP7_75t_R _21267_ (.A1(net5864),
    .A2(net5863),
    .B(net5857),
    .Y(_13020_));
 AOI21x1_ASAP7_75t_R _21268_ (.A1(net6216),
    .A2(net6215),
    .B(net4989),
    .Y(_13021_));
 INVx1_ASAP7_75t_R _21269_ (.A(_13021_),
    .Y(_13022_));
 AO21x1_ASAP7_75t_R _21270_ (.A1(_13020_),
    .A2(_13022_),
    .B(net6211),
    .Y(_13023_));
 NOR2x1_ASAP7_75t_R _21271_ (.A(net4932),
    .B(net5862),
    .Y(_13024_));
 INVx1_ASAP7_75t_R _21272_ (.A(_13024_),
    .Y(_13025_));
 NAND2x1_ASAP7_75t_R _21273_ (.A(_12971_),
    .B(_13025_),
    .Y(_13026_));
 AOI21x1_ASAP7_75t_R _21274_ (.A1(net6211),
    .A2(_13026_),
    .B(net5853),
    .Y(_13027_));
 AO21x1_ASAP7_75t_R _21275_ (.A1(_13023_),
    .A2(_13027_),
    .B(net5848),
    .Y(_13028_));
 NAND2x1_ASAP7_75t_R _21276_ (.A(net5860),
    .B(net5864),
    .Y(_13029_));
 NOR2x1p5_ASAP7_75t_R _21277_ (.A(net6212),
    .B(_13021_),
    .Y(_13030_));
 NAND2x1_ASAP7_75t_R _21278_ (.A(_13029_),
    .B(_13030_),
    .Y(_13031_));
 AOI21x1_ASAP7_75t_R _21279_ (.A1(net6218),
    .A2(net6217),
    .B(_12947_),
    .Y(_13032_));
 NOR2x2_ASAP7_75t_R _21280_ (.A(_13032_),
    .B(net6206),
    .Y(_13033_));
 NOR2x1p5_ASAP7_75t_R _21281_ (.A(net6207),
    .B(_13033_),
    .Y(_13034_));
 NAND2x1_ASAP7_75t_R _21282_ (.A(_13031_),
    .B(_13034_),
    .Y(_13035_));
 AOI21x1_ASAP7_75t_R _21283_ (.A1(_13022_),
    .A2(_12971_),
    .B(net6205),
    .Y(_13036_));
 AOI21x1_ASAP7_75t_R _21284_ (.A1(net4524),
    .A2(_12981_),
    .B(net6211),
    .Y(_13037_));
 OAI21x1_ASAP7_75t_R _21286_ (.A1(_13036_),
    .A2(_13037_),
    .B(net6207),
    .Y(_13039_));
 NAND2x1_ASAP7_75t_R _21287_ (.A(_13035_),
    .B(_13039_),
    .Y(_13040_));
 AOI21x1_ASAP7_75t_R _21288_ (.A1(net5848),
    .A2(_13040_),
    .B(_12935_),
    .Y(_13041_));
 OAI21x1_ASAP7_75t_R _21289_ (.A1(_13019_),
    .A2(_13028_),
    .B(_13041_),
    .Y(_13042_));
 AOI21x1_ASAP7_75t_R _21290_ (.A1(net5859),
    .A2(net5862),
    .B(_12894_),
    .Y(_13043_));
 NOR2x1_ASAP7_75t_R _21291_ (.A(net5853),
    .B(net5502),
    .Y(_13044_));
 NOR2x1_ASAP7_75t_R _21292_ (.A(net5295),
    .B(net5860),
    .Y(_13045_));
 AOI21x1_ASAP7_75t_R _21293_ (.A1(net5859),
    .A2(net5864),
    .B(net5857),
    .Y(_13046_));
 OAI21x1_ASAP7_75t_R _21295_ (.A1(net5186),
    .A2(_13046_),
    .B(net6210),
    .Y(_13048_));
 AOI21x1_ASAP7_75t_R _21297_ (.A1(_13044_),
    .A2(_13048_),
    .B(net5848),
    .Y(_13050_));
 NOR2x1_ASAP7_75t_R _21298_ (.A(net5863),
    .B(net5861),
    .Y(_13051_));
 NOR2x1_ASAP7_75t_R _21299_ (.A(_12894_),
    .B(net5864),
    .Y(_13052_));
 NOR2x1_ASAP7_75t_R _21300_ (.A(_13052_),
    .B(_13043_),
    .Y(_13053_));
 INVx1_ASAP7_75t_R _21301_ (.A(_01135_),
    .Y(_13054_));
 AO21x1_ASAP7_75t_R _21302_ (.A1(net6217),
    .A2(net6218),
    .B(_13054_),
    .Y(_13055_));
 OA21x2_ASAP7_75t_R _21303_ (.A1(net5860),
    .A2(_12947_),
    .B(net6211),
    .Y(_13056_));
 AOI21x1_ASAP7_75t_R _21304_ (.A1(net4931),
    .A2(_13056_),
    .B(net6207),
    .Y(_13057_));
 OAI21x1_ASAP7_75t_R _21305_ (.A1(_13051_),
    .A2(net5185),
    .B(_13057_),
    .Y(_13058_));
 AOI21x1_ASAP7_75t_R _21307_ (.A1(_13050_),
    .A2(_13058_),
    .B(net6200),
    .Y(_13060_));
 INVx1_ASAP7_75t_R _21308_ (.A(_12945_),
    .Y(_13061_));
 NOR2x1_ASAP7_75t_R _21309_ (.A(_12874_),
    .B(net5864),
    .Y(_13062_));
 NAND2x1_ASAP7_75t_R _21310_ (.A(net6204),
    .B(_13062_),
    .Y(_13063_));
 AND2x2_ASAP7_75t_R _21311_ (.A(_12993_),
    .B(_13063_),
    .Y(_13064_));
 NAND2x1_ASAP7_75t_R _21312_ (.A(_13061_),
    .B(_13064_),
    .Y(_13065_));
 INVx4_ASAP7_75t_R _21313_ (.A(_12832_),
    .Y(_01125_));
 NOR2x1_ASAP7_75t_R _21314_ (.A(net5860),
    .B(net5496),
    .Y(_13066_));
 OAI21x1_ASAP7_75t_R _21316_ (.A1(_13046_),
    .A2(_13066_),
    .B(net6201),
    .Y(_13068_));
 NAND2x1_ASAP7_75t_R _21317_ (.A(net5859),
    .B(net5860),
    .Y(_13069_));
 AO21x2_ASAP7_75t_R _21318_ (.A1(net6215),
    .A2(net6216),
    .B(_13054_),
    .Y(_13070_));
 AND2x2_ASAP7_75t_R _21319_ (.A(_13070_),
    .B(net6211),
    .Y(_13071_));
 AOI21x1_ASAP7_75t_R _21320_ (.A1(_13069_),
    .A2(_13071_),
    .B(net6207),
    .Y(_13072_));
 INVx1_ASAP7_75t_R _21321_ (.A(_12966_),
    .Y(_13073_));
 AOI21x1_ASAP7_75t_R _21322_ (.A1(_13068_),
    .A2(_13072_),
    .B(net5494),
    .Y(_13074_));
 NAND2x1_ASAP7_75t_R _21323_ (.A(_13065_),
    .B(_13074_),
    .Y(_13075_));
 INVx1_ASAP7_75t_R _21324_ (.A(_13010_),
    .Y(_13076_));
 AOI21x1_ASAP7_75t_R _21325_ (.A1(_13060_),
    .A2(_13075_),
    .B(_13076_),
    .Y(_13077_));
 NAND2x1_ASAP7_75t_R _21326_ (.A(_13042_),
    .B(_13077_),
    .Y(_13078_));
 NAND2x1_ASAP7_75t_R _21327_ (.A(_13012_),
    .B(_13078_),
    .Y(_00056_));
 NOR2x1_ASAP7_75t_R _21328_ (.A(_13062_),
    .B(_12970_),
    .Y(_13079_));
 INVx1_ASAP7_75t_R _21329_ (.A(_12971_),
    .Y(_13080_));
 OA21x2_ASAP7_75t_R _21331_ (.A1(_13080_),
    .A2(_13051_),
    .B(net6203),
    .Y(_13082_));
 OAI21x1_ASAP7_75t_R _21333_ (.A1(net4930),
    .A2(_13082_),
    .B(net6207),
    .Y(_13084_));
 AO21x1_ASAP7_75t_R _21334_ (.A1(net5505),
    .A2(net4933),
    .B(net6214),
    .Y(_13085_));
 AO21x1_ASAP7_75t_R _21335_ (.A1(net4581),
    .A2(net4524),
    .B(net6203),
    .Y(_13086_));
 AO21x1_ASAP7_75t_R _21336_ (.A1(_13085_),
    .A2(_13086_),
    .B(net6207),
    .Y(_13087_));
 AOI21x1_ASAP7_75t_R _21337_ (.A1(_13084_),
    .A2(_13087_),
    .B(net5848),
    .Y(_13088_));
 NAND2x1_ASAP7_75t_R _21338_ (.A(net5859),
    .B(net6206),
    .Y(_13089_));
 INVx1_ASAP7_75t_R _21339_ (.A(_12977_),
    .Y(_13090_));
 NAND2x1_ASAP7_75t_R _21340_ (.A(_13089_),
    .B(_13090_),
    .Y(_13091_));
 AO21x1_ASAP7_75t_R _21341_ (.A1(_12948_),
    .A2(net6211),
    .B(net5854),
    .Y(_13092_));
 AOI21x1_ASAP7_75t_R _21342_ (.A1(_13069_),
    .A2(_13091_),
    .B(_13092_),
    .Y(_13093_));
 AND3x1_ASAP7_75t_R _21343_ (.A(net6215),
    .B(net6216),
    .C(net5069),
    .Y(_13094_));
 NAND2x1_ASAP7_75t_R _21344_ (.A(net6202),
    .B(_13070_),
    .Y(_13095_));
 OAI21x1_ASAP7_75t_R _21346_ (.A1(_13094_),
    .A2(_13095_),
    .B(_12916_),
    .Y(_13097_));
 NAND2x1_ASAP7_75t_R _21348_ (.A(net5863),
    .B(net5864),
    .Y(_13099_));
 NOR2x1p5_ASAP7_75t_R _21349_ (.A(net5860),
    .B(net4765),
    .Y(_13100_));
 AOI21x1_ASAP7_75t_R _21350_ (.A1(net5862),
    .A2(net5491),
    .B(net4577),
    .Y(_13101_));
 NOR2x1_ASAP7_75t_R _21351_ (.A(net6202),
    .B(_13101_),
    .Y(_13102_));
 OAI21x1_ASAP7_75t_R _21352_ (.A1(_13097_),
    .A2(_13102_),
    .B(net5848),
    .Y(_13103_));
 OAI21x1_ASAP7_75t_R _21354_ (.A1(_13093_),
    .A2(_13103_),
    .B(net5849),
    .Y(_13105_));
 OAI21x1_ASAP7_75t_R _21355_ (.A1(_13088_),
    .A2(_13105_),
    .B(net6199),
    .Y(_13106_));
 AND2x2_ASAP7_75t_R _21357_ (.A(net5848),
    .B(_01142_),
    .Y(_13108_));
 AO21x1_ASAP7_75t_R _21358_ (.A1(net6217),
    .A2(net6218),
    .B(net5068),
    .Y(_13109_));
 NAND2x1_ASAP7_75t_R _21359_ (.A(net6202),
    .B(_13109_),
    .Y(_13110_));
 NOR2x1_ASAP7_75t_R _21360_ (.A(net5861),
    .B(_13099_),
    .Y(_13111_));
 OAI21x1_ASAP7_75t_R _21361_ (.A1(_13110_),
    .A2(_13111_),
    .B(net6207),
    .Y(_13112_));
 AO21x1_ASAP7_75t_R _21362_ (.A1(net6214),
    .A2(_13108_),
    .B(_13112_),
    .Y(_13113_));
 INVx1_ASAP7_75t_R _21363_ (.A(_13046_),
    .Y(_13114_));
 NAND2x1_ASAP7_75t_R _21364_ (.A(_13114_),
    .B(net5504),
    .Y(_13115_));
 AO21x1_ASAP7_75t_R _21365_ (.A1(net5862),
    .A2(_12903_),
    .B(net6212),
    .Y(_13116_));
 OAI21x1_ASAP7_75t_R _21367_ (.A1(_13051_),
    .A2(_13116_),
    .B(net5493),
    .Y(_13118_));
 AOI21x1_ASAP7_75t_R _21368_ (.A1(net6214),
    .A2(_13115_),
    .B(_13118_),
    .Y(_13119_));
 AND3x1_ASAP7_75t_R _21369_ (.A(_13029_),
    .B(net6203),
    .C(_12979_),
    .Y(_13120_));
 NOR3x1_ASAP7_75t_R _21371_ (.A(_13120_),
    .B(net5493),
    .C(_13079_),
    .Y(_13122_));
 OAI21x1_ASAP7_75t_R _21372_ (.A1(_13119_),
    .A2(_13122_),
    .B(net5851),
    .Y(_13123_));
 AOI21x1_ASAP7_75t_R _21373_ (.A1(_13113_),
    .A2(_13123_),
    .B(net5850),
    .Y(_13124_));
 AOI21x1_ASAP7_75t_R _21374_ (.A1(net5190),
    .A2(_12881_),
    .B(net6209),
    .Y(_13125_));
 AO21x1_ASAP7_75t_R _21375_ (.A1(_13070_),
    .A2(net4477),
    .B(net5854),
    .Y(_13126_));
 NOR2x1_ASAP7_75t_R _21376_ (.A(net5860),
    .B(net5864),
    .Y(_13127_));
 AOI21x1_ASAP7_75t_R _21377_ (.A1(net6212),
    .A2(_13029_),
    .B(_13127_),
    .Y(_13128_));
 OA21x2_ASAP7_75t_R _21378_ (.A1(net5191),
    .A2(net6211),
    .B(net5856),
    .Y(_13129_));
 AOI21x1_ASAP7_75t_R _21379_ (.A1(_13128_),
    .A2(_13129_),
    .B(net5494),
    .Y(_13130_));
 OAI21x1_ASAP7_75t_R _21380_ (.A1(_13125_),
    .A2(_13126_),
    .B(_13130_),
    .Y(_13131_));
 NOR2x1_ASAP7_75t_R _21381_ (.A(net5863),
    .B(net5864),
    .Y(_13132_));
 INVx1_ASAP7_75t_R _21382_ (.A(_13132_),
    .Y(_13133_));
 NAND2x1_ASAP7_75t_R _21383_ (.A(_12977_),
    .B(_13133_),
    .Y(_13134_));
 NAND2x1_ASAP7_75t_R _21384_ (.A(net5861),
    .B(net6213),
    .Y(_13135_));
 INVx1_ASAP7_75t_R _21385_ (.A(_13135_),
    .Y(_13136_));
 AOI21x1_ASAP7_75t_R _21386_ (.A1(net5503),
    .A2(_13136_),
    .B(net5852),
    .Y(_13137_));
 AOI21x1_ASAP7_75t_R _21387_ (.A1(_13134_),
    .A2(_13137_),
    .B(net5848),
    .Y(_13138_));
 INVx1_ASAP7_75t_R _21388_ (.A(net5295),
    .Y(_13139_));
 OA21x2_ASAP7_75t_R _21389_ (.A1(net5862),
    .A2(_13139_),
    .B(net6205),
    .Y(_13140_));
 NAND2x1_ASAP7_75t_R _21390_ (.A(net5505),
    .B(_13140_),
    .Y(_13141_));
 AOI21x1_ASAP7_75t_R _21391_ (.A1(_13069_),
    .A2(_13056_),
    .B(net6207),
    .Y(_13142_));
 NAND2x1_ASAP7_75t_R _21392_ (.A(_13141_),
    .B(_13142_),
    .Y(_13143_));
 AOI21x1_ASAP7_75t_R _21393_ (.A1(_13138_),
    .A2(_13143_),
    .B(net5849),
    .Y(_13144_));
 AOI21x1_ASAP7_75t_R _21394_ (.A1(_13131_),
    .A2(_13144_),
    .B(net6199),
    .Y(_13145_));
 NAND2x1_ASAP7_75t_R _21395_ (.A(net5859),
    .B(net5857),
    .Y(_13146_));
 NOR2x1_ASAP7_75t_R _21396_ (.A(net6212),
    .B(_12924_),
    .Y(_13147_));
 AOI21x1_ASAP7_75t_R _21397_ (.A1(_13146_),
    .A2(_13147_),
    .B(net5856),
    .Y(_13148_));
 AO21x1_ASAP7_75t_R _21398_ (.A1(net5491),
    .A2(_13146_),
    .B(net6202),
    .Y(_13149_));
 AOI21x1_ASAP7_75t_R _21399_ (.A1(_13148_),
    .A2(_13149_),
    .B(net5495),
    .Y(_13150_));
 NOR2x1_ASAP7_75t_R _21400_ (.A(net6211),
    .B(_12906_),
    .Y(_13151_));
 AND3x1_ASAP7_75t_R _21401_ (.A(net5191),
    .B(_12948_),
    .C(net6211),
    .Y(_13152_));
 OAI21x1_ASAP7_75t_R _21402_ (.A1(_13151_),
    .A2(_13152_),
    .B(net5855),
    .Y(_13153_));
 NAND2x1_ASAP7_75t_R _21403_ (.A(_13150_),
    .B(_13153_),
    .Y(_13154_));
 INVx1_ASAP7_75t_R _21404_ (.A(_13045_),
    .Y(_13155_));
 OA21x2_ASAP7_75t_R _21405_ (.A1(_13155_),
    .A2(net6211),
    .B(net6207),
    .Y(_13156_));
 OAI21x1_ASAP7_75t_R _21406_ (.A1(net6202),
    .A2(_13101_),
    .B(_13156_),
    .Y(_13157_));
 OA21x2_ASAP7_75t_R _21407_ (.A1(_12823_),
    .A2(_12811_),
    .B(_12830_),
    .Y(_13158_));
 OA21x2_ASAP7_75t_R _21408_ (.A1(_12829_),
    .A2(_12826_),
    .B(_00951_),
    .Y(_13159_));
 OAI21x1_ASAP7_75t_R _21409_ (.A1(_13158_),
    .A2(_13159_),
    .B(_12874_),
    .Y(_13160_));
 AO21x1_ASAP7_75t_R _21410_ (.A1(net5488),
    .A2(_13146_),
    .B(net6211),
    .Y(_13161_));
 OA21x2_ASAP7_75t_R _21411_ (.A1(net5857),
    .A2(_13054_),
    .B(net6211),
    .Y(_13162_));
 AOI21x1_ASAP7_75t_R _21412_ (.A1(net5488),
    .A2(_13162_),
    .B(net6207),
    .Y(_13163_));
 AOI21x1_ASAP7_75t_R _21413_ (.A1(_13161_),
    .A2(_13163_),
    .B(net5848),
    .Y(_13164_));
 AOI21x1_ASAP7_75t_R _21414_ (.A1(_13157_),
    .A2(_13164_),
    .B(net6200),
    .Y(_13165_));
 NAND2x1_ASAP7_75t_R _21415_ (.A(_13154_),
    .B(_13165_),
    .Y(_13166_));
 NAND2x1_ASAP7_75t_R _21416_ (.A(_13166_),
    .B(_13145_),
    .Y(_13167_));
 OAI21x1_ASAP7_75t_R _21417_ (.A1(_13106_),
    .A2(_13124_),
    .B(_13167_),
    .Y(_00057_));
 INVx1_ASAP7_75t_R _21418_ (.A(_13066_),
    .Y(_13168_));
 AOI21x1_ASAP7_75t_R _21419_ (.A1(net4582),
    .A2(_13168_),
    .B(net6211),
    .Y(_13169_));
 AOI21x1_ASAP7_75t_R _21420_ (.A1(net5190),
    .A2(_12881_),
    .B(net6201),
    .Y(_13170_));
 OAI21x1_ASAP7_75t_R _21421_ (.A1(_13169_),
    .A2(_13170_),
    .B(net6207),
    .Y(_13171_));
 INVx1_ASAP7_75t_R _21422_ (.A(_13055_),
    .Y(_13172_));
 AO21x1_ASAP7_75t_R _21423_ (.A1(net5857),
    .A2(net5295),
    .B(net6211),
    .Y(_13173_));
 NOR2x1_ASAP7_75t_R _21424_ (.A(_13172_),
    .B(_13173_),
    .Y(_13174_));
 OAI21x1_ASAP7_75t_R _21425_ (.A1(_13127_),
    .A2(_13046_),
    .B(net6211),
    .Y(_13175_));
 INVx1_ASAP7_75t_R _21426_ (.A(_13175_),
    .Y(_13176_));
 OAI21x1_ASAP7_75t_R _21427_ (.A1(_13174_),
    .A2(_13176_),
    .B(net5853),
    .Y(_13177_));
 NAND3x1_ASAP7_75t_R _21428_ (.A(_13171_),
    .B(_13177_),
    .C(net5848),
    .Y(_13178_));
 NOR2x1_ASAP7_75t_R _21429_ (.A(net5294),
    .B(net5860),
    .Y(_13179_));
 INVx1_ASAP7_75t_R _21430_ (.A(_13179_),
    .Y(_13180_));
 AOI21x1_ASAP7_75t_R _21431_ (.A1(_13180_),
    .A2(_13020_),
    .B(net6201),
    .Y(_13181_));
 NAND2x1_ASAP7_75t_R _21433_ (.A(net6207),
    .B(net5185),
    .Y(_13183_));
 AOI22x1_ASAP7_75t_R _21434_ (.A1(net6219),
    .A2(_12847_),
    .B1(net6215),
    .B2(net6216),
    .Y(_13184_));
 OAI21x1_ASAP7_75t_R _21435_ (.A1(net5069),
    .A2(net5857),
    .B(net6211),
    .Y(_13185_));
 NOR2x1_ASAP7_75t_R _21436_ (.A(_13184_),
    .B(_13185_),
    .Y(_13186_));
 AOI21x1_ASAP7_75t_R _21437_ (.A1(_12948_),
    .A2(_13029_),
    .B(net6211),
    .Y(_13187_));
 OAI21x1_ASAP7_75t_R _21438_ (.A1(_13186_),
    .A2(_13187_),
    .B(net5855),
    .Y(_13188_));
 OAI21x1_ASAP7_75t_R _21439_ (.A1(_13181_),
    .A2(_13183_),
    .B(_13188_),
    .Y(_13189_));
 AOI21x1_ASAP7_75t_R _21440_ (.A1(net5495),
    .A2(_13189_),
    .B(net5849),
    .Y(_13190_));
 OAI21x1_ASAP7_75t_R _21441_ (.A1(net5066),
    .A2(net5860),
    .B(net6211),
    .Y(_13191_));
 NOR2x1_ASAP7_75t_R _21442_ (.A(net5497),
    .B(_13191_),
    .Y(_13192_));
 OAI21x1_ASAP7_75t_R _21443_ (.A1(net5294),
    .A2(net5857),
    .B(net6202),
    .Y(_13193_));
 OAI21x1_ASAP7_75t_R _21444_ (.A1(_13184_),
    .A2(_13193_),
    .B(net5856),
    .Y(_13194_));
 NOR2x1_ASAP7_75t_R _21445_ (.A(_13192_),
    .B(_13194_),
    .Y(_13195_));
 OAI21x1_ASAP7_75t_R _21446_ (.A1(net4578),
    .A2(net4764),
    .B(net6209),
    .Y(_13196_));
 NOR2x1_ASAP7_75t_R _21447_ (.A(net5066),
    .B(net5857),
    .Y(_13197_));
 OAI21x1_ASAP7_75t_R _21448_ (.A1(_13184_),
    .A2(_13197_),
    .B(net6201),
    .Y(_13198_));
 AOI21x1_ASAP7_75t_R _21449_ (.A1(_13196_),
    .A2(_13198_),
    .B(net5855),
    .Y(_13199_));
 OAI21x1_ASAP7_75t_R _21450_ (.A1(_13195_),
    .A2(_13199_),
    .B(net5495),
    .Y(_13200_));
 NOR2x1_ASAP7_75t_R _21451_ (.A(net5294),
    .B(net5857),
    .Y(_13201_));
 OAI21x1_ASAP7_75t_R _21452_ (.A1(net4935),
    .A2(_13201_),
    .B(net6202),
    .Y(_13202_));
 AOI21x1_ASAP7_75t_R _21453_ (.A1(net5295),
    .A2(net5860),
    .B(net6202),
    .Y(_13203_));
 NAND2x1_ASAP7_75t_R _21454_ (.A(_13146_),
    .B(_13203_),
    .Y(_13204_));
 AOI21x1_ASAP7_75t_R _21455_ (.A1(_13202_),
    .A2(_13204_),
    .B(net6207),
    .Y(_13205_));
 NAND2x1_ASAP7_75t_R _21456_ (.A(net5488),
    .B(_13203_),
    .Y(_13206_));
 AOI21x1_ASAP7_75t_R _21457_ (.A1(_13206_),
    .A2(net4693),
    .B(net5855),
    .Y(_13207_));
 OAI21x1_ASAP7_75t_R _21458_ (.A1(_13205_),
    .A2(_13207_),
    .B(net5848),
    .Y(_13208_));
 AOI21x1_ASAP7_75t_R _21460_ (.A1(_13200_),
    .A2(_13208_),
    .B(net6200),
    .Y(_13210_));
 AOI21x1_ASAP7_75t_R _21461_ (.A1(_13178_),
    .A2(_13190_),
    .B(_13210_),
    .Y(_13211_));
 AO21x1_ASAP7_75t_R _21462_ (.A1(net6215),
    .A2(net6216),
    .B(_12878_),
    .Y(_13212_));
 AOI21x1_ASAP7_75t_R _21463_ (.A1(net4688),
    .A2(_13020_),
    .B(net6201),
    .Y(_13213_));
 OAI21x1_ASAP7_75t_R _21464_ (.A1(net4690),
    .A2(_13111_),
    .B(net5856),
    .Y(_13214_));
 OAI21x1_ASAP7_75t_R _21465_ (.A1(net4764),
    .A2(net4936),
    .B(net6208),
    .Y(_13215_));
 OA21x2_ASAP7_75t_R _21466_ (.A1(net4524),
    .A2(net6208),
    .B(net6207),
    .Y(_13216_));
 AOI21x1_ASAP7_75t_R _21467_ (.A1(_13215_),
    .A2(_13216_),
    .B(net5848),
    .Y(_13217_));
 OAI21x1_ASAP7_75t_R _21468_ (.A1(_13213_),
    .A2(_13214_),
    .B(_13217_),
    .Y(_13218_));
 OA21x2_ASAP7_75t_R _21469_ (.A1(_01144_),
    .A2(net6211),
    .B(net5853),
    .Y(_13219_));
 AOI21x1_ASAP7_75t_R _21470_ (.A1(_13219_),
    .A2(_13175_),
    .B(net5494),
    .Y(_13220_));
 NAND2x1_ASAP7_75t_R _21471_ (.A(_01139_),
    .B(net6211),
    .Y(_13221_));
 NAND3x1_ASAP7_75t_R _21472_ (.A(net5185),
    .B(net6207),
    .C(_13221_),
    .Y(_13222_));
 NAND2x1_ASAP7_75t_R _21473_ (.A(_13220_),
    .B(_13222_),
    .Y(_13223_));
 AOI21x1_ASAP7_75t_R _21474_ (.A1(_13218_),
    .A2(_13223_),
    .B(net5849),
    .Y(_13224_));
 NAND2x1_ASAP7_75t_R _21475_ (.A(net5863),
    .B(net6212),
    .Y(_13225_));
 AO21x1_ASAP7_75t_R _21476_ (.A1(_13225_),
    .A2(_13135_),
    .B(net5500),
    .Y(_13226_));
 NAND2x1_ASAP7_75t_R _21477_ (.A(_12978_),
    .B(_13226_),
    .Y(_13227_));
 OA21x2_ASAP7_75t_R _21478_ (.A1(_01140_),
    .A2(net6211),
    .B(net6207),
    .Y(_13228_));
 OAI21x1_ASAP7_75t_R _21479_ (.A1(net5860),
    .A2(net5503),
    .B(net4476),
    .Y(_13229_));
 AOI21x1_ASAP7_75t_R _21480_ (.A1(_13229_),
    .A2(_13228_),
    .B(net5848),
    .Y(_13230_));
 OAI21x1_ASAP7_75t_R _21481_ (.A1(net6207),
    .A2(_13227_),
    .B(_13230_),
    .Y(_13231_));
 NOR3x1_ASAP7_75t_R _21482_ (.A(_13024_),
    .B(net6205),
    .C(net4766),
    .Y(_13232_));
 NOR2x1_ASAP7_75t_R _21483_ (.A(_13080_),
    .B(_13090_),
    .Y(_13233_));
 OAI21x1_ASAP7_75t_R _21484_ (.A1(_13232_),
    .A2(_13233_),
    .B(net5852),
    .Y(_13234_));
 NAND2x1_ASAP7_75t_R _21485_ (.A(_01142_),
    .B(net6204),
    .Y(_13235_));
 AOI21x1_ASAP7_75t_R _21486_ (.A1(net5858),
    .A2(net5864),
    .B(net6204),
    .Y(_13236_));
 AOI21x1_ASAP7_75t_R _21487_ (.A1(_13236_),
    .A2(_13133_),
    .B(net5851),
    .Y(_13237_));
 AOI21x1_ASAP7_75t_R _21488_ (.A1(_13235_),
    .A2(_13237_),
    .B(net5493),
    .Y(_13238_));
 NAND2x1_ASAP7_75t_R _21489_ (.A(_13234_),
    .B(_13238_),
    .Y(_13239_));
 AOI21x1_ASAP7_75t_R _21490_ (.A1(_13231_),
    .A2(_13239_),
    .B(net6200),
    .Y(_13240_));
 OAI21x1_ASAP7_75t_R _21491_ (.A1(_13240_),
    .A2(_13224_),
    .B(_13076_),
    .Y(_13241_));
 OAI21x1_ASAP7_75t_R _21492_ (.A1(_13076_),
    .A2(_13211_),
    .B(_13241_),
    .Y(_00058_));
 AO21x1_ASAP7_75t_R _21493_ (.A1(net6217),
    .A2(net6218),
    .B(net5294),
    .Y(_13242_));
 AO21x1_ASAP7_75t_R _21494_ (.A1(_13212_),
    .A2(_13242_),
    .B(net6202),
    .Y(_13243_));
 NAND2x1_ASAP7_75t_R _21495_ (.A(_12948_),
    .B(net5502),
    .Y(_13244_));
 NAND3x1_ASAP7_75t_R _21496_ (.A(_13243_),
    .B(_13244_),
    .C(net5848),
    .Y(_13245_));
 INVx1_ASAP7_75t_R _21497_ (.A(_12951_),
    .Y(_13246_));
 OA21x2_ASAP7_75t_R _21498_ (.A1(net6201),
    .A2(_13246_),
    .B(_13073_),
    .Y(_13247_));
 AOI21x1_ASAP7_75t_R _21499_ (.A1(_13198_),
    .A2(_13247_),
    .B(net5855),
    .Y(_13248_));
 AOI21x1_ASAP7_75t_R _21500_ (.A1(_13245_),
    .A2(_13248_),
    .B(net5849),
    .Y(_13249_));
 INVx1_ASAP7_75t_R _21501_ (.A(net4578),
    .Y(_13250_));
 NOR2x1_ASAP7_75t_R _21502_ (.A(net6201),
    .B(_13250_),
    .Y(_13251_));
 NOR2x1_ASAP7_75t_R _21503_ (.A(_13066_),
    .B(_13110_),
    .Y(_13252_));
 OAI21x1_ASAP7_75t_R _21504_ (.A1(_13251_),
    .A2(_13252_),
    .B(net5848),
    .Y(_13253_));
 NAND2x1p5_ASAP7_75t_R _21505_ (.A(_13100_),
    .B(net6205),
    .Y(_13254_));
 INVx1_ASAP7_75t_R _21506_ (.A(_12996_),
    .Y(_13255_));
 OA21x2_ASAP7_75t_R _21507_ (.A1(_13254_),
    .A2(net5848),
    .B(_13255_),
    .Y(_13256_));
 AO21x1_ASAP7_75t_R _21508_ (.A1(_13253_),
    .A2(_13256_),
    .B(net6207),
    .Y(_13257_));
 NAND2x1_ASAP7_75t_R _21509_ (.A(_13249_),
    .B(_13257_),
    .Y(_13258_));
 AO21x1_ASAP7_75t_R _21510_ (.A1(net6217),
    .A2(net6218),
    .B(net5067),
    .Y(_13259_));
 AOI21x1_ASAP7_75t_R _21511_ (.A1(_13259_),
    .A2(_13212_),
    .B(net6202),
    .Y(_13260_));
 INVx1_ASAP7_75t_R _21512_ (.A(_13193_),
    .Y(_13261_));
 NAND2x1_ASAP7_75t_R _21513_ (.A(_12979_),
    .B(_13261_),
    .Y(_13262_));
 OA21x2_ASAP7_75t_R _21514_ (.A1(_13262_),
    .A2(net6207),
    .B(net5848),
    .Y(_13263_));
 OAI21x1_ASAP7_75t_R _21515_ (.A1(_13112_),
    .A2(net4523),
    .B(_13263_),
    .Y(_13264_));
 NAND2x1p5_ASAP7_75t_R _21516_ (.A(_13254_),
    .B(_13191_),
    .Y(_13265_));
 OA21x2_ASAP7_75t_R _21517_ (.A1(_13135_),
    .A2(net5863),
    .B(net5856),
    .Y(_13266_));
 OAI21x1_ASAP7_75t_R _21518_ (.A1(net4689),
    .A2(_13265_),
    .B(_13266_),
    .Y(_13267_));
 AOI21x1_ASAP7_75t_R _21519_ (.A1(_13134_),
    .A2(_12919_),
    .B(net5848),
    .Y(_13268_));
 AOI21x1_ASAP7_75t_R _21520_ (.A1(_13267_),
    .A2(_13268_),
    .B(net6200),
    .Y(_13269_));
 AOI21x1_ASAP7_75t_R _21521_ (.A1(_13264_),
    .A2(_13269_),
    .B(_13076_),
    .Y(_13270_));
 NAND2x1_ASAP7_75t_R _21522_ (.A(_13258_),
    .B(_13270_),
    .Y(_13271_));
 NOR2x1_ASAP7_75t_R _21523_ (.A(_13024_),
    .B(_13013_),
    .Y(_13272_));
 AOI22x1_ASAP7_75t_R _21524_ (.A1(_13272_),
    .A2(net6202),
    .B1(net4524),
    .B2(net4477),
    .Y(_13273_));
 NOR2x1_ASAP7_75t_R _21525_ (.A(net6207),
    .B(_13273_),
    .Y(_13274_));
 AO21x1_ASAP7_75t_R _21526_ (.A1(_13070_),
    .A2(_13203_),
    .B(_13187_),
    .Y(_13275_));
 OAI21x1_ASAP7_75t_R _21527_ (.A1(net5856),
    .A2(_13275_),
    .B(net6200),
    .Y(_13276_));
 NOR2x1_ASAP7_75t_R _21528_ (.A(_13274_),
    .B(_13276_),
    .Y(_13277_));
 NOR2x1_ASAP7_75t_R _21529_ (.A(net6213),
    .B(net4577),
    .Y(_13278_));
 AOI21x1_ASAP7_75t_R _21530_ (.A1(_12981_),
    .A2(_13278_),
    .B(net6207),
    .Y(_13279_));
 AOI21x1_ASAP7_75t_R _21531_ (.A1(net4576),
    .A2(net5504),
    .B(net5851),
    .Y(_13280_));
 NOR2x1_ASAP7_75t_R _21532_ (.A(net6203),
    .B(net5498),
    .Y(_13281_));
 NAND2x1_ASAP7_75t_R _21533_ (.A(_13272_),
    .B(_13281_),
    .Y(_13282_));
 AOI22x1_ASAP7_75t_R _21534_ (.A1(_13016_),
    .A2(_13279_),
    .B1(_13280_),
    .B2(_13282_),
    .Y(_13283_));
 OAI21x1_ASAP7_75t_R _21535_ (.A1(net6200),
    .A2(_13283_),
    .B(net5494),
    .Y(_13284_));
 AND3x1_ASAP7_75t_R _21536_ (.A(net5503),
    .B(net6204),
    .C(_12979_),
    .Y(_13285_));
 INVx1_ASAP7_75t_R _21537_ (.A(net5500),
    .Y(_13286_));
 AO21x1_ASAP7_75t_R _21538_ (.A1(_13056_),
    .A2(_13286_),
    .B(net5852),
    .Y(_13287_));
 AO21x1_ASAP7_75t_R _21539_ (.A1(_13029_),
    .A2(_12979_),
    .B(net6213),
    .Y(_13288_));
 AOI21x1_ASAP7_75t_R _21540_ (.A1(net4434),
    .A2(_13288_),
    .B(_12935_),
    .Y(_13289_));
 OAI21x1_ASAP7_75t_R _21541_ (.A1(_13285_),
    .A2(_13287_),
    .B(_13289_),
    .Y(_13290_));
 NAND2x1_ASAP7_75t_R _21542_ (.A(net4692),
    .B(net4580),
    .Y(_13291_));
 NAND2x1_ASAP7_75t_R _21543_ (.A(_13291_),
    .B(_13163_),
    .Y(_13292_));
 NAND2x1_ASAP7_75t_R _21544_ (.A(net5858),
    .B(net6212),
    .Y(_13293_));
 OAI21x1_ASAP7_75t_R _21545_ (.A1(net5859),
    .A2(net5858),
    .B(net6207),
    .Y(_13294_));
 NOR2x1_ASAP7_75t_R _21546_ (.A(net5489),
    .B(_13294_),
    .Y(_13295_));
 AOI21x1_ASAP7_75t_R _21547_ (.A1(_13293_),
    .A2(_13295_),
    .B(net6200),
    .Y(_13296_));
 AOI21x1_ASAP7_75t_R _21548_ (.A1(_13292_),
    .A2(_13296_),
    .B(net5493),
    .Y(_13297_));
 AOI21x1_ASAP7_75t_R _21549_ (.A1(_13290_),
    .A2(_13297_),
    .B(net6199),
    .Y(_13298_));
 OAI21x1_ASAP7_75t_R _21550_ (.A1(_13277_),
    .A2(_13284_),
    .B(_13298_),
    .Y(_13299_));
 NAND2x1_ASAP7_75t_R _21551_ (.A(_13271_),
    .B(_13299_),
    .Y(_00059_));
 INVx1_ASAP7_75t_R _21552_ (.A(_01134_),
    .Y(_13300_));
 NAND2x1_ASAP7_75t_R _21553_ (.A(_13300_),
    .B(net6203),
    .Y(_13301_));
 OAI21x1_ASAP7_75t_R _21554_ (.A1(net6203),
    .A2(net4581),
    .B(_13301_),
    .Y(_13302_));
 AO21x1_ASAP7_75t_R _21555_ (.A1(_13302_),
    .A2(net6207),
    .B(net5848),
    .Y(_13303_));
 OA21x2_ASAP7_75t_R _21556_ (.A1(net5857),
    .A2(_12987_),
    .B(net6212),
    .Y(_13304_));
 NAND2x1_ASAP7_75t_R _21557_ (.A(_13160_),
    .B(_13304_),
    .Y(_13305_));
 INVx1_ASAP7_75t_R _21558_ (.A(_13305_),
    .Y(_13306_));
 AOI21x1_ASAP7_75t_R _21559_ (.A1(net6202),
    .A2(_13184_),
    .B(net6207),
    .Y(_13307_));
 OAI21x1_ASAP7_75t_R _21560_ (.A1(net6211),
    .A2(_13160_),
    .B(_13307_),
    .Y(_13308_));
 NOR2x1_ASAP7_75t_R _21561_ (.A(_13306_),
    .B(_13308_),
    .Y(_13309_));
 OAI21x1_ASAP7_75t_R _21562_ (.A1(_13303_),
    .A2(_13309_),
    .B(net6200),
    .Y(_13310_));
 NOR2x1_ASAP7_75t_R _21563_ (.A(net6212),
    .B(net5499),
    .Y(_13311_));
 NOR2x1_ASAP7_75t_R _21564_ (.A(_13184_),
    .B(_12989_),
    .Y(_13312_));
 AOI211x1_ASAP7_75t_R _21565_ (.A1(_12990_),
    .A2(_13311_),
    .B(_13312_),
    .C(net6207),
    .Y(_13313_));
 OAI21x1_ASAP7_75t_R _21566_ (.A1(net6212),
    .A2(_12971_),
    .B(net4691),
    .Y(_13314_));
 OAI21x1_ASAP7_75t_R _21567_ (.A1(net5187),
    .A2(_13314_),
    .B(net5848),
    .Y(_13315_));
 NOR2x1_ASAP7_75t_R _21568_ (.A(_13313_),
    .B(_13315_),
    .Y(_13316_));
 OAI21x1_ASAP7_75t_R _21569_ (.A1(_13310_),
    .A2(_13316_),
    .B(net6199),
    .Y(_13317_));
 OAI21x1_ASAP7_75t_R _21570_ (.A1(net6211),
    .A2(_13094_),
    .B(_12916_),
    .Y(_13318_));
 OA21x2_ASAP7_75t_R _21571_ (.A1(net5491),
    .A2(net5857),
    .B(net6211),
    .Y(_13319_));
 NOR2x1_ASAP7_75t_R _21572_ (.A(_13318_),
    .B(_13319_),
    .Y(_13320_));
 OAI21x1_ASAP7_75t_R _21573_ (.A1(_12924_),
    .A2(_13173_),
    .B(net6207),
    .Y(_13321_));
 NOR2x1_ASAP7_75t_R _21574_ (.A(_13321_),
    .B(net5189),
    .Y(_13322_));
 OAI21x1_ASAP7_75t_R _21575_ (.A1(_13320_),
    .A2(_13322_),
    .B(net5493),
    .Y(_13323_));
 NOR2x1_ASAP7_75t_R _21576_ (.A(net5493),
    .B(_13079_),
    .Y(_13324_));
 AO21x1_ASAP7_75t_R _21577_ (.A1(net6204),
    .A2(_12904_),
    .B(net6207),
    .Y(_13325_));
 AOI21x1_ASAP7_75t_R _21578_ (.A1(net6204),
    .A2(net5499),
    .B(_13325_),
    .Y(_13326_));
 AO21x1_ASAP7_75t_R _21579_ (.A1(_13146_),
    .A2(_13242_),
    .B(net6211),
    .Y(_13327_));
 AND3x1_ASAP7_75t_R _21580_ (.A(net5848),
    .B(_13135_),
    .C(net6207),
    .Y(_13328_));
 AOI22x1_ASAP7_75t_R _21581_ (.A1(_13324_),
    .A2(_13326_),
    .B1(_13327_),
    .B2(_13328_),
    .Y(_13329_));
 AOI21x1_ASAP7_75t_R _21582_ (.A1(_13323_),
    .A2(_13329_),
    .B(net6200),
    .Y(_13330_));
 OAI21x1_ASAP7_75t_R _21583_ (.A1(net5858),
    .A2(net5496),
    .B(net6214),
    .Y(_13331_));
 OA21x2_ASAP7_75t_R _21584_ (.A1(_13331_),
    .A2(_13051_),
    .B(net6207),
    .Y(_13332_));
 INVx1_ASAP7_75t_R _21585_ (.A(_13118_),
    .Y(_13333_));
 AND3x1_ASAP7_75t_R _21586_ (.A(net5493),
    .B(net5851),
    .C(net4933),
    .Y(_13334_));
 AOI22x1_ASAP7_75t_R _21587_ (.A1(_13332_),
    .A2(_13333_),
    .B1(_13334_),
    .B2(_12989_),
    .Y(_13335_));
 NAND2x1_ASAP7_75t_R _21588_ (.A(_12971_),
    .B(_13236_),
    .Y(_13336_));
 AO21x1_ASAP7_75t_R _21589_ (.A1(_13160_),
    .A2(net5492),
    .B(net6214),
    .Y(_13337_));
 AOI21x1_ASAP7_75t_R _21590_ (.A1(_13336_),
    .A2(_13337_),
    .B(net6207),
    .Y(_13338_));
 INVx1_ASAP7_75t_R _21591_ (.A(_13237_),
    .Y(_13339_));
 NOR2x1_ASAP7_75t_R _21592_ (.A(_13339_),
    .B(_13120_),
    .Y(_13340_));
 OAI21x1_ASAP7_75t_R _21593_ (.A1(_13338_),
    .A2(_13340_),
    .B(net5848),
    .Y(_13341_));
 AOI21x1_ASAP7_75t_R _21594_ (.A1(_13335_),
    .A2(_13341_),
    .B(net6200),
    .Y(_13342_));
 OAI21x1_ASAP7_75t_R _21595_ (.A1(net5861),
    .A2(net5503),
    .B(net6213),
    .Y(_13343_));
 INVx1_ASAP7_75t_R _21596_ (.A(_13343_),
    .Y(_13344_));
 OAI21x1_ASAP7_75t_R _21597_ (.A1(net4689),
    .A2(_13173_),
    .B(net5856),
    .Y(_13345_));
 AOI21x1_ASAP7_75t_R _21598_ (.A1(_13286_),
    .A2(_13344_),
    .B(_13345_),
    .Y(_13346_));
 AOI21x1_ASAP7_75t_R _21599_ (.A1(net5864),
    .A2(net5862),
    .B(_12904_),
    .Y(_13347_));
 OAI21x1_ASAP7_75t_R _21600_ (.A1(net6202),
    .A2(_13347_),
    .B(net6207),
    .Y(_13348_));
 OAI21x1_ASAP7_75t_R _21601_ (.A1(_13348_),
    .A2(_13125_),
    .B(net5848),
    .Y(_13349_));
 NOR2x1_ASAP7_75t_R _21602_ (.A(_13346_),
    .B(_13349_),
    .Y(_13350_));
 OAI21x1_ASAP7_75t_R _21603_ (.A1(_13095_),
    .A2(net4578),
    .B(net6207),
    .Y(_13351_));
 NOR2x1_ASAP7_75t_R _21604_ (.A(_12989_),
    .B(_12991_),
    .Y(_13352_));
 NOR2x1_ASAP7_75t_R _21605_ (.A(_13351_),
    .B(_13352_),
    .Y(_13353_));
 AO21x1_ASAP7_75t_R _21606_ (.A1(_12924_),
    .A2(net6211),
    .B(net4934),
    .Y(_13354_));
 INVx1_ASAP7_75t_R _21607_ (.A(_13129_),
    .Y(_13355_));
 OAI21x1_ASAP7_75t_R _21608_ (.A1(_13354_),
    .A2(_13355_),
    .B(net5495),
    .Y(_13356_));
 OAI21x1_ASAP7_75t_R _21609_ (.A1(_13353_),
    .A2(_13356_),
    .B(net6200),
    .Y(_13357_));
 OAI21x1_ASAP7_75t_R _21610_ (.A1(_13350_),
    .A2(_13357_),
    .B(_13076_),
    .Y(_13358_));
 OAI22x1_ASAP7_75t_R _21611_ (.A1(_13317_),
    .A2(_13330_),
    .B1(_13342_),
    .B2(_13358_),
    .Y(_00060_));
 OA21x2_ASAP7_75t_R _21612_ (.A1(net5864),
    .A2(net6203),
    .B(net6207),
    .Y(_13359_));
 AND2x2_ASAP7_75t_R _21613_ (.A(_13337_),
    .B(_13359_),
    .Y(_13360_));
 NAND2x1_ASAP7_75t_R _21614_ (.A(net6213),
    .B(_12981_),
    .Y(_13361_));
 INVx1_ASAP7_75t_R _21615_ (.A(_13361_),
    .Y(_13362_));
 AO21x1_ASAP7_75t_R _21616_ (.A1(_13043_),
    .A2(net5490),
    .B(net6207),
    .Y(_13363_));
 AOI21x1_ASAP7_75t_R _21617_ (.A1(net5504),
    .A2(_13362_),
    .B(_13363_),
    .Y(_13364_));
 OAI21x1_ASAP7_75t_R _21618_ (.A1(_13360_),
    .A2(_13364_),
    .B(net5493),
    .Y(_13365_));
 NOR2x1_ASAP7_75t_R _21619_ (.A(net5069),
    .B(net5857),
    .Y(_13366_));
 OAI21x1_ASAP7_75t_R _21620_ (.A1(net4929),
    .A2(_13127_),
    .B(net6204),
    .Y(_13367_));
 OA21x2_ASAP7_75t_R _21621_ (.A1(_12925_),
    .A2(net6204),
    .B(net5851),
    .Y(_13368_));
 AOI21x1_ASAP7_75t_R _21622_ (.A1(_13367_),
    .A2(_13368_),
    .B(net5493),
    .Y(_13369_));
 AO21x1_ASAP7_75t_R _21623_ (.A1(_13056_),
    .A2(_12971_),
    .B(_13261_),
    .Y(_13370_));
 NAND2x1_ASAP7_75t_R _21624_ (.A(net6207),
    .B(_13370_),
    .Y(_13371_));
 AOI21x1_ASAP7_75t_R _21625_ (.A1(_13369_),
    .A2(_13371_),
    .B(net5850),
    .Y(_13372_));
 NAND2x1_ASAP7_75t_R _21626_ (.A(_13365_),
    .B(_13372_),
    .Y(_13373_));
 NOR2x1_ASAP7_75t_R _21627_ (.A(net6207),
    .B(_13140_),
    .Y(_13374_));
 OAI21x1_ASAP7_75t_R _21628_ (.A1(net6205),
    .A2(_13114_),
    .B(_13374_),
    .Y(_13375_));
 OA21x2_ASAP7_75t_R _21629_ (.A1(_13135_),
    .A2(net5863),
    .B(net6207),
    .Y(_13376_));
 AOI21x1_ASAP7_75t_R _21630_ (.A1(_13265_),
    .A2(_13376_),
    .B(net5494),
    .Y(_13377_));
 AOI21x1_ASAP7_75t_R _21631_ (.A1(_13375_),
    .A2(_13377_),
    .B(net6200),
    .Y(_13378_));
 INVx1_ASAP7_75t_R _21632_ (.A(net4937),
    .Y(_13379_));
 AOI21x1_ASAP7_75t_R _21633_ (.A1(net4687),
    .A2(_13203_),
    .B(net6207),
    .Y(_13380_));
 AND2x2_ASAP7_75t_R _21634_ (.A(_12988_),
    .B(net6202),
    .Y(_13381_));
 OAI21x1_ASAP7_75t_R _21635_ (.A1(net5860),
    .A2(net5503),
    .B(_13381_),
    .Y(_13382_));
 AOI21x1_ASAP7_75t_R _21636_ (.A1(_13380_),
    .A2(_13382_),
    .B(net5848),
    .Y(_13383_));
 AO21x1_ASAP7_75t_R _21637_ (.A1(_13155_),
    .A2(_13242_),
    .B(net6202),
    .Y(_13384_));
 NAND2x1_ASAP7_75t_R _21638_ (.A(_13384_),
    .B(_13064_),
    .Y(_13385_));
 NAND2x1_ASAP7_75t_R _21639_ (.A(_13383_),
    .B(_13385_),
    .Y(_13386_));
 AOI21x1_ASAP7_75t_R _21640_ (.A1(_13378_),
    .A2(_13386_),
    .B(net6199),
    .Y(_13387_));
 NAND2x1_ASAP7_75t_R _21641_ (.A(_13387_),
    .B(_13373_),
    .Y(_13388_));
 AOI211x1_ASAP7_75t_R _21642_ (.A1(net6201),
    .A2(_13184_),
    .B(_12942_),
    .C(net5189),
    .Y(_13389_));
 AO21x1_ASAP7_75t_R _21643_ (.A1(_13090_),
    .A2(_13089_),
    .B(_13172_),
    .Y(_13390_));
 OA21x2_ASAP7_75t_R _21644_ (.A1(_12981_),
    .A2(net6205),
    .B(net5853),
    .Y(_13391_));
 AO21x1_ASAP7_75t_R _21645_ (.A1(_13390_),
    .A2(_13391_),
    .B(net5494),
    .Y(_13392_));
 AND2x2_ASAP7_75t_R _21646_ (.A(_13225_),
    .B(net6207),
    .Y(_13393_));
 AOI21x1_ASAP7_75t_R _21647_ (.A1(_13393_),
    .A2(_13018_),
    .B(net5848),
    .Y(_13394_));
 OAI21x1_ASAP7_75t_R _21648_ (.A1(net4764),
    .A2(_13046_),
    .B(net6210),
    .Y(_13395_));
 AOI21x1_ASAP7_75t_R _21649_ (.A1(net5488),
    .A2(_13381_),
    .B(net6207),
    .Y(_13396_));
 NAND2x1_ASAP7_75t_R _21650_ (.A(_13395_),
    .B(_13396_),
    .Y(_13397_));
 AOI21x1_ASAP7_75t_R _21651_ (.A1(_13394_),
    .A2(_13397_),
    .B(net6200),
    .Y(_13398_));
 OAI21x1_ASAP7_75t_R _21652_ (.A1(_13389_),
    .A2(_13392_),
    .B(_13398_),
    .Y(_13399_));
 AO21x1_ASAP7_75t_R _21653_ (.A1(net6215),
    .A2(net6216),
    .B(_13379_),
    .Y(_13400_));
 AOI21x1_ASAP7_75t_R _21654_ (.A1(net6211),
    .A2(_13400_),
    .B(net5856),
    .Y(_13401_));
 OAI21x1_ASAP7_75t_R _21655_ (.A1(_13111_),
    .A2(net5185),
    .B(_13401_),
    .Y(_13402_));
 NAND2x1_ASAP7_75t_R _21656_ (.A(net6211),
    .B(net4931),
    .Y(_13403_));
 AOI21x1_ASAP7_75t_R _21657_ (.A1(_13403_),
    .A2(_13129_),
    .B(net5848),
    .Y(_13404_));
 AOI21x1_ASAP7_75t_R _21658_ (.A1(_13402_),
    .A2(_13404_),
    .B(net5849),
    .Y(_13405_));
 AO21x1_ASAP7_75t_R _21659_ (.A1(_12981_),
    .A2(_13022_),
    .B(net6205),
    .Y(_13406_));
 AOI21x1_ASAP7_75t_R _21660_ (.A1(net4931),
    .A2(net4579),
    .B(net6207),
    .Y(_13407_));
 AO21x1_ASAP7_75t_R _21661_ (.A1(net5068),
    .A2(net6211),
    .B(net5853),
    .Y(_13408_));
 OAI21x1_ASAP7_75t_R _21662_ (.A1(_13408_),
    .A2(_13091_),
    .B(net5848),
    .Y(_13409_));
 AO21x1_ASAP7_75t_R _21663_ (.A1(_13406_),
    .A2(_13407_),
    .B(_13409_),
    .Y(_13410_));
 AOI21x1_ASAP7_75t_R _21664_ (.A1(_13405_),
    .A2(_13410_),
    .B(_13076_),
    .Y(_13411_));
 NAND2x1_ASAP7_75t_R _21665_ (.A(_13399_),
    .B(_13411_),
    .Y(_13412_));
 NAND2x1_ASAP7_75t_R _21666_ (.A(_13412_),
    .B(_13388_),
    .Y(_00061_));
 OAI21x1_ASAP7_75t_R _21667_ (.A1(net6213),
    .A2(_12981_),
    .B(net5852),
    .Y(_13413_));
 OA21x2_ASAP7_75t_R _21668_ (.A1(_13184_),
    .A2(net5496),
    .B(net6212),
    .Y(_13414_));
 OAI21x1_ASAP7_75t_R _21669_ (.A1(_13413_),
    .A2(_13414_),
    .B(net5848),
    .Y(_13415_));
 AO21x1_ASAP7_75t_R _21670_ (.A1(_13147_),
    .A2(_13400_),
    .B(net5856),
    .Y(_13416_));
 AOI21x1_ASAP7_75t_R _21671_ (.A1(net5505),
    .A2(_13344_),
    .B(_13416_),
    .Y(_13417_));
 OAI21x1_ASAP7_75t_R _21672_ (.A1(_13415_),
    .A2(_13417_),
    .B(net6200),
    .Y(_13418_));
 AO21x1_ASAP7_75t_R _21673_ (.A1(net4577),
    .A2(net6206),
    .B(net6207),
    .Y(_13419_));
 AO21x1_ASAP7_75t_R _21674_ (.A1(net5185),
    .A2(_13221_),
    .B(_13419_),
    .Y(_13420_));
 OA21x2_ASAP7_75t_R _21675_ (.A1(net4577),
    .A2(net4929),
    .B(net6206),
    .Y(_13421_));
 AOI21x1_ASAP7_75t_R _21676_ (.A1(_13114_),
    .A2(_13168_),
    .B(net6206),
    .Y(_13422_));
 OAI21x1_ASAP7_75t_R _21677_ (.A1(_13421_),
    .A2(_13422_),
    .B(net6207),
    .Y(_13423_));
 AOI21x1_ASAP7_75t_R _21678_ (.A1(_13420_),
    .A2(_13423_),
    .B(net5848),
    .Y(_13424_));
 OAI21x1_ASAP7_75t_R _21679_ (.A1(_13418_),
    .A2(_13424_),
    .B(_13076_),
    .Y(_13425_));
 AO21x1_ASAP7_75t_R _21680_ (.A1(_13146_),
    .A2(_13250_),
    .B(net6211),
    .Y(_13426_));
 AO21x1_ASAP7_75t_R _21681_ (.A1(_12879_),
    .A2(_13246_),
    .B(net6201),
    .Y(_13427_));
 AO21x1_ASAP7_75t_R _21682_ (.A1(_13426_),
    .A2(_13427_),
    .B(net6207),
    .Y(_13428_));
 NOR2x1_ASAP7_75t_R _21683_ (.A(net6201),
    .B(_13020_),
    .Y(_13429_));
 OAI21x1_ASAP7_75t_R _21684_ (.A1(_13197_),
    .A2(_13179_),
    .B(net6201),
    .Y(_13430_));
 NAND2x1_ASAP7_75t_R _21685_ (.A(_13255_),
    .B(_13430_),
    .Y(_13431_));
 OAI21x1_ASAP7_75t_R _21686_ (.A1(_13429_),
    .A2(_13431_),
    .B(net6207),
    .Y(_13432_));
 AOI21x1_ASAP7_75t_R _21687_ (.A1(_13428_),
    .A2(_13432_),
    .B(net5495),
    .Y(_13433_));
 OA21x2_ASAP7_75t_R _21688_ (.A1(net4929),
    .A2(net4934),
    .B(net6212),
    .Y(_13434_));
 NOR2x1_ASAP7_75t_R _21689_ (.A(_13325_),
    .B(_13434_),
    .Y(_13435_));
 AO21x1_ASAP7_75t_R _21690_ (.A1(_13160_),
    .A2(net5491),
    .B(net6202),
    .Y(_13436_));
 AND2x2_ASAP7_75t_R _21691_ (.A(_01137_),
    .B(_01143_),
    .Y(_13437_));
 OA21x2_ASAP7_75t_R _21692_ (.A1(net6211),
    .A2(_13437_),
    .B(net6207),
    .Y(_13438_));
 AO21x1_ASAP7_75t_R _21693_ (.A1(_13436_),
    .A2(_13438_),
    .B(net5848),
    .Y(_13439_));
 OAI21x1_ASAP7_75t_R _21694_ (.A1(_13435_),
    .A2(_13439_),
    .B(net5849),
    .Y(_13440_));
 NOR2x1_ASAP7_75t_R _21695_ (.A(_13433_),
    .B(_13440_),
    .Y(_13441_));
 AO21x1_ASAP7_75t_R _21696_ (.A1(_13305_),
    .A2(_13110_),
    .B(net6207),
    .Y(_13442_));
 AO21x1_ASAP7_75t_R _21697_ (.A1(net6217),
    .A2(net6218),
    .B(_13139_),
    .Y(_13443_));
 INVx1_ASAP7_75t_R _21698_ (.A(_13443_),
    .Y(_13444_));
 OAI21x1_ASAP7_75t_R _21699_ (.A1(_13444_),
    .A2(_12991_),
    .B(net6212),
    .Y(_13445_));
 AOI21x1_ASAP7_75t_R _21700_ (.A1(net6207),
    .A2(_13445_),
    .B(net5849),
    .Y(_13446_));
 NAND2x1_ASAP7_75t_R _21701_ (.A(_13442_),
    .B(_13446_),
    .Y(_13447_));
 AO21x1_ASAP7_75t_R _21702_ (.A1(net6211),
    .A2(_13246_),
    .B(net4580),
    .Y(_13448_));
 AND2x2_ASAP7_75t_R _21703_ (.A(_13448_),
    .B(_13376_),
    .Y(_13449_));
 NAND2x1_ASAP7_75t_R _21704_ (.A(net5851),
    .B(_13331_),
    .Y(_13450_));
 NOR2x1_ASAP7_75t_R _21705_ (.A(_13051_),
    .B(net5185),
    .Y(_13451_));
 NOR2x1_ASAP7_75t_R _21706_ (.A(_13450_),
    .B(_13451_),
    .Y(_13452_));
 OAI21x1_ASAP7_75t_R _21707_ (.A1(_13449_),
    .A2(_13452_),
    .B(net5849),
    .Y(_13453_));
 AOI21x1_ASAP7_75t_R _21708_ (.A1(_13447_),
    .A2(_13453_),
    .B(net5493),
    .Y(_13454_));
 AO21x1_ASAP7_75t_R _21709_ (.A1(_01138_),
    .A2(net6212),
    .B(_12916_),
    .Y(_13455_));
 AOI21x1_ASAP7_75t_R _21710_ (.A1(_13160_),
    .A2(_13381_),
    .B(_13455_),
    .Y(_13456_));
 NOR2x1_ASAP7_75t_R _21711_ (.A(net4764),
    .B(_13403_),
    .Y(_13457_));
 AO21x1_ASAP7_75t_R _21712_ (.A1(_13013_),
    .A2(net6204),
    .B(net6207),
    .Y(_13458_));
 OAI21x1_ASAP7_75t_R _21713_ (.A1(_13457_),
    .A2(_13458_),
    .B(net6200),
    .Y(_13459_));
 OAI21x1_ASAP7_75t_R _21714_ (.A1(_13456_),
    .A2(_13459_),
    .B(net5493),
    .Y(_13460_));
 OAI21x1_ASAP7_75t_R _21715_ (.A1(net6204),
    .A2(net5489),
    .B(_13095_),
    .Y(_13461_));
 AOI21x1_ASAP7_75t_R _21716_ (.A1(net5505),
    .A2(_13461_),
    .B(net6207),
    .Y(_13462_));
 INVx1_ASAP7_75t_R _21717_ (.A(net5501),
    .Y(_13463_));
 AO21x1_ASAP7_75t_R _21718_ (.A1(_13295_),
    .A2(_13463_),
    .B(net6200),
    .Y(_13464_));
 NOR2x1_ASAP7_75t_R _21719_ (.A(_13462_),
    .B(_13464_),
    .Y(_13465_));
 OAI21x1_ASAP7_75t_R _21720_ (.A1(_13460_),
    .A2(_13465_),
    .B(net6199),
    .Y(_13466_));
 OAI22x1_ASAP7_75t_R _21721_ (.A1(_13425_),
    .A2(_13441_),
    .B1(_13454_),
    .B2(_13466_),
    .Y(_00062_));
 NAND2x1_ASAP7_75t_R _21722_ (.A(_13430_),
    .B(_13226_),
    .Y(_13467_));
 AOI21x1_ASAP7_75t_R _21723_ (.A1(_13070_),
    .A2(net4477),
    .B(net6207),
    .Y(_13468_));
 AOI21x1_ASAP7_75t_R _21724_ (.A1(_13244_),
    .A2(_13468_),
    .B(net5495),
    .Y(_13469_));
 OAI21x1_ASAP7_75t_R _21725_ (.A1(net5854),
    .A2(_13467_),
    .B(_13469_),
    .Y(_13470_));
 AOI21x1_ASAP7_75t_R _21726_ (.A1(net4524),
    .A2(_13020_),
    .B(net6201),
    .Y(_13471_));
 INVx1_ASAP7_75t_R _21727_ (.A(net5502),
    .Y(_13472_));
 OAI21x1_ASAP7_75t_R _21728_ (.A1(_13472_),
    .A2(_12991_),
    .B(net5856),
    .Y(_13473_));
 AOI21x1_ASAP7_75t_R _21729_ (.A1(net6202),
    .A2(_13070_),
    .B(_12916_),
    .Y(_13474_));
 AOI21x1_ASAP7_75t_R _21730_ (.A1(_13474_),
    .A2(_13305_),
    .B(net5848),
    .Y(_13475_));
 OAI21x1_ASAP7_75t_R _21731_ (.A1(_13471_),
    .A2(_13473_),
    .B(_13475_),
    .Y(_13476_));
 AOI21x1_ASAP7_75t_R _21732_ (.A1(_13470_),
    .A2(_13476_),
    .B(net6200),
    .Y(_13477_));
 OAI21x1_ASAP7_75t_R _21733_ (.A1(_13051_),
    .A2(_13127_),
    .B(net6213),
    .Y(_13478_));
 AOI21x1_ASAP7_75t_R _21734_ (.A1(net4475),
    .A2(_13478_),
    .B(net5852),
    .Y(_13479_));
 OAI21x1_ASAP7_75t_R _21735_ (.A1(net5858),
    .A2(net5490),
    .B(net4579),
    .Y(_13480_));
 AOI21x1_ASAP7_75t_R _21736_ (.A1(_13343_),
    .A2(_13480_),
    .B(net6207),
    .Y(_13481_));
 OAI21x1_ASAP7_75t_R _21737_ (.A1(_13479_),
    .A2(_13481_),
    .B(net5848),
    .Y(_13482_));
 OAI21x1_ASAP7_75t_R _21738_ (.A1(net5858),
    .A2(net5492),
    .B(net6204),
    .Y(_13483_));
 OAI21x1_ASAP7_75t_R _21739_ (.A1(_13127_),
    .A2(_13483_),
    .B(_13237_),
    .Y(_13484_));
 OAI21x1_ASAP7_75t_R _21740_ (.A1(_13051_),
    .A2(_13331_),
    .B(_13089_),
    .Y(_13485_));
 AOI21x1_ASAP7_75t_R _21741_ (.A1(net5851),
    .A2(_13485_),
    .B(net5848),
    .Y(_13486_));
 NAND2x1_ASAP7_75t_R _21742_ (.A(_13484_),
    .B(_13486_),
    .Y(_13487_));
 AOI21x1_ASAP7_75t_R _21743_ (.A1(_13482_),
    .A2(_13487_),
    .B(net5850),
    .Y(_13488_));
 OAI21x1_ASAP7_75t_R _21744_ (.A1(_13477_),
    .A2(_13488_),
    .B(net6199),
    .Y(_13489_));
 NOR2x1_ASAP7_75t_R _21745_ (.A(net6207),
    .B(net5501),
    .Y(_13490_));
 OAI21x1_ASAP7_75t_R _21746_ (.A1(net6214),
    .A2(_12979_),
    .B(_13490_),
    .Y(_13491_));
 NAND2x1_ASAP7_75t_R _21747_ (.A(net6203),
    .B(net4929),
    .Y(_13492_));
 OA21x2_ASAP7_75t_R _21748_ (.A1(_13300_),
    .A2(net6203),
    .B(net6207),
    .Y(_13493_));
 AOI21x1_ASAP7_75t_R _21749_ (.A1(_13492_),
    .A2(_13493_),
    .B(net5848),
    .Y(_13494_));
 OAI21x1_ASAP7_75t_R _21750_ (.A1(net4930),
    .A2(_13491_),
    .B(_13494_),
    .Y(_13495_));
 NAND2x1p5_ASAP7_75t_R _21751_ (.A(net4476),
    .B(_13022_),
    .Y(_13496_));
 NAND2x1_ASAP7_75t_R _21752_ (.A(net5488),
    .B(net5502),
    .Y(_13497_));
 AOI21x1_ASAP7_75t_R _21753_ (.A1(_13496_),
    .A2(_13497_),
    .B(net6207),
    .Y(_13498_));
 NOR2x1_ASAP7_75t_R _21754_ (.A(net4934),
    .B(net4578),
    .Y(_13499_));
 AO21x1_ASAP7_75t_R _21755_ (.A1(_01143_),
    .A2(net6212),
    .B(_12916_),
    .Y(_13500_));
 AOI21x1_ASAP7_75t_R _21756_ (.A1(net6202),
    .A2(_13499_),
    .B(_13500_),
    .Y(_13501_));
 OAI21x1_ASAP7_75t_R _21757_ (.A1(_13498_),
    .A2(_13501_),
    .B(net5848),
    .Y(_13502_));
 AOI21x1_ASAP7_75t_R _21758_ (.A1(_13502_),
    .A2(_13495_),
    .B(net5849),
    .Y(_13503_));
 AO21x1_ASAP7_75t_R _21759_ (.A1(_13139_),
    .A2(net6203),
    .B(net6207),
    .Y(_13504_));
 AO21x1_ASAP7_75t_R _21760_ (.A1(_12990_),
    .A2(_13281_),
    .B(_13504_),
    .Y(_13505_));
 NAND2x1_ASAP7_75t_R _21761_ (.A(net6212),
    .B(net5498),
    .Y(_13506_));
 NAND2x1_ASAP7_75t_R _21762_ (.A(net6207),
    .B(net4524),
    .Y(_13507_));
 AOI21x1_ASAP7_75t_R _21763_ (.A1(net6203),
    .A2(net4929),
    .B(_13507_),
    .Y(_13508_));
 AOI21x1_ASAP7_75t_R _21764_ (.A1(_13506_),
    .A2(_13508_),
    .B(net5493),
    .Y(_13509_));
 NAND2x1_ASAP7_75t_R _21765_ (.A(_13505_),
    .B(_13509_),
    .Y(_13510_));
 NOR2x1_ASAP7_75t_R _21766_ (.A(net4577),
    .B(_13361_),
    .Y(_13511_));
 NAND2x1_ASAP7_75t_R _21767_ (.A(net6204),
    .B(net4524),
    .Y(_13512_));
 AOI21x1_ASAP7_75t_R _21768_ (.A1(net5861),
    .A2(net5490),
    .B(_13512_),
    .Y(_13513_));
 OAI21x1_ASAP7_75t_R _21769_ (.A1(_13511_),
    .A2(_13513_),
    .B(net6207),
    .Y(_13514_));
 NOR2x1_ASAP7_75t_R _21770_ (.A(net5858),
    .B(_13089_),
    .Y(_13515_));
 NOR2x1_ASAP7_75t_R _21771_ (.A(_13515_),
    .B(_13260_),
    .Y(_13516_));
 AOI21x1_ASAP7_75t_R _21772_ (.A1(_13490_),
    .A2(_13516_),
    .B(net5848),
    .Y(_13517_));
 NAND2x1_ASAP7_75t_R _21773_ (.A(_13514_),
    .B(_13517_),
    .Y(_13518_));
 AOI21x1_ASAP7_75t_R _21774_ (.A1(_13510_),
    .A2(_13518_),
    .B(net6200),
    .Y(_13519_));
 OAI21x1_ASAP7_75t_R _21775_ (.A1(_13503_),
    .A2(_13519_),
    .B(_13076_),
    .Y(_13520_));
 NAND2x1_ASAP7_75t_R _21776_ (.A(_13520_),
    .B(_13489_),
    .Y(_00063_));
 INVx1_ASAP7_75t_R _21777_ (.A(net6649),
    .Y(_13521_));
 XOR2x2_ASAP7_75t_R _21778_ (.A(_10682_),
    .B(_13521_),
    .Y(_13522_));
 XNOR2x2_ASAP7_75t_R _21779_ (.A(_00646_),
    .B(_00639_),
    .Y(_13523_));
 XOR2x2_ASAP7_75t_R _21780_ (.A(_00672_),
    .B(_00640_),
    .Y(_13524_));
 XOR2x2_ASAP7_75t_R _21781_ (.A(_13523_),
    .B(_13524_),
    .Y(_13525_));
 NOR2x1p5_ASAP7_75t_R _21782_ (.A(_13522_),
    .B(_13525_),
    .Y(_13526_));
 XOR2x2_ASAP7_75t_R _21783_ (.A(_10682_),
    .B(net6649),
    .Y(_13527_));
 XOR2x2_ASAP7_75t_R _21784_ (.A(_00646_),
    .B(_00639_),
    .Y(_13528_));
 XOR2x2_ASAP7_75t_R _21785_ (.A(_13528_),
    .B(_13524_),
    .Y(_13529_));
 OAI21x1_ASAP7_75t_R _21786_ (.A1(_13527_),
    .A2(_13529_),
    .B(net6673),
    .Y(_13530_));
 NAND2x1_ASAP7_75t_R _21787_ (.A(_00456_),
    .B(_10676_),
    .Y(_13531_));
 OAI21x1_ASAP7_75t_R _21788_ (.A1(_13530_),
    .A2(_13526_),
    .B(_13531_),
    .Y(_13532_));
 XOR2x2_ASAP7_75t_R _21789_ (.A(net6359),
    .B(net6532),
    .Y(_13533_));
 XOR2x2_ASAP7_75t_R _21791_ (.A(_00575_),
    .B(net6618),
    .Y(_13534_));
 NAND2x1_ASAP7_75t_R _21792_ (.A(_10696_),
    .B(_13534_),
    .Y(_13535_));
 XNOR2x2_ASAP7_75t_R _21793_ (.A(_00575_),
    .B(net6618),
    .Y(_13536_));
 NAND2x1_ASAP7_75t_R _21794_ (.A(net6567),
    .B(_13536_),
    .Y(_13537_));
 AOI21x1_ASAP7_75t_R _21795_ (.A1(_13535_),
    .A2(_13537_),
    .B(_13523_),
    .Y(_13538_));
 XOR2x2_ASAP7_75t_R _21796_ (.A(net6618),
    .B(net6569),
    .Y(_13539_));
 NAND2x1_ASAP7_75t_R _21797_ (.A(net6651),
    .B(_13539_),
    .Y(_13540_));
 INVx1_ASAP7_75t_R _21798_ (.A(net6651),
    .Y(_13541_));
 XNOR2x2_ASAP7_75t_R _21799_ (.A(net6618),
    .B(net6569),
    .Y(_13542_));
 NAND2x1_ASAP7_75t_R _21800_ (.A(_13541_),
    .B(_13542_),
    .Y(_13543_));
 AOI21x1_ASAP7_75t_R _21801_ (.A1(_13540_),
    .A2(_13543_),
    .B(_13528_),
    .Y(_13544_));
 OAI21x1_ASAP7_75t_R _21803_ (.A1(_13538_),
    .A2(_13544_),
    .B(net6673),
    .Y(_13546_));
 INVx1_ASAP7_75t_R _21804_ (.A(net6533),
    .Y(_13547_));
 NOR2x1_ASAP7_75t_R _21805_ (.A(net6664),
    .B(_00457_),
    .Y(_13548_));
 INVx1_ASAP7_75t_R _21806_ (.A(_13548_),
    .Y(_13549_));
 NAND3x1_ASAP7_75t_R _21807_ (.A(_13546_),
    .B(_13547_),
    .C(_13549_),
    .Y(_13550_));
 AO21x1_ASAP7_75t_R _21808_ (.A1(_13546_),
    .A2(_13549_),
    .B(_13547_),
    .Y(_13551_));
 NAND2x1_ASAP7_75t_R _21809_ (.A(_13550_),
    .B(_13551_),
    .Y(_01152_));
 OR2x2_ASAP7_75t_R _21810_ (.A(net6660),
    .B(_00458_),
    .Y(_13552_));
 INVx1_ASAP7_75t_R _21811_ (.A(_00577_),
    .Y(_13553_));
 NOR2x1_ASAP7_75t_R _21812_ (.A(_13553_),
    .B(_10725_),
    .Y(_13554_));
 NOR2x1_ASAP7_75t_R _21813_ (.A(net6646),
    .B(_10721_),
    .Y(_13555_));
 OAI21x1_ASAP7_75t_R _21814_ (.A1(_13554_),
    .A2(_13555_),
    .B(net6451),
    .Y(_13556_));
 INVx1_ASAP7_75t_R _21815_ (.A(_13556_),
    .Y(_13557_));
 NAND2x1_ASAP7_75t_R _21816_ (.A(_13553_),
    .B(_10725_),
    .Y(_13558_));
 INVx1_ASAP7_75t_R _21817_ (.A(net6451),
    .Y(_13559_));
 NOR2x1_ASAP7_75t_R _21818_ (.A(_00641_),
    .B(_00673_),
    .Y(_13560_));
 AND2x2_ASAP7_75t_R _21819_ (.A(_00641_),
    .B(_00673_),
    .Y(_13561_));
 OAI21x1_ASAP7_75t_R _21820_ (.A1(_13560_),
    .A2(_13561_),
    .B(net6646),
    .Y(_13562_));
 NAND3x1_ASAP7_75t_R _21821_ (.A(_13558_),
    .B(_13559_),
    .C(_13562_),
    .Y(_13563_));
 INVx1_ASAP7_75t_R _21822_ (.A(_13563_),
    .Y(_13564_));
 OAI21x1_ASAP7_75t_R _21823_ (.A1(_13557_),
    .A2(_13564_),
    .B(net6653),
    .Y(_13565_));
 INVx1_ASAP7_75t_R _21824_ (.A(net6531),
    .Y(_13566_));
 AOI21x1_ASAP7_75t_R _21825_ (.A1(_13552_),
    .A2(_13565_),
    .B(_13566_),
    .Y(_13567_));
 NAND2x1_ASAP7_75t_R _21826_ (.A(_00458_),
    .B(net6456),
    .Y(_13568_));
 NAND3x1_ASAP7_75t_R _21827_ (.A(_13563_),
    .B(net6653),
    .C(_13556_),
    .Y(_13569_));
 AOI21x1_ASAP7_75t_R _21828_ (.A1(_13568_),
    .A2(_13569_),
    .B(net6531),
    .Y(_13570_));
 NOR2x1_ASAP7_75t_R _21829_ (.A(_13567_),
    .B(_13570_),
    .Y(_13571_));
 INVx1_ASAP7_75t_R _21832_ (.A(_13546_),
    .Y(_13573_));
 OAI21x1_ASAP7_75t_R _21833_ (.A1(_13548_),
    .A2(_13573_),
    .B(_13547_),
    .Y(_13574_));
 NAND3x1_ASAP7_75t_R _21834_ (.A(_13546_),
    .B(net6533),
    .C(_13549_),
    .Y(_13575_));
 NAND2x1_ASAP7_75t_R _21835_ (.A(_13574_),
    .B(_13575_),
    .Y(_13576_));
 AOI21x1_ASAP7_75t_R _21838_ (.A1(_13552_),
    .A2(_13565_),
    .B(net6531),
    .Y(_13578_));
 AOI21x1_ASAP7_75t_R _21839_ (.A1(_13568_),
    .A2(_13569_),
    .B(_13566_),
    .Y(_13579_));
 NOR2x1_ASAP7_75t_R _21840_ (.A(_13578_),
    .B(_13579_),
    .Y(_13580_));
 XOR2x2_ASAP7_75t_R _21843_ (.A(_10761_),
    .B(net6645),
    .Y(_13582_));
 XOR2x2_ASAP7_75t_R _21844_ (.A(_00641_),
    .B(net6593),
    .Y(_13583_));
 XNOR2x2_ASAP7_75t_R _21845_ (.A(_13583_),
    .B(_10760_),
    .Y(_13584_));
 NOR2x1_ASAP7_75t_R _21846_ (.A(_13582_),
    .B(_13584_),
    .Y(_13585_));
 XNOR2x2_ASAP7_75t_R _21847_ (.A(net6645),
    .B(_10761_),
    .Y(_13586_));
 XOR2x2_ASAP7_75t_R _21848_ (.A(_10760_),
    .B(_13583_),
    .Y(_13587_));
 NOR2x1_ASAP7_75t_R _21849_ (.A(_13586_),
    .B(_13587_),
    .Y(_13588_));
 OAI21x1_ASAP7_75t_R _21850_ (.A1(_13585_),
    .A2(_13588_),
    .B(net6669),
    .Y(_13589_));
 INVx1_ASAP7_75t_R _21851_ (.A(net6530),
    .Y(_13590_));
 NOR2x1_ASAP7_75t_R _21852_ (.A(net6663),
    .B(_00559_),
    .Y(_13591_));
 INVx1_ASAP7_75t_R _21853_ (.A(_13591_),
    .Y(_13592_));
 NAND3x1_ASAP7_75t_R _21854_ (.A(_13589_),
    .B(_13590_),
    .C(_13592_),
    .Y(_13593_));
 AO21x1_ASAP7_75t_R _21855_ (.A1(_13589_),
    .A2(_13592_),
    .B(_13590_),
    .Y(_13594_));
 NAND2x1_ASAP7_75t_R _21856_ (.A(_13593_),
    .B(_13594_),
    .Y(_13595_));
 INVx1_ASAP7_75t_R _21858_ (.A(_01154_),
    .Y(_13597_));
 OAI21x1_ASAP7_75t_R _21859_ (.A1(net5845),
    .A2(net6196),
    .B(_13597_),
    .Y(_13598_));
 NOR2x1_ASAP7_75t_R _21860_ (.A(net6668),
    .B(_00558_),
    .Y(_13599_));
 XOR2x2_ASAP7_75t_R _21861_ (.A(_00579_),
    .B(_00643_),
    .Y(_13600_));
 XOR2x2_ASAP7_75t_R _21862_ (.A(_10775_),
    .B(_13600_),
    .Y(_13601_));
 XOR2x2_ASAP7_75t_R _21863_ (.A(net6595),
    .B(net6593),
    .Y(_13602_));
 XOR2x2_ASAP7_75t_R _21864_ (.A(_13602_),
    .B(net6562),
    .Y(_13603_));
 XOR2x2_ASAP7_75t_R _21865_ (.A(_13601_),
    .B(_13603_),
    .Y(_13604_));
 NOR2x1_ASAP7_75t_R _21866_ (.A(net6461),
    .B(_13604_),
    .Y(_13605_));
 INVx1_ASAP7_75t_R _21867_ (.A(_00850_),
    .Y(_13606_));
 OAI21x1_ASAP7_75t_R _21868_ (.A1(_13599_),
    .A2(_13605_),
    .B(_13606_),
    .Y(_13607_));
 AND2x2_ASAP7_75t_R _21869_ (.A(net6461),
    .B(_00558_),
    .Y(_13608_));
 XNOR2x2_ASAP7_75t_R _21870_ (.A(_13603_),
    .B(_13601_),
    .Y(_13609_));
 NOR2x1_ASAP7_75t_R _21871_ (.A(net6461),
    .B(_13609_),
    .Y(_13610_));
 OAI21x1_ASAP7_75t_R _21872_ (.A1(_13608_),
    .A2(_13610_),
    .B(_00850_),
    .Y(_13611_));
 NAND2x1_ASAP7_75t_R _21873_ (.A(_13607_),
    .B(_13611_),
    .Y(_13612_));
 INVx2_ASAP7_75t_R _21874_ (.A(_13612_),
    .Y(_13613_));
 OA21x2_ASAP7_75t_R _21875_ (.A1(net5839),
    .A2(net4928),
    .B(net5479),
    .Y(_13614_));
 INVx1_ASAP7_75t_R _21876_ (.A(_01151_),
    .Y(_13615_));
 OAI21x1_ASAP7_75t_R _21877_ (.A1(net5844),
    .A2(net6195),
    .B(_13615_),
    .Y(_13616_));
 NOR2x1_ASAP7_75t_R _21879_ (.A(_13616_),
    .B(net5840),
    .Y(_13618_));
 OAI21x1_ASAP7_75t_R _21880_ (.A1(net5845),
    .A2(net6196),
    .B(net4988),
    .Y(_13619_));
 NAND2x1_ASAP7_75t_R _21881_ (.A(_13619_),
    .B(_13595_),
    .Y(_13620_));
 INVx1_ASAP7_75t_R _21882_ (.A(_13620_),
    .Y(_13621_));
 NOR2x1_ASAP7_75t_R _21883_ (.A(net4522),
    .B(net4474),
    .Y(_13622_));
 XOR2x2_ASAP7_75t_R _21884_ (.A(_00645_),
    .B(_00677_),
    .Y(_13623_));
 XOR2x2_ASAP7_75t_R _21885_ (.A(_10802_),
    .B(_00581_),
    .Y(_13624_));
 XNOR2x2_ASAP7_75t_R _21886_ (.A(_13623_),
    .B(_13624_),
    .Y(_13625_));
 NOR2x1_ASAP7_75t_R _21887_ (.A(net6668),
    .B(_00556_),
    .Y(_13626_));
 AO21x1_ASAP7_75t_R _21888_ (.A1(_13625_),
    .A2(net6668),
    .B(_13626_),
    .Y(_13627_));
 XOR2x2_ASAP7_75t_R _21889_ (.A(_13627_),
    .B(_00852_),
    .Y(_13628_));
 AOI21x1_ASAP7_75t_R _21891_ (.A1(net4686),
    .A2(_13622_),
    .B(net6194),
    .Y(_13630_));
 OAI21x1_ASAP7_75t_R _21893_ (.A1(net4685),
    .A2(net5840),
    .B(net5834),
    .Y(_13632_));
 NAND2x1_ASAP7_75t_R _21894_ (.A(net5847),
    .B(net5487),
    .Y(_13633_));
 XNOR2x2_ASAP7_75t_R _21895_ (.A(_13532_),
    .B(net6532),
    .Y(_13634_));
 OAI21x1_ASAP7_75t_R _21896_ (.A1(net5483),
    .A2(net6193),
    .B(net5481),
    .Y(_13635_));
 INVx1_ASAP7_75t_R _21897_ (.A(_13589_),
    .Y(_13636_));
 OAI21x1_ASAP7_75t_R _21898_ (.A1(_13591_),
    .A2(_13636_),
    .B(_13590_),
    .Y(_13637_));
 NAND3x1_ASAP7_75t_R _21899_ (.A(_13589_),
    .B(net6530),
    .C(_13592_),
    .Y(_13638_));
 NAND2x1_ASAP7_75t_R _21900_ (.A(_13637_),
    .B(_13638_),
    .Y(_13639_));
 AOI21x1_ASAP7_75t_R _21902_ (.A1(_13633_),
    .A2(_13635_),
    .B(net5468),
    .Y(_13641_));
 OR2x2_ASAP7_75t_R _21903_ (.A(_13632_),
    .B(_13641_),
    .Y(_13642_));
 OAI21x1_ASAP7_75t_R _21905_ (.A1(net5846),
    .A2(net6193),
    .B(net5480),
    .Y(_13643_));
 AOI21x1_ASAP7_75t_R _21906_ (.A1(_13616_),
    .A2(_13643_),
    .B(net5839),
    .Y(_13644_));
 INVx1_ASAP7_75t_R _21907_ (.A(_13644_),
    .Y(_13645_));
 OAI21x1_ASAP7_75t_R _21910_ (.A1(net5845),
    .A2(net6196),
    .B(_01147_),
    .Y(_13648_));
 OAI21x1_ASAP7_75t_R _21911_ (.A1(net5483),
    .A2(net5480),
    .B(net4925),
    .Y(_13649_));
 INVx1_ASAP7_75t_R _21913_ (.A(net5065),
    .Y(_13651_));
 NAND2x1_ASAP7_75t_R _21914_ (.A(_13651_),
    .B(net5485),
    .Y(_13652_));
 OAI21x1_ASAP7_75t_R _21916_ (.A1(net5838),
    .A2(_13652_),
    .B(net5829),
    .Y(_13654_));
 AOI21x1_ASAP7_75t_R _21917_ (.A1(net5839),
    .A2(_13649_),
    .B(_13654_),
    .Y(_13655_));
 NOR2x1_ASAP7_75t_R _21919_ (.A(_01161_),
    .B(net5466),
    .Y(_13657_));
 INVx1_ASAP7_75t_R _21920_ (.A(_01148_),
    .Y(_13658_));
 OAI21x1_ASAP7_75t_R _21921_ (.A1(net5844),
    .A2(net6195),
    .B(_13658_),
    .Y(_13659_));
 OAI21x1_ASAP7_75t_R _21923_ (.A1(net4575),
    .A2(net5838),
    .B(net5478),
    .Y(_13661_));
 OAI21x1_ASAP7_75t_R _21925_ (.A1(_13657_),
    .A2(_13661_),
    .B(net6194),
    .Y(_13663_));
 AOI21x1_ASAP7_75t_R _21926_ (.A1(net4448),
    .A2(_13655_),
    .B(_13663_),
    .Y(_13664_));
 XNOR2x2_ASAP7_75t_R _21927_ (.A(_00580_),
    .B(_00611_),
    .Y(_13665_));
 INVx1_ASAP7_75t_R _21928_ (.A(_13665_),
    .Y(_13666_));
 XOR2x2_ASAP7_75t_R _21929_ (.A(_00643_),
    .B(net6594),
    .Y(_13667_));
 XOR2x2_ASAP7_75t_R _21930_ (.A(_13667_),
    .B(net6561),
    .Y(_13668_));
 NOR2x1_ASAP7_75t_R _21931_ (.A(_13666_),
    .B(_13668_),
    .Y(_13669_));
 XOR2x2_ASAP7_75t_R _21932_ (.A(_13667_),
    .B(_10803_),
    .Y(_13670_));
 NOR2x1_ASAP7_75t_R _21933_ (.A(_13665_),
    .B(_13670_),
    .Y(_13671_));
 OAI21x1_ASAP7_75t_R _21934_ (.A1(_13669_),
    .A2(_13671_),
    .B(net6666),
    .Y(_13672_));
 NOR2x1_ASAP7_75t_R _21935_ (.A(net6665),
    .B(_00557_),
    .Y(_13673_));
 INVx1_ASAP7_75t_R _21936_ (.A(_13673_),
    .Y(_13674_));
 NAND3x1_ASAP7_75t_R _21937_ (.A(_13672_),
    .B(_00851_),
    .C(_13674_),
    .Y(_13675_));
 AO21x1_ASAP7_75t_R _21938_ (.A1(_13672_),
    .A2(_13674_),
    .B(_00851_),
    .Y(_13676_));
 NAND2x1_ASAP7_75t_R _21939_ (.A(_13675_),
    .B(_13676_),
    .Y(_13677_));
 INVx1_ASAP7_75t_R _21940_ (.A(_13677_),
    .Y(_13678_));
 AOI211x1_ASAP7_75t_R _21943_ (.A1(_13630_),
    .A2(net4449),
    .B(_13664_),
    .C(net5463),
    .Y(_13681_));
 NOR2x1_ASAP7_75t_R _21944_ (.A(_01149_),
    .B(net5486),
    .Y(_13682_));
 AO21x1_ASAP7_75t_R _21947_ (.A1(net4924),
    .A2(net5470),
    .B(net5479),
    .Y(_13685_));
 NAND2x1_ASAP7_75t_R _21948_ (.A(net5483),
    .B(net6197),
    .Y(_13686_));
 INVx1_ASAP7_75t_R _21949_ (.A(_13686_),
    .Y(_13687_));
 OAI21x1_ASAP7_75t_R _21951_ (.A1(net5183),
    .A2(net5480),
    .B(net5840),
    .Y(_13689_));
 AOI21x1_ASAP7_75t_R _21952_ (.A1(net5480),
    .A2(_13687_),
    .B(_13689_),
    .Y(_13690_));
 NOR2x1_ASAP7_75t_R _21953_ (.A(_13685_),
    .B(_13690_),
    .Y(_13691_));
 NAND2x1_ASAP7_75t_R _21954_ (.A(net5293),
    .B(net5487),
    .Y(_13692_));
 AOI21x1_ASAP7_75t_R _21956_ (.A1(net5180),
    .A2(_13643_),
    .B(net5838),
    .Y(_13694_));
 AO21x1_ASAP7_75t_R _21958_ (.A1(net4924),
    .A2(net5838),
    .B(net5829),
    .Y(_13696_));
 OAI21x1_ASAP7_75t_R _21959_ (.A1(_13694_),
    .A2(_13696_),
    .B(net6194),
    .Y(_13697_));
 OAI21x1_ASAP7_75t_R _21960_ (.A1(_13691_),
    .A2(_13697_),
    .B(net5463),
    .Y(_13698_));
 AOI21x1_ASAP7_75t_R _21962_ (.A1(net5064),
    .A2(net5480),
    .B(net5466),
    .Y(_13700_));
 OAI21x1_ASAP7_75t_R _21963_ (.A1(net5844),
    .A2(net6195),
    .B(_01147_),
    .Y(_13701_));
 INVx1_ASAP7_75t_R _21964_ (.A(_13701_),
    .Y(_13702_));
 OA21x2_ASAP7_75t_R _21966_ (.A1(net4922),
    .A2(_13702_),
    .B(net5468),
    .Y(_13704_));
 OAI21x1_ASAP7_75t_R _21968_ (.A1(_13700_),
    .A2(_13704_),
    .B(net5478),
    .Y(_13706_));
 NAND2x1_ASAP7_75t_R _21969_ (.A(net5846),
    .B(net5480),
    .Y(_13707_));
 AOI21x1_ASAP7_75t_R _21972_ (.A1(_13707_),
    .A2(net5180),
    .B(net5466),
    .Y(_13710_));
 INVx2_ASAP7_75t_R _21973_ (.A(net4574),
    .Y(_13711_));
 NAND2x1_ASAP7_75t_R _21974_ (.A(net6197),
    .B(net5482),
    .Y(_13712_));
 NAND2x1_ASAP7_75t_R _21975_ (.A(net5471),
    .B(_13712_),
    .Y(_13713_));
 NOR2x1p5_ASAP7_75t_R _21976_ (.A(net4472),
    .B(_13713_),
    .Y(_13714_));
 OAI21x1_ASAP7_75t_R _21978_ (.A1(_13710_),
    .A2(_13714_),
    .B(net5834),
    .Y(_13716_));
 AOI21x1_ASAP7_75t_R _21979_ (.A1(_13706_),
    .A2(_13716_),
    .B(net6194),
    .Y(_13717_));
 XOR2x2_ASAP7_75t_R _21980_ (.A(_00645_),
    .B(net6593),
    .Y(_13718_));
 XOR2x2_ASAP7_75t_R _21981_ (.A(_13718_),
    .B(net6445),
    .Y(_13719_));
 XOR2x2_ASAP7_75t_R _21982_ (.A(net6644),
    .B(_00613_),
    .Y(_13720_));
 XOR2x2_ASAP7_75t_R _21983_ (.A(_13719_),
    .B(_13720_),
    .Y(_13721_));
 NOR2x1_ASAP7_75t_R _21984_ (.A(net6657),
    .B(_00555_),
    .Y(_13722_));
 AO21x1_ASAP7_75t_R _21985_ (.A1(_13721_),
    .A2(net6664),
    .B(_13722_),
    .Y(_13723_));
 XOR2x2_ASAP7_75t_R _21986_ (.A(_13723_),
    .B(_00853_),
    .Y(_13724_));
 INVx1_ASAP7_75t_R _21987_ (.A(_13724_),
    .Y(_13725_));
 OAI21x1_ASAP7_75t_R _21988_ (.A1(_13698_),
    .A2(_13717_),
    .B(_13725_),
    .Y(_13726_));
 NOR2x1_ASAP7_75t_R _21989_ (.A(net6197),
    .B(net5480),
    .Y(_13727_));
 OA21x2_ASAP7_75t_R _21990_ (.A1(net4922),
    .A2(_13727_),
    .B(net5468),
    .Y(_13728_));
 OAI21x1_ASAP7_75t_R _21992_ (.A1(net4926),
    .A2(_13728_),
    .B(net5833),
    .Y(_13730_));
 NOR2x1_ASAP7_75t_R _21993_ (.A(net5483),
    .B(net5482),
    .Y(_13731_));
 NOR2x1_ASAP7_75t_R _21995_ (.A(net5291),
    .B(net5486),
    .Y(_13733_));
 OA21x2_ASAP7_75t_R _21996_ (.A1(net5178),
    .A2(_13733_),
    .B(net5843),
    .Y(_13734_));
 NOR2x1_ASAP7_75t_R _21997_ (.A(net5481),
    .B(_13686_),
    .Y(_13735_));
 NAND2x1_ASAP7_75t_R _21998_ (.A(net6193),
    .B(net5482),
    .Y(_13736_));
 NAND2x1_ASAP7_75t_R _21999_ (.A(net5467),
    .B(_13736_),
    .Y(_13737_));
 NOR2x1_ASAP7_75t_R _22000_ (.A(net4920),
    .B(_13737_),
    .Y(_13738_));
 OAI21x1_ASAP7_75t_R _22002_ (.A1(_13734_),
    .A2(_13738_),
    .B(net5476),
    .Y(_13740_));
 AOI21x1_ASAP7_75t_R _22003_ (.A1(_13730_),
    .A2(_13740_),
    .B(net5464),
    .Y(_13741_));
 NAND2x1_ASAP7_75t_R _22004_ (.A(net5291),
    .B(net5486),
    .Y(_13742_));
 AND3x1_ASAP7_75t_R _22007_ (.A(_13742_),
    .B(net5843),
    .C(net4762),
    .Y(_13745_));
 NAND2x1_ASAP7_75t_R _22008_ (.A(net5483),
    .B(net5480),
    .Y(_13746_));
 NAND2x1_ASAP7_75t_R _22009_ (.A(net5475),
    .B(_13746_),
    .Y(_13747_));
 OAI21x1_ASAP7_75t_R _22011_ (.A1(_13687_),
    .A2(_13747_),
    .B(net5479),
    .Y(_13749_));
 NOR2x1_ASAP7_75t_R _22012_ (.A(_13745_),
    .B(_13749_),
    .Y(_13750_));
 NAND2x1_ASAP7_75t_R _22013_ (.A(net5483),
    .B(net5486),
    .Y(_13751_));
 AO21x1_ASAP7_75t_R _22015_ (.A1(_13751_),
    .A2(net5469),
    .B(net5479),
    .Y(_13753_));
 OAI21x1_ASAP7_75t_R _22016_ (.A1(net5845),
    .A2(net6196),
    .B(net4927),
    .Y(_13754_));
 AO21x1_ASAP7_75t_R _22017_ (.A1(net6197),
    .A2(net5483),
    .B(net5482),
    .Y(_13755_));
 AOI21x1_ASAP7_75t_R _22018_ (.A1(net4682),
    .A2(_13755_),
    .B(net5468),
    .Y(_13756_));
 OAI21x1_ASAP7_75t_R _22020_ (.A1(_13753_),
    .A2(_13756_),
    .B(net5465),
    .Y(_13758_));
 INVx1_ASAP7_75t_R _22021_ (.A(_13628_),
    .Y(_13759_));
 OAI21x1_ASAP7_75t_R _22023_ (.A1(_13750_),
    .A2(_13758_),
    .B(net5825),
    .Y(_13761_));
 OAI21x1_ASAP7_75t_R _22024_ (.A1(_13741_),
    .A2(_13761_),
    .B(net6192),
    .Y(_13762_));
 AO21x1_ASAP7_75t_R _22025_ (.A1(_13633_),
    .A2(_13686_),
    .B(net5840),
    .Y(_13763_));
 NAND2x1_ASAP7_75t_R _22026_ (.A(net5483),
    .B(net6193),
    .Y(_13764_));
 AOI21x1_ASAP7_75t_R _22027_ (.A1(net5177),
    .A2(_13707_),
    .B(net5466),
    .Y(_13765_));
 NOR2x1_ASAP7_75t_R _22028_ (.A(net5834),
    .B(_13765_),
    .Y(_13766_));
 NAND2x1_ASAP7_75t_R _22029_ (.A(_13763_),
    .B(_13766_),
    .Y(_13767_));
 INVx1_ASAP7_75t_R _22030_ (.A(_01153_),
    .Y(_13768_));
 OAI21x1_ASAP7_75t_R _22031_ (.A1(net5176),
    .A2(net5486),
    .B(net4921),
    .Y(_13769_));
 AOI21x1_ASAP7_75t_R _22032_ (.A1(net5835),
    .A2(_13769_),
    .B(net5477),
    .Y(_13770_));
 OAI21x1_ASAP7_75t_R _22033_ (.A1(net5483),
    .A2(net6193),
    .B(net5486),
    .Y(_13771_));
 OAI21x1_ASAP7_75t_R _22034_ (.A1(net5845),
    .A2(net6196),
    .B(_13658_),
    .Y(_13772_));
 AO21x1_ASAP7_75t_R _22035_ (.A1(_13771_),
    .A2(net4573),
    .B(net5835),
    .Y(_13773_));
 AOI21x1_ASAP7_75t_R _22038_ (.A1(_13770_),
    .A2(_13773_),
    .B(net5828),
    .Y(_13776_));
 NAND2x1_ASAP7_75t_R _22040_ (.A(net6197),
    .B(net5486),
    .Y(_13778_));
 NAND2x1_ASAP7_75t_R _22041_ (.A(_13778_),
    .B(net4573),
    .Y(_13779_));
 OAI21x1_ASAP7_75t_R _22042_ (.A1(net5844),
    .A2(net6195),
    .B(net4988),
    .Y(_13780_));
 AOI21x1_ASAP7_75t_R _22044_ (.A1(net5840),
    .A2(_13780_),
    .B(net5834),
    .Y(_13782_));
 OAI21x1_ASAP7_75t_R _22045_ (.A1(net5836),
    .A2(_13779_),
    .B(_13782_),
    .Y(_13783_));
 AOI21x1_ASAP7_75t_R _22046_ (.A1(net4921),
    .A2(net4573),
    .B(net5466),
    .Y(_13784_));
 AOI21x1_ASAP7_75t_R _22047_ (.A1(net4925),
    .A2(_13692_),
    .B(net5836),
    .Y(_13785_));
 OAI21x1_ASAP7_75t_R _22048_ (.A1(_13784_),
    .A2(_13785_),
    .B(net5830),
    .Y(_13786_));
 AOI21x1_ASAP7_75t_R _22049_ (.A1(_13783_),
    .A2(_13786_),
    .B(net5465),
    .Y(_13787_));
 AOI211x1_ASAP7_75t_R _22050_ (.A1(_13767_),
    .A2(_13776_),
    .B(_13787_),
    .C(_13759_),
    .Y(_13788_));
 OAI22x1_ASAP7_75t_R _22051_ (.A1(_13681_),
    .A2(_13726_),
    .B1(_13762_),
    .B2(_13788_),
    .Y(_00064_));
 INVx1_ASAP7_75t_R _22053_ (.A(_13751_),
    .Y(_13790_));
 NOR2x1_ASAP7_75t_R _22054_ (.A(net5843),
    .B(_13790_),
    .Y(_13791_));
 NOR2x1_ASAP7_75t_R _22055_ (.A(net5483),
    .B(net6193),
    .Y(_13792_));
 NAND2x1_ASAP7_75t_R _22056_ (.A(net5481),
    .B(_13792_),
    .Y(_13793_));
 AOI211x1_ASAP7_75t_R _22057_ (.A1(net4681),
    .A2(_13793_),
    .B(net4473),
    .C(net5476),
    .Y(_13794_));
 INVx1_ASAP7_75t_R _22058_ (.A(net4763),
    .Y(_13795_));
 AOI21x1_ASAP7_75t_R _22059_ (.A1(net6197),
    .A2(net5847),
    .B(net5481),
    .Y(_13796_));
 NOR2x1_ASAP7_75t_R _22060_ (.A(_13795_),
    .B(_13796_),
    .Y(_13797_));
 NOR2x1_ASAP7_75t_R _22061_ (.A(net5065),
    .B(net5480),
    .Y(_13798_));
 OAI21x1_ASAP7_75t_R _22062_ (.A1(_13798_),
    .A2(_13733_),
    .B(net5473),
    .Y(_13799_));
 OAI21x1_ASAP7_75t_R _22063_ (.A1(net5473),
    .A2(_13797_),
    .B(_13799_),
    .Y(_13800_));
 OAI21x1_ASAP7_75t_R _22064_ (.A1(net5832),
    .A2(_13800_),
    .B(net5828),
    .Y(_13801_));
 NOR2x1_ASAP7_75t_R _22065_ (.A(net5847),
    .B(net5487),
    .Y(_13802_));
 OAI21x1_ASAP7_75t_R _22066_ (.A1(_13702_),
    .A2(_13802_),
    .B(net5474),
    .Y(_13803_));
 INVx1_ASAP7_75t_R _22067_ (.A(_13754_),
    .Y(_13804_));
 NOR2x1_ASAP7_75t_R _22068_ (.A(net6193),
    .B(net5482),
    .Y(_13805_));
 OAI21x1_ASAP7_75t_R _22069_ (.A1(_13804_),
    .A2(_13805_),
    .B(net5843),
    .Y(_13806_));
 AOI21x1_ASAP7_75t_R _22070_ (.A1(_13803_),
    .A2(net4447),
    .B(net5476),
    .Y(_13807_));
 AO21x1_ASAP7_75t_R _22071_ (.A1(net4925),
    .A2(net4574),
    .B(net5474),
    .Y(_13808_));
 OAI21x1_ASAP7_75t_R _22072_ (.A1(net5178),
    .A2(net4922),
    .B(net5474),
    .Y(_13809_));
 AOI21x1_ASAP7_75t_R _22073_ (.A1(_13808_),
    .A2(_13809_),
    .B(net5832),
    .Y(_13810_));
 OAI21x1_ASAP7_75t_R _22074_ (.A1(_13807_),
    .A2(_13810_),
    .B(net5465),
    .Y(_13811_));
 OAI21x1_ASAP7_75t_R _22075_ (.A1(_13794_),
    .A2(_13801_),
    .B(_13811_),
    .Y(_13812_));
 AOI21x1_ASAP7_75t_R _22076_ (.A1(net5182),
    .A2(_13755_),
    .B(net5472),
    .Y(_13813_));
 OAI21x1_ASAP7_75t_R _22077_ (.A1(_01147_),
    .A2(net5480),
    .B(net5466),
    .Y(_13814_));
 OAI21x1_ASAP7_75t_R _22078_ (.A1(_13802_),
    .A2(_13814_),
    .B(net5465),
    .Y(_13815_));
 OAI21x1_ASAP7_75t_R _22079_ (.A1(net5483),
    .A2(net5487),
    .B(net5472),
    .Y(_13816_));
 OAI21x1_ASAP7_75t_R _22080_ (.A1(net5174),
    .A2(_13816_),
    .B(net5828),
    .Y(_13817_));
 INVx1_ASAP7_75t_R _22081_ (.A(_13806_),
    .Y(_13818_));
 OAI22x1_ASAP7_75t_R _22082_ (.A1(_13813_),
    .A2(_13815_),
    .B1(_13817_),
    .B2(_13818_),
    .Y(_13819_));
 NAND2x1_ASAP7_75t_R _22083_ (.A(net5847),
    .B(net6197),
    .Y(_13820_));
 NOR2x1_ASAP7_75t_R _22084_ (.A(net5486),
    .B(_13820_),
    .Y(_13821_));
 AOI21x1_ASAP7_75t_R _22085_ (.A1(_13768_),
    .A2(net5486),
    .B(net5843),
    .Y(_13822_));
 INVx1_ASAP7_75t_R _22086_ (.A(_13822_),
    .Y(_13823_));
 NAND3x1_ASAP7_75t_R _22087_ (.A(net5835),
    .B(net5828),
    .C(_01163_),
    .Y(_13824_));
 OAI21x1_ASAP7_75t_R _22088_ (.A1(_13821_),
    .A2(_13823_),
    .B(_13824_),
    .Y(_13825_));
 OAI21x1_ASAP7_75t_R _22089_ (.A1(net5476),
    .A2(_13825_),
    .B(net6194),
    .Y(_13826_));
 AOI21x1_ASAP7_75t_R _22090_ (.A1(net5476),
    .A2(_13819_),
    .B(_13826_),
    .Y(_13827_));
 AOI21x1_ASAP7_75t_R _22091_ (.A1(net5826),
    .A2(_13812_),
    .B(_13827_),
    .Y(_13828_));
 NAND3x1_ASAP7_75t_R _22093_ (.A(net5179),
    .B(net5177),
    .C(net5469),
    .Y(_13830_));
 NOR2x1_ASAP7_75t_R _22094_ (.A(net5480),
    .B(net5475),
    .Y(_13831_));
 AOI21x1_ASAP7_75t_R _22095_ (.A1(net5181),
    .A2(_13831_),
    .B(net5479),
    .Y(_13832_));
 AOI21x1_ASAP7_75t_R _22096_ (.A1(_13830_),
    .A2(_13832_),
    .B(_13759_),
    .Y(_13833_));
 AO21x1_ASAP7_75t_R _22097_ (.A1(_13751_),
    .A2(net4682),
    .B(net5843),
    .Y(_13834_));
 OA21x2_ASAP7_75t_R _22098_ (.A1(_13620_),
    .A2(_13790_),
    .B(net5479),
    .Y(_13835_));
 NAND2x1_ASAP7_75t_R _22099_ (.A(_13834_),
    .B(_13835_),
    .Y(_13836_));
 AOI21x1_ASAP7_75t_R _22100_ (.A1(_13833_),
    .A2(_13836_),
    .B(net5828),
    .Y(_13837_));
 NOR2x1_ASAP7_75t_R _22101_ (.A(net5473),
    .B(_13797_),
    .Y(_13838_));
 AO21x1_ASAP7_75t_R _22102_ (.A1(net4520),
    .A2(net5473),
    .B(net5476),
    .Y(_13839_));
 INVx1_ASAP7_75t_R _22103_ (.A(_13635_),
    .Y(_13840_));
 NAND2x1_ASAP7_75t_R _22104_ (.A(net5472),
    .B(_13840_),
    .Y(_13841_));
 AOI21x1_ASAP7_75t_R _22105_ (.A1(net5291),
    .A2(net5486),
    .B(net5475),
    .Y(_13842_));
 AOI21x1_ASAP7_75t_R _22106_ (.A1(_13736_),
    .A2(_13842_),
    .B(net5834),
    .Y(_13843_));
 AOI21x1_ASAP7_75t_R _22107_ (.A1(_13841_),
    .A2(_13843_),
    .B(net6194),
    .Y(_13844_));
 OAI21x1_ASAP7_75t_R _22108_ (.A1(_13838_),
    .A2(_13839_),
    .B(_13844_),
    .Y(_13845_));
 NAND2x1_ASAP7_75t_R _22109_ (.A(_13837_),
    .B(_13845_),
    .Y(_13846_));
 NOR2x1_ASAP7_75t_R _22110_ (.A(net6197),
    .B(net5486),
    .Y(_13847_));
 AOI21x1_ASAP7_75t_R _22111_ (.A1(net5837),
    .A2(_13778_),
    .B(_13847_),
    .Y(_13848_));
 NOR2x1_ASAP7_75t_R _22112_ (.A(net5834),
    .B(_13618_),
    .Y(_13849_));
 AOI21x1_ASAP7_75t_R _22113_ (.A1(_13848_),
    .A2(_13849_),
    .B(_13759_),
    .Y(_13850_));
 OAI21x1_ASAP7_75t_R _22114_ (.A1(net5291),
    .A2(net5485),
    .B(net4575),
    .Y(_13851_));
 AOI21x1_ASAP7_75t_R _22115_ (.A1(net5839),
    .A2(_13851_),
    .B(net5479),
    .Y(_13852_));
 NAND2x1_ASAP7_75t_R _22116_ (.A(_13852_),
    .B(_13645_),
    .Y(_13853_));
 AOI21x1_ASAP7_75t_R _22117_ (.A1(_13850_),
    .A2(_13853_),
    .B(net5465),
    .Y(_13854_));
 AO21x1_ASAP7_75t_R _22118_ (.A1(_13746_),
    .A2(_13820_),
    .B(net5473),
    .Y(_13855_));
 NAND2x1p5_ASAP7_75t_R _22119_ (.A(net5474),
    .B(net4574),
    .Y(_13856_));
 OA21x2_ASAP7_75t_R _22120_ (.A1(_13856_),
    .A2(_13802_),
    .B(net5834),
    .Y(_13857_));
 NAND2x1_ASAP7_75t_R _22121_ (.A(_13855_),
    .B(_13857_),
    .Y(_13858_));
 AOI21x1_ASAP7_75t_R _22122_ (.A1(net4684),
    .A2(net4762),
    .B(net5469),
    .Y(_13859_));
 AOI21x1_ASAP7_75t_R _22123_ (.A1(net5469),
    .A2(_13649_),
    .B(_13859_),
    .Y(_13860_));
 AOI21x1_ASAP7_75t_R _22124_ (.A1(net5479),
    .A2(_13860_),
    .B(net6194),
    .Y(_13861_));
 NAND2x1_ASAP7_75t_R _22125_ (.A(_13858_),
    .B(_13861_),
    .Y(_13862_));
 AOI21x1_ASAP7_75t_R _22126_ (.A1(_13854_),
    .A2(_13862_),
    .B(net6192),
    .Y(_13863_));
 NAND2x1_ASAP7_75t_R _22127_ (.A(_13846_),
    .B(_13863_),
    .Y(_13864_));
 OAI21x1_ASAP7_75t_R _22128_ (.A1(_13725_),
    .A2(_13828_),
    .B(_13864_),
    .Y(_00065_));
 NAND3x1_ASAP7_75t_R _22129_ (.A(net5179),
    .B(net5177),
    .C(net5835),
    .Y(_13865_));
 AOI21x1_ASAP7_75t_R _22130_ (.A1(net5831),
    .A2(_13865_),
    .B(net5465),
    .Y(_13866_));
 AND3x1_ASAP7_75t_R _22131_ (.A(net5471),
    .B(net5828),
    .C(_01163_),
    .Y(_13867_));
 NOR2x1_ASAP7_75t_R _22132_ (.A(_13768_),
    .B(net5487),
    .Y(_13868_));
 NOR3x1_ASAP7_75t_R _22133_ (.A(_13868_),
    .B(net5471),
    .C(_13711_),
    .Y(_13869_));
 NOR2x1_ASAP7_75t_R _22134_ (.A(_13702_),
    .B(_13713_),
    .Y(_13870_));
 OAI21x1_ASAP7_75t_R _22135_ (.A1(_13869_),
    .A2(_13870_),
    .B(net5476),
    .Y(_13871_));
 OAI21x1_ASAP7_75t_R _22136_ (.A1(_13866_),
    .A2(_13867_),
    .B(_13871_),
    .Y(_13872_));
 OA21x2_ASAP7_75t_R _22137_ (.A1(net5836),
    .A2(_01161_),
    .B(net5834),
    .Y(_13873_));
 AO21x1_ASAP7_75t_R _22138_ (.A1(_13643_),
    .A2(net4575),
    .B(net5466),
    .Y(_13874_));
 AOI21x1_ASAP7_75t_R _22139_ (.A1(_13873_),
    .A2(_13874_),
    .B(net5828),
    .Y(_13875_));
 NAND2x1_ASAP7_75t_R _22140_ (.A(net6193),
    .B(net5486),
    .Y(_13876_));
 NAND2x1_ASAP7_75t_R _22141_ (.A(net5840),
    .B(_13876_),
    .Y(_13877_));
 NAND2x1_ASAP7_75t_R _22142_ (.A(_13780_),
    .B(_13736_),
    .Y(_13878_));
 AOI21x1_ASAP7_75t_R _22143_ (.A1(net5466),
    .A2(_13878_),
    .B(net5831),
    .Y(_13879_));
 OAI21x1_ASAP7_75t_R _22144_ (.A1(_13802_),
    .A2(_13877_),
    .B(_13879_),
    .Y(_13880_));
 AOI21x1_ASAP7_75t_R _22145_ (.A1(_13875_),
    .A2(_13880_),
    .B(net6194),
    .Y(_13881_));
 NAND2x1_ASAP7_75t_R _22146_ (.A(_13872_),
    .B(_13881_),
    .Y(_13882_));
 INVx1_ASAP7_75t_R _22148_ (.A(_13735_),
    .Y(_13884_));
 AND3x1_ASAP7_75t_R _22150_ (.A(_13638_),
    .B(_13637_),
    .C(_01160_),
    .Y(_13886_));
 AO21x1_ASAP7_75t_R _22151_ (.A1(_13884_),
    .A2(net5475),
    .B(_13886_),
    .Y(_13887_));
 AO21x1_ASAP7_75t_R _22152_ (.A1(net4683),
    .A2(net4573),
    .B(net5466),
    .Y(_13888_));
 OA21x2_ASAP7_75t_R _22153_ (.A1(net5835),
    .A2(_13648_),
    .B(net5465),
    .Y(_13889_));
 AOI21x1_ASAP7_75t_R _22154_ (.A1(_13888_),
    .A2(_13889_),
    .B(net5476),
    .Y(_13890_));
 OAI21x1_ASAP7_75t_R _22155_ (.A1(net5465),
    .A2(_13887_),
    .B(_13890_),
    .Y(_13891_));
 OA21x2_ASAP7_75t_R _22156_ (.A1(net5835),
    .A2(_01165_),
    .B(net5828),
    .Y(_13892_));
 AO21x1_ASAP7_75t_R _22157_ (.A1(net5487),
    .A2(net5847),
    .B(net6193),
    .Y(_13893_));
 NAND2x1_ASAP7_75t_R _22158_ (.A(net5835),
    .B(_13893_),
    .Y(_13894_));
 AOI21x1_ASAP7_75t_R _22159_ (.A1(_13892_),
    .A2(_13894_),
    .B(net5831),
    .Y(_13895_));
 AND2x2_ASAP7_75t_R _22160_ (.A(_01149_),
    .B(net5064),
    .Y(_13896_));
 NOR2x1_ASAP7_75t_R _22161_ (.A(_13896_),
    .B(net5486),
    .Y(_13897_));
 OAI21x1_ASAP7_75t_R _22162_ (.A1(_13897_),
    .A2(_13796_),
    .B(net5842),
    .Y(_13898_));
 AOI21x1_ASAP7_75t_R _22163_ (.A1(_13822_),
    .A2(_13793_),
    .B(net5828),
    .Y(_13899_));
 NAND2x1_ASAP7_75t_R _22164_ (.A(_13898_),
    .B(_13899_),
    .Y(_13900_));
 AOI21x1_ASAP7_75t_R _22165_ (.A1(_13895_),
    .A2(_13900_),
    .B(net5827),
    .Y(_13901_));
 AOI21x1_ASAP7_75t_R _22166_ (.A1(_13891_),
    .A2(_13901_),
    .B(net6192),
    .Y(_13902_));
 NAND2x1_ASAP7_75t_R _22167_ (.A(_13882_),
    .B(_13902_),
    .Y(_13903_));
 NAND2x1_ASAP7_75t_R _22168_ (.A(_13598_),
    .B(net5840),
    .Y(_13904_));
 NOR2x1_ASAP7_75t_R _22169_ (.A(_13727_),
    .B(_13904_),
    .Y(_13905_));
 NOR2x1_ASAP7_75t_R _22170_ (.A(net5483),
    .B(net5486),
    .Y(_13906_));
 INVx1_ASAP7_75t_R _22171_ (.A(_01156_),
    .Y(_13907_));
 OAI21x1_ASAP7_75t_R _22172_ (.A1(net5844),
    .A2(net6195),
    .B(_13907_),
    .Y(_13908_));
 NAND2x1_ASAP7_75t_R _22173_ (.A(_13908_),
    .B(net5475),
    .Y(_13909_));
 OAI21x1_ASAP7_75t_R _22174_ (.A1(_13906_),
    .A2(_13909_),
    .B(net5479),
    .Y(_13910_));
 NOR2x1_ASAP7_75t_R _22175_ (.A(_13905_),
    .B(_13910_),
    .Y(_13911_));
 AO21x1_ASAP7_75t_R _22176_ (.A1(_13780_),
    .A2(net4573),
    .B(net5468),
    .Y(_13912_));
 NOR2x1_ASAP7_75t_R _22177_ (.A(net5292),
    .B(net5482),
    .Y(_13913_));
 OAI21x1_ASAP7_75t_R _22178_ (.A1(_13906_),
    .A2(_13913_),
    .B(net5468),
    .Y(_13914_));
 AOI21x1_ASAP7_75t_R _22179_ (.A1(_13912_),
    .A2(_13914_),
    .B(net5476),
    .Y(_13915_));
 OAI21x1_ASAP7_75t_R _22180_ (.A1(_13911_),
    .A2(_13915_),
    .B(net5464),
    .Y(_13916_));
 NOR2x1_ASAP7_75t_R _22181_ (.A(net6193),
    .B(net5487),
    .Y(_13917_));
 INVx1_ASAP7_75t_R _22182_ (.A(_13616_),
    .Y(_13918_));
 OA21x2_ASAP7_75t_R _22183_ (.A1(_13917_),
    .A2(_13918_),
    .B(net5841),
    .Y(_13919_));
 INVx1_ASAP7_75t_R _22184_ (.A(net4928),
    .Y(_13920_));
 AO21x1_ASAP7_75t_R _22185_ (.A1(net5475),
    .A2(_13920_),
    .B(_13632_),
    .Y(_13921_));
 NAND2x1_ASAP7_75t_R _22186_ (.A(net4685),
    .B(net5840),
    .Y(_13922_));
 OAI21x1_ASAP7_75t_R _22187_ (.A1(_13906_),
    .A2(_13922_),
    .B(_13909_),
    .Y(_13923_));
 AOI21x1_ASAP7_75t_R _22188_ (.A1(_13614_),
    .A2(_13923_),
    .B(net5465),
    .Y(_13924_));
 OAI21x1_ASAP7_75t_R _22189_ (.A1(_13919_),
    .A2(_13921_),
    .B(_13924_),
    .Y(_13925_));
 AOI21x1_ASAP7_75t_R _22190_ (.A1(_13916_),
    .A2(_13925_),
    .B(net6194),
    .Y(_13926_));
 AO21x1_ASAP7_75t_R _22191_ (.A1(net5179),
    .A2(net4574),
    .B(net5840),
    .Y(_13927_));
 AO21x1_ASAP7_75t_R _22192_ (.A1(_13643_),
    .A2(net4683),
    .B(net5466),
    .Y(_13928_));
 AOI21x1_ASAP7_75t_R _22193_ (.A1(_13927_),
    .A2(_13928_),
    .B(net5477),
    .Y(_13929_));
 AOI21x1_ASAP7_75t_R _22194_ (.A1(net4918),
    .A2(_13754_),
    .B(net5843),
    .Y(_13930_));
 AOI21x1_ASAP7_75t_R _22195_ (.A1(net5843),
    .A2(_13893_),
    .B(_13930_),
    .Y(_13931_));
 OAI21x1_ASAP7_75t_R _22196_ (.A1(net5830),
    .A2(_13931_),
    .B(net5828),
    .Y(_13932_));
 NOR2x1_ASAP7_75t_R _22197_ (.A(_13929_),
    .B(_13932_),
    .Y(_13933_));
 OAI21x1_ASAP7_75t_R _22198_ (.A1(_13733_),
    .A2(_13796_),
    .B(net5843),
    .Y(_13934_));
 AO21x1_ASAP7_75t_R _22199_ (.A1(_13805_),
    .A2(net5483),
    .B(net5843),
    .Y(_13935_));
 AOI21x1_ASAP7_75t_R _22200_ (.A1(_13934_),
    .A2(_13935_),
    .B(net5476),
    .Y(_13936_));
 NAND2x1p5_ASAP7_75t_R _22201_ (.A(net5475),
    .B(_13772_),
    .Y(_13937_));
 OAI21x1_ASAP7_75t_R _22202_ (.A1(_13727_),
    .A2(_13937_),
    .B(net5476),
    .Y(_13938_));
 NOR3x1_ASAP7_75t_R _22203_ (.A(_13906_),
    .B(_13798_),
    .C(net5468),
    .Y(_13939_));
 OAI21x1_ASAP7_75t_R _22204_ (.A1(_13939_),
    .A2(_13938_),
    .B(net5464),
    .Y(_13940_));
 OAI21x1_ASAP7_75t_R _22205_ (.A1(_13936_),
    .A2(_13940_),
    .B(net6194),
    .Y(_13941_));
 NOR2x1_ASAP7_75t_R _22206_ (.A(_13933_),
    .B(_13941_),
    .Y(_13942_));
 OAI21x1_ASAP7_75t_R _22207_ (.A1(_13926_),
    .A2(_13942_),
    .B(net6192),
    .Y(_13943_));
 NAND2x1_ASAP7_75t_R _22208_ (.A(_13903_),
    .B(_13943_),
    .Y(_00066_));
 NAND2x1_ASAP7_75t_R _22209_ (.A(_13768_),
    .B(net5486),
    .Y(_13944_));
 NAND2x1_ASAP7_75t_R _22210_ (.A(net5179),
    .B(_13944_),
    .Y(_13945_));
 AO21x1_ASAP7_75t_R _22211_ (.A1(net5842),
    .A2(_13780_),
    .B(net5465),
    .Y(_13946_));
 AO21x1_ASAP7_75t_R _22212_ (.A1(net5469),
    .A2(_13945_),
    .B(_13946_),
    .Y(_13947_));
 OR3x1_ASAP7_75t_R _22213_ (.A(net5840),
    .B(net5828),
    .C(net4762),
    .Y(_13948_));
 NAND2x1_ASAP7_75t_R _22214_ (.A(net5840),
    .B(net4924),
    .Y(_13949_));
 AND2x2_ASAP7_75t_R _22215_ (.A(_13948_),
    .B(_13949_),
    .Y(_13950_));
 AOI21x1_ASAP7_75t_R _22216_ (.A1(_13947_),
    .A2(_13950_),
    .B(net5833),
    .Y(_13951_));
 OA21x2_ASAP7_75t_R _22217_ (.A1(net5470),
    .A2(net4928),
    .B(net5465),
    .Y(_13952_));
 AO21x1_ASAP7_75t_R _22218_ (.A1(_13914_),
    .A2(_13952_),
    .B(net5479),
    .Y(_13953_));
 AO21x1_ASAP7_75t_R _22219_ (.A1(net5169),
    .A2(net5486),
    .B(_13897_),
    .Y(_13954_));
 AND3x1_ASAP7_75t_R _22220_ (.A(_13751_),
    .B(net5469),
    .C(net4763),
    .Y(_13955_));
 AOI211x1_ASAP7_75t_R _22221_ (.A1(_13954_),
    .A2(net5842),
    .B(_13955_),
    .C(net5464),
    .Y(_13956_));
 OAI21x1_ASAP7_75t_R _22222_ (.A1(_13953_),
    .A2(_13956_),
    .B(net6194),
    .Y(_13957_));
 NOR2x1_ASAP7_75t_R _22223_ (.A(_13951_),
    .B(_13957_),
    .Y(_13958_));
 NAND2x1_ASAP7_75t_R _22224_ (.A(net5843),
    .B(_13649_),
    .Y(_13959_));
 AO21x1_ASAP7_75t_R _22225_ (.A1(_13830_),
    .A2(_13959_),
    .B(net5479),
    .Y(_13960_));
 AND3x1_ASAP7_75t_R _22226_ (.A(_13742_),
    .B(net5469),
    .C(net4763),
    .Y(_13961_));
 OA21x2_ASAP7_75t_R _22227_ (.A1(_13790_),
    .A2(_13920_),
    .B(net5843),
    .Y(_13962_));
 OAI21x1_ASAP7_75t_R _22228_ (.A1(_13961_),
    .A2(_13962_),
    .B(net5479),
    .Y(_13963_));
 AOI21x1_ASAP7_75t_R _22229_ (.A1(_13960_),
    .A2(_13963_),
    .B(net5828),
    .Y(_13964_));
 OAI21x1_ASAP7_75t_R _22230_ (.A1(_13913_),
    .A2(_13897_),
    .B(net5842),
    .Y(_13965_));
 OAI21x1_ASAP7_75t_R _22231_ (.A1(_13821_),
    .A2(_13823_),
    .B(_13965_),
    .Y(_13966_));
 INVx1_ASAP7_75t_R _22232_ (.A(_13910_),
    .Y(_13967_));
 AOI21x1_ASAP7_75t_R _22233_ (.A1(net5832),
    .A2(_13966_),
    .B(_13967_),
    .Y(_13968_));
 OAI21x1_ASAP7_75t_R _22234_ (.A1(net5464),
    .A2(_13968_),
    .B(net5826),
    .Y(_13969_));
 OAI21x1_ASAP7_75t_R _22235_ (.A1(_13964_),
    .A2(_13969_),
    .B(net6192),
    .Y(_13970_));
 OAI21x1_ASAP7_75t_R _22236_ (.A1(_13856_),
    .A2(_13840_),
    .B(net5830),
    .Y(_13971_));
 AOI211x1_ASAP7_75t_R _22237_ (.A1(net5181),
    .A2(net5487),
    .B(_13868_),
    .C(net5472),
    .Y(_13972_));
 NOR2x1_ASAP7_75t_R _22238_ (.A(_13972_),
    .B(_13971_),
    .Y(_13973_));
 AO21x1_ASAP7_75t_R _22239_ (.A1(_13633_),
    .A2(net5181),
    .B(net5467),
    .Y(_13974_));
 AO21x1_ASAP7_75t_R _22240_ (.A1(_13692_),
    .A2(net4761),
    .B(net5843),
    .Y(_13975_));
 AOI21x1_ASAP7_75t_R _22241_ (.A1(_13974_),
    .A2(_13975_),
    .B(net5830),
    .Y(_13976_));
 OAI21x1_ASAP7_75t_R _22242_ (.A1(_13973_),
    .A2(_13976_),
    .B(net5465),
    .Y(_13977_));
 NAND2x1_ASAP7_75t_R _22243_ (.A(net5482),
    .B(net5835),
    .Y(_13978_));
 INVx1_ASAP7_75t_R _22244_ (.A(_13764_),
    .Y(_13979_));
 OAI21x1_ASAP7_75t_R _22245_ (.A1(net5483),
    .A2(net5482),
    .B(net5834),
    .Y(_13980_));
 NOR2x1_ASAP7_75t_R _22246_ (.A(_13979_),
    .B(_13980_),
    .Y(_13981_));
 AOI21x1_ASAP7_75t_R _22247_ (.A1(_13978_),
    .A2(_13981_),
    .B(net5465),
    .Y(_13982_));
 NOR2x1_ASAP7_75t_R _22248_ (.A(net5184),
    .B(net5482),
    .Y(_13983_));
 OAI21x1_ASAP7_75t_R _22249_ (.A1(net4916),
    .A2(_13937_),
    .B(_13843_),
    .Y(_13984_));
 AOI21x1_ASAP7_75t_R _22250_ (.A1(_13982_),
    .A2(_13984_),
    .B(net6194),
    .Y(_13985_));
 NAND2x1_ASAP7_75t_R _22251_ (.A(_13985_),
    .B(_13977_),
    .Y(_13986_));
 OAI21x1_ASAP7_75t_R _22252_ (.A1(_13795_),
    .A2(_13805_),
    .B(net5474),
    .Y(_13987_));
 OAI21x1_ASAP7_75t_R _22253_ (.A1(_13918_),
    .A2(_13733_),
    .B(net5843),
    .Y(_13988_));
 AOI21x1_ASAP7_75t_R _22254_ (.A1(_13987_),
    .A2(_13988_),
    .B(net5476),
    .Y(_13989_));
 AO21x1_ASAP7_75t_R _22255_ (.A1(net4925),
    .A2(_13780_),
    .B(net5467),
    .Y(_13990_));
 OAI21x1_ASAP7_75t_R _22256_ (.A1(net5178),
    .A2(_13868_),
    .B(net5472),
    .Y(_13991_));
 AOI21x1_ASAP7_75t_R _22257_ (.A1(_13990_),
    .A2(_13991_),
    .B(net5830),
    .Y(_13992_));
 OAI21x1_ASAP7_75t_R _22258_ (.A1(_13989_),
    .A2(_13992_),
    .B(net5465),
    .Y(_13993_));
 OAI21x1_ASAP7_75t_R _22259_ (.A1(_13906_),
    .A2(net5174),
    .B(net5468),
    .Y(_13994_));
 AOI21x1_ASAP7_75t_R _22260_ (.A1(_13782_),
    .A2(_13994_),
    .B(net5465),
    .Y(_13995_));
 AO21x1_ASAP7_75t_R _22261_ (.A1(_13633_),
    .A2(net5177),
    .B(net5843),
    .Y(_13996_));
 AOI21x1_ASAP7_75t_R _22262_ (.A1(net5171),
    .A2(_13621_),
    .B(net5477),
    .Y(_13997_));
 NAND2x1_ASAP7_75t_R _22263_ (.A(_13996_),
    .B(_13997_),
    .Y(_13998_));
 AOI21x1_ASAP7_75t_R _22264_ (.A1(_13995_),
    .A2(_13998_),
    .B(_13759_),
    .Y(_13999_));
 AOI21x1_ASAP7_75t_R _22265_ (.A1(_13993_),
    .A2(_13999_),
    .B(net6192),
    .Y(_14000_));
 NAND2x1_ASAP7_75t_R _22266_ (.A(_14000_),
    .B(_13986_),
    .Y(_14001_));
 OAI21x1_ASAP7_75t_R _22267_ (.A1(_13958_),
    .A2(_13970_),
    .B(_14001_),
    .Y(_00067_));
 NOR2x1_ASAP7_75t_R _22268_ (.A(net5479),
    .B(net4926),
    .Y(_14002_));
 AO21x1_ASAP7_75t_R _22269_ (.A1(_13780_),
    .A2(net4682),
    .B(net5842),
    .Y(_14003_));
 NAND2x1_ASAP7_75t_R _22270_ (.A(net5065),
    .B(net5485),
    .Y(_14004_));
 AO21x1_ASAP7_75t_R _22271_ (.A1(_14004_),
    .A2(net5475),
    .B(net5833),
    .Y(_14005_));
 NOR2x1_ASAP7_75t_R _22272_ (.A(net5481),
    .B(_13820_),
    .Y(_14006_));
 NOR2x1_ASAP7_75t_R _22273_ (.A(net5473),
    .B(_14006_),
    .Y(_14007_));
 OAI21x1_ASAP7_75t_R _22274_ (.A1(_14005_),
    .A2(_14007_),
    .B(net5464),
    .Y(_14008_));
 AOI21x1_ASAP7_75t_R _22275_ (.A1(_14002_),
    .A2(_14003_),
    .B(_14008_),
    .Y(_14009_));
 INVx1_ASAP7_75t_R _22276_ (.A(_13648_),
    .Y(_14010_));
 AO21x1_ASAP7_75t_R _22277_ (.A1(_14010_),
    .A2(net5468),
    .B(net5833),
    .Y(_14011_));
 NOR2x1_ASAP7_75t_R _22278_ (.A(net5837),
    .B(net5171),
    .Y(_14012_));
 NOR3x1_ASAP7_75t_R _22279_ (.A(_13818_),
    .B(_14011_),
    .C(_14012_),
    .Y(_14013_));
 AO21x1_ASAP7_75t_R _22280_ (.A1(_13746_),
    .A2(net4917),
    .B(net5842),
    .Y(_14014_));
 NOR2x1_ASAP7_75t_R _22281_ (.A(net5479),
    .B(_13831_),
    .Y(_14015_));
 AO21x1_ASAP7_75t_R _22282_ (.A1(_14014_),
    .A2(_14015_),
    .B(net5465),
    .Y(_14016_));
 OAI21x1_ASAP7_75t_R _22283_ (.A1(_14013_),
    .A2(_14016_),
    .B(net5825),
    .Y(_14017_));
 NOR2x1_ASAP7_75t_R _22284_ (.A(_14009_),
    .B(_14017_),
    .Y(_14018_));
 NOR2x1_ASAP7_75t_R _22285_ (.A(net5838),
    .B(_13643_),
    .Y(_14019_));
 OAI21x1_ASAP7_75t_R _22286_ (.A1(_13847_),
    .A2(_13689_),
    .B(net5478),
    .Y(_14020_));
 NOR2x1_ASAP7_75t_R _22287_ (.A(_14019_),
    .B(_14020_),
    .Y(_14021_));
 INVx1_ASAP7_75t_R _22288_ (.A(_01155_),
    .Y(_14022_));
 NOR2x1p5_ASAP7_75t_R _22289_ (.A(net5466),
    .B(net4575),
    .Y(_14023_));
 AOI21x1_ASAP7_75t_R _22290_ (.A1(_14022_),
    .A2(net5466),
    .B(_14023_),
    .Y(_14024_));
 OAI21x1_ASAP7_75t_R _22291_ (.A1(net5478),
    .A2(_14024_),
    .B(net5463),
    .Y(_14025_));
 OAI21x1_ASAP7_75t_R _22292_ (.A1(_14021_),
    .A2(_14025_),
    .B(net6194),
    .Y(_14026_));
 NOR2x1_ASAP7_75t_R _22293_ (.A(net5170),
    .B(_13689_),
    .Y(_14027_));
 OA21x2_ASAP7_75t_R _22294_ (.A1(_13847_),
    .A2(net5175),
    .B(net5468),
    .Y(_14028_));
 OAI21x1_ASAP7_75t_R _22295_ (.A1(_14027_),
    .A2(_14028_),
    .B(net5478),
    .Y(_14029_));
 OAI21x1_ASAP7_75t_R _22296_ (.A1(_13765_),
    .A2(_13704_),
    .B(net5834),
    .Y(_14030_));
 AOI21x1_ASAP7_75t_R _22297_ (.A1(_14029_),
    .A2(_14030_),
    .B(net5463),
    .Y(_14031_));
 OAI21x1_ASAP7_75t_R _22298_ (.A1(_14026_),
    .A2(_14031_),
    .B(net6192),
    .Y(_14032_));
 NOR2x1_ASAP7_75t_R _22299_ (.A(net5829),
    .B(net4923),
    .Y(_14033_));
 AO21x1_ASAP7_75t_R _22300_ (.A1(_14033_),
    .A2(_13689_),
    .B(net5828),
    .Y(_14034_));
 NAND2x1_ASAP7_75t_R _22301_ (.A(net5836),
    .B(_13778_),
    .Y(_14035_));
 AOI21x1_ASAP7_75t_R _22302_ (.A1(_13814_),
    .A2(_14035_),
    .B(_13802_),
    .Y(_14036_));
 NOR2x1_ASAP7_75t_R _22303_ (.A(net5477),
    .B(_14036_),
    .Y(_14037_));
 OAI21x1_ASAP7_75t_R _22304_ (.A1(_14034_),
    .A2(_14037_),
    .B(net5825),
    .Y(_14038_));
 NOR2x1_ASAP7_75t_R _22305_ (.A(net5174),
    .B(_13816_),
    .Y(_14039_));
 NAND2x1_ASAP7_75t_R _22306_ (.A(net5843),
    .B(net5177),
    .Y(_14040_));
 NOR2x1_ASAP7_75t_R _22307_ (.A(_13917_),
    .B(_14040_),
    .Y(_14041_));
 OAI21x1_ASAP7_75t_R _22308_ (.A1(_14039_),
    .A2(_14041_),
    .B(net5830),
    .Y(_14042_));
 OA21x2_ASAP7_75t_R _22309_ (.A1(_13917_),
    .A2(_13702_),
    .B(net5841),
    .Y(_14043_));
 NOR2x1_ASAP7_75t_R _22310_ (.A(net5175),
    .B(_13737_),
    .Y(_14044_));
 OAI21x1_ASAP7_75t_R _22311_ (.A1(_14043_),
    .A2(_14044_),
    .B(net5476),
    .Y(_14045_));
 AOI21x1_ASAP7_75t_R _22312_ (.A1(_14042_),
    .A2(_14045_),
    .B(net5464),
    .Y(_14046_));
 OAI21x1_ASAP7_75t_R _22313_ (.A1(_14038_),
    .A2(_14046_),
    .B(_13725_),
    .Y(_14047_));
 NOR2x1_ASAP7_75t_R _22314_ (.A(_13920_),
    .B(_14023_),
    .Y(_14048_));
 AO21x1_ASAP7_75t_R _22315_ (.A1(_14048_),
    .A2(_13849_),
    .B(net5828),
    .Y(_14049_));
 AO21x1_ASAP7_75t_R _22316_ (.A1(_13851_),
    .A2(net5470),
    .B(net5479),
    .Y(_14050_));
 NOR2x1_ASAP7_75t_R _22317_ (.A(_13690_),
    .B(_14050_),
    .Y(_14051_));
 OAI21x1_ASAP7_75t_R _22318_ (.A1(_14051_),
    .A2(_14049_),
    .B(net6194),
    .Y(_14052_));
 OA21x2_ASAP7_75t_R _22319_ (.A1(net5174),
    .A2(_14010_),
    .B(net5841),
    .Y(_14053_));
 OAI21x1_ASAP7_75t_R _22320_ (.A1(net4521),
    .A2(_14053_),
    .B(net5834),
    .Y(_14054_));
 OAI21x1_ASAP7_75t_R _22321_ (.A1(net5486),
    .A2(net5181),
    .B(net5843),
    .Y(_14055_));
 NOR2x1_ASAP7_75t_R _22322_ (.A(_13727_),
    .B(_14055_),
    .Y(_14056_));
 OAI21x1_ASAP7_75t_R _22323_ (.A1(net4519),
    .A2(_14056_),
    .B(net5476),
    .Y(_14057_));
 AOI21x1_ASAP7_75t_R _22324_ (.A1(_14054_),
    .A2(_14057_),
    .B(net5465),
    .Y(_14058_));
 NOR2x1_ASAP7_75t_R _22325_ (.A(_14058_),
    .B(_14052_),
    .Y(_14059_));
 OAI22x1_ASAP7_75t_R _22326_ (.A1(_14018_),
    .A2(_14032_),
    .B1(_14059_),
    .B2(_14047_),
    .Y(_00068_));
 NAND2x1_ASAP7_75t_R _22327_ (.A(net5064),
    .B(net5480),
    .Y(_14060_));
 AOI22x1_ASAP7_75t_R _22328_ (.A1(_13831_),
    .A2(net5181),
    .B1(net5470),
    .B2(_14060_),
    .Y(_14061_));
 AOI21x1_ASAP7_75t_R _22329_ (.A1(net5483),
    .A2(_13831_),
    .B(net5479),
    .Y(_14062_));
 OAI21x1_ASAP7_75t_R _22330_ (.A1(net5840),
    .A2(net4761),
    .B(_13904_),
    .Y(_14063_));
 AO21x1_ASAP7_75t_R _22331_ (.A1(_14062_),
    .A2(_14063_),
    .B(net5465),
    .Y(_14064_));
 AOI21x1_ASAP7_75t_R _22332_ (.A1(net5479),
    .A2(_14061_),
    .B(_14064_),
    .Y(_14065_));
 AOI211x1_ASAP7_75t_R _22333_ (.A1(_14060_),
    .A2(net5172),
    .B(_14012_),
    .C(_13685_),
    .Y(_14066_));
 AOI211x1_ASAP7_75t_R _22334_ (.A1(_13917_),
    .A2(net5483),
    .B(net4916),
    .C(net5841),
    .Y(_14067_));
 OA21x2_ASAP7_75t_R _22335_ (.A1(net5470),
    .A2(net5064),
    .B(net5479),
    .Y(_14068_));
 NAND2x1_ASAP7_75t_R _22336_ (.A(_13949_),
    .B(_14068_),
    .Y(_14069_));
 OAI21x1_ASAP7_75t_R _22337_ (.A1(_14067_),
    .A2(_14069_),
    .B(net5465),
    .Y(_14070_));
 OAI21x1_ASAP7_75t_R _22338_ (.A1(_14066_),
    .A2(_14070_),
    .B(net5825),
    .Y(_14071_));
 OAI21x1_ASAP7_75t_R _22339_ (.A1(_14065_),
    .A2(_14071_),
    .B(_13725_),
    .Y(_14072_));
 AND3x1_ASAP7_75t_R _22340_ (.A(net5179),
    .B(_14004_),
    .C(net5470),
    .Y(_14073_));
 OAI21x1_ASAP7_75t_R _22341_ (.A1(net4469),
    .A2(_14073_),
    .B(net5478),
    .Y(_14074_));
 NAND2x1_ASAP7_75t_R _22342_ (.A(net5829),
    .B(_13909_),
    .Y(_14075_));
 AO21x1_ASAP7_75t_R _22343_ (.A1(net4474),
    .A2(net4921),
    .B(_14075_),
    .Y(_14076_));
 NAND3x1_ASAP7_75t_R _22344_ (.A(_14074_),
    .B(net5828),
    .C(_14076_),
    .Y(_14077_));
 NAND2x1_ASAP7_75t_R _22345_ (.A(_13820_),
    .B(_13791_),
    .Y(_14078_));
 AO21x1_ASAP7_75t_R _22346_ (.A1(_13793_),
    .A2(_13944_),
    .B(net5473),
    .Y(_14079_));
 AOI21x1_ASAP7_75t_R _22347_ (.A1(_14078_),
    .A2(_14079_),
    .B(net5832),
    .Y(_14080_));
 AOI211x1_ASAP7_75t_R _22348_ (.A1(net6197),
    .A2(net5842),
    .B(_14044_),
    .C(net5476),
    .Y(_14081_));
 OAI21x1_ASAP7_75t_R _22349_ (.A1(_14080_),
    .A2(_14081_),
    .B(net5464),
    .Y(_14082_));
 AOI21x1_ASAP7_75t_R _22350_ (.A1(_14077_),
    .A2(_14082_),
    .B(net5825),
    .Y(_14083_));
 AND2x2_ASAP7_75t_R _22351_ (.A(net5480),
    .B(_13896_),
    .Y(_14084_));
 OAI21x1_ASAP7_75t_R _22352_ (.A1(net5468),
    .A2(_14084_),
    .B(net5833),
    .Y(_14085_));
 NOR2x1_ASAP7_75t_R _22353_ (.A(_13821_),
    .B(_13935_),
    .Y(_14086_));
 INVx1_ASAP7_75t_R _22354_ (.A(net5173),
    .Y(_14087_));
 AOI21x1_ASAP7_75t_R _22355_ (.A1(_14087_),
    .A2(_13849_),
    .B(net5828),
    .Y(_14088_));
 OAI21x1_ASAP7_75t_R _22356_ (.A1(_14085_),
    .A2(_14086_),
    .B(_14088_),
    .Y(_14089_));
 NAND2x1_ASAP7_75t_R _22357_ (.A(net4762),
    .B(net4917),
    .Y(_14090_));
 AOI21x1_ASAP7_75t_R _22358_ (.A1(net5473),
    .A2(_14090_),
    .B(net5832),
    .Y(_14091_));
 NAND2x1_ASAP7_75t_R _22359_ (.A(_13944_),
    .B(_13621_),
    .Y(_14092_));
 NAND2x1_ASAP7_75t_R _22360_ (.A(_14091_),
    .B(_14092_),
    .Y(_14093_));
 OA21x2_ASAP7_75t_R _22361_ (.A1(net5474),
    .A2(_13768_),
    .B(net5834),
    .Y(_14094_));
 AO21x1_ASAP7_75t_R _22362_ (.A1(net5175),
    .A2(net5481),
    .B(net5843),
    .Y(_14095_));
 AOI21x1_ASAP7_75t_R _22363_ (.A1(_14094_),
    .A2(_14095_),
    .B(net5465),
    .Y(_14096_));
 AOI21x1_ASAP7_75t_R _22364_ (.A1(_14093_),
    .A2(_14096_),
    .B(_13759_),
    .Y(_14097_));
 AOI21x1_ASAP7_75t_R _22365_ (.A1(_14089_),
    .A2(_14097_),
    .B(_13725_),
    .Y(_14098_));
 NOR2x1_ASAP7_75t_R _22366_ (.A(net5840),
    .B(_13707_),
    .Y(_14099_));
 OA21x2_ASAP7_75t_R _22367_ (.A1(_13692_),
    .A2(net5466),
    .B(net5478),
    .Y(_14100_));
 AO21x1_ASAP7_75t_R _22368_ (.A1(_13635_),
    .A2(net4917),
    .B(net5837),
    .Y(_14101_));
 AOI21x1_ASAP7_75t_R _22369_ (.A1(_14100_),
    .A2(_14101_),
    .B(net5465),
    .Y(_14102_));
 OAI21x1_ASAP7_75t_R _22370_ (.A1(_13642_),
    .A2(_14099_),
    .B(_14102_),
    .Y(_14103_));
 OA21x2_ASAP7_75t_R _22371_ (.A1(net5467),
    .A2(net5483),
    .B(net5834),
    .Y(_14104_));
 AOI21x1_ASAP7_75t_R _22372_ (.A1(_14104_),
    .A2(_13763_),
    .B(net5828),
    .Y(_14105_));
 NAND2x1_ASAP7_75t_R _22373_ (.A(_13621_),
    .B(_13884_),
    .Y(_14106_));
 NOR2x1_ASAP7_75t_R _22374_ (.A(net5843),
    .B(_13983_),
    .Y(_14107_));
 AOI21x1_ASAP7_75t_R _22375_ (.A1(_13736_),
    .A2(_14107_),
    .B(net5830),
    .Y(_14108_));
 NAND2x1_ASAP7_75t_R _22376_ (.A(_14106_),
    .B(_14108_),
    .Y(_14109_));
 AOI21x1_ASAP7_75t_R _22377_ (.A1(_14105_),
    .A2(_14109_),
    .B(net6194),
    .Y(_14110_));
 NAND2x1_ASAP7_75t_R _22378_ (.A(_14103_),
    .B(_14110_),
    .Y(_14111_));
 NAND2x1_ASAP7_75t_R _22379_ (.A(_14098_),
    .B(_14111_),
    .Y(_14112_));
 OAI21x1_ASAP7_75t_R _22380_ (.A1(_14072_),
    .A2(_14083_),
    .B(_14112_),
    .Y(_00069_));
 OAI21x1_ASAP7_75t_R _22381_ (.A1(net5169),
    .A2(net5486),
    .B(net5467),
    .Y(_14113_));
 NOR2x1_ASAP7_75t_R _22382_ (.A(net4916),
    .B(_14113_),
    .Y(_14114_));
 OA21x2_ASAP7_75t_R _22383_ (.A1(_13796_),
    .A2(net4922),
    .B(net5841),
    .Y(_14115_));
 NOR2x1_ASAP7_75t_R _22384_ (.A(_14114_),
    .B(_14115_),
    .Y(_14116_));
 AND4x1_ASAP7_75t_R _22385_ (.A(_13652_),
    .B(net5838),
    .C(_13616_),
    .D(net4928),
    .Y(_14117_));
 AO21x1_ASAP7_75t_R _22386_ (.A1(net5466),
    .A2(net5170),
    .B(_13661_),
    .Y(_14118_));
 OAI22x1_ASAP7_75t_R _22387_ (.A1(_14116_),
    .A2(net5478),
    .B1(_14117_),
    .B2(_14118_),
    .Y(_14119_));
 NAND2x1_ASAP7_75t_R _22388_ (.A(_01158_),
    .B(_01164_),
    .Y(_14120_));
 AO21x1_ASAP7_75t_R _22389_ (.A1(net5466),
    .A2(_14120_),
    .B(net5477),
    .Y(_14121_));
 NOR2x1_ASAP7_75t_R _22390_ (.A(_13687_),
    .B(_13877_),
    .Y(_14122_));
 NOR2x1_ASAP7_75t_R _22391_ (.A(_14121_),
    .B(_14122_),
    .Y(_14123_));
 OA21x2_ASAP7_75t_R _22392_ (.A1(_13798_),
    .A2(_13920_),
    .B(net5840),
    .Y(_14124_));
 OAI21x1_ASAP7_75t_R _22393_ (.A1(_14011_),
    .A2(_14124_),
    .B(net5463),
    .Y(_14125_));
 OAI21x1_ASAP7_75t_R _22394_ (.A1(_14123_),
    .A2(_14125_),
    .B(net5824),
    .Y(_14126_));
 AOI21x1_ASAP7_75t_R _22395_ (.A1(net5828),
    .A2(_14119_),
    .B(_14126_),
    .Y(_14127_));
 AOI21x1_ASAP7_75t_R _22396_ (.A1(net4573),
    .A2(_13755_),
    .B(net5835),
    .Y(_14128_));
 OAI21x1_ASAP7_75t_R _22397_ (.A1(_13886_),
    .A2(_14128_),
    .B(net5476),
    .Y(_14129_));
 AOI21x1_ASAP7_75t_R _22398_ (.A1(net5179),
    .A2(_13755_),
    .B(net5467),
    .Y(_14130_));
 AND3x1_ASAP7_75t_R _22399_ (.A(_14004_),
    .B(net5467),
    .C(net4573),
    .Y(_14131_));
 OAI21x1_ASAP7_75t_R _22400_ (.A1(_14130_),
    .A2(_14131_),
    .B(net5830),
    .Y(_14132_));
 AOI21x1_ASAP7_75t_R _22401_ (.A1(_14129_),
    .A2(_14132_),
    .B(net5828),
    .Y(_14133_));
 OA21x2_ASAP7_75t_R _22402_ (.A1(_13692_),
    .A2(net5836),
    .B(net5477),
    .Y(_14134_));
 AO21x1_ASAP7_75t_R _22403_ (.A1(_13707_),
    .A2(net6197),
    .B(net5466),
    .Y(_14135_));
 AO21x1_ASAP7_75t_R _22404_ (.A1(_14134_),
    .A2(_14135_),
    .B(net5465),
    .Y(_14136_));
 INVx1_ASAP7_75t_R _22405_ (.A(_14062_),
    .Y(_14137_));
 NOR2x1_ASAP7_75t_R _22406_ (.A(_13856_),
    .B(_14084_),
    .Y(_14138_));
 NOR3x1_ASAP7_75t_R _22407_ (.A(_14137_),
    .B(_13765_),
    .C(_14138_),
    .Y(_14139_));
 OAI21x1_ASAP7_75t_R _22408_ (.A1(_14136_),
    .A2(_14139_),
    .B(net6194),
    .Y(_14140_));
 OAI21x1_ASAP7_75t_R _22409_ (.A1(_14133_),
    .A2(_14140_),
    .B(_13725_),
    .Y(_14141_));
 AOI21x1_ASAP7_75t_R _22410_ (.A1(_01159_),
    .A2(net5835),
    .B(net5476),
    .Y(_14142_));
 OAI21x1_ASAP7_75t_R _22411_ (.A1(_13913_),
    .A2(_13917_),
    .B(net5466),
    .Y(_14143_));
 AOI21x1_ASAP7_75t_R _22412_ (.A1(_14142_),
    .A2(_14143_),
    .B(_13759_),
    .Y(_14144_));
 AO21x1_ASAP7_75t_R _22413_ (.A1(net4763),
    .A2(net4918),
    .B(net5472),
    .Y(_14145_));
 NAND2x1_ASAP7_75t_R _22414_ (.A(net5472),
    .B(_13731_),
    .Y(_14146_));
 NAND3x1_ASAP7_75t_R _22415_ (.A(_14145_),
    .B(_14146_),
    .C(net5476),
    .Y(_14147_));
 AOI21x1_ASAP7_75t_R _22416_ (.A1(_14144_),
    .A2(_14147_),
    .B(net5828),
    .Y(_14148_));
 AOI21x1_ASAP7_75t_R _22417_ (.A1(_14113_),
    .A2(_14040_),
    .B(net5178),
    .Y(_14149_));
 NAND2x1_ASAP7_75t_R _22418_ (.A(net6193),
    .B(net5471),
    .Y(_14150_));
 AOI21x1_ASAP7_75t_R _22419_ (.A1(_14150_),
    .A2(_13981_),
    .B(net6194),
    .Y(_14151_));
 OAI21x1_ASAP7_75t_R _22420_ (.A1(net5830),
    .A2(_14149_),
    .B(_14151_),
    .Y(_14152_));
 AOI21x1_ASAP7_75t_R _22421_ (.A1(_14148_),
    .A2(_14152_),
    .B(_13725_),
    .Y(_14153_));
 NOR2x1_ASAP7_75t_R _22422_ (.A(net4919),
    .B(_14020_),
    .Y(_14154_));
 AND3x1_ASAP7_75t_R _22423_ (.A(_13643_),
    .B(net5838),
    .C(_13616_),
    .Y(_14155_));
 AO21x1_ASAP7_75t_R _22424_ (.A1(_14155_),
    .A2(net5829),
    .B(net5824),
    .Y(_14156_));
 NAND2x1p5_ASAP7_75t_R _22425_ (.A(net4470),
    .B(net4680),
    .Y(_14157_));
 AOI21x1_ASAP7_75t_R _22426_ (.A1(_14157_),
    .A2(_14062_),
    .B(net6194),
    .Y(_14158_));
 AO21x1_ASAP7_75t_R _22427_ (.A1(net5486),
    .A2(net6193),
    .B(net5846),
    .Y(_14159_));
 AOI21x1_ASAP7_75t_R _22428_ (.A1(net5466),
    .A2(_14159_),
    .B(net5834),
    .Y(_14160_));
 NAND2x1_ASAP7_75t_R _22429_ (.A(_14035_),
    .B(_14160_),
    .Y(_14161_));
 AOI21x1_ASAP7_75t_R _22430_ (.A1(_14161_),
    .A2(_14158_),
    .B(net5463),
    .Y(_14162_));
 OAI21x1_ASAP7_75t_R _22431_ (.A1(_14154_),
    .A2(_14156_),
    .B(_14162_),
    .Y(_14163_));
 NAND2x1_ASAP7_75t_R _22432_ (.A(_14153_),
    .B(_14163_),
    .Y(_14164_));
 OAI21x1_ASAP7_75t_R _22433_ (.A1(_14127_),
    .A2(_14141_),
    .B(_14164_),
    .Y(_00070_));
 AOI211x1_ASAP7_75t_R _22434_ (.A1(net5837),
    .A2(_13727_),
    .B(_13654_),
    .C(_14010_),
    .Y(_14165_));
 AO21x1_ASAP7_75t_R _22435_ (.A1(net4927),
    .A2(net5466),
    .B(net5834),
    .Y(_14166_));
 OAI21x1_ASAP7_75t_R _22436_ (.A1(_14166_),
    .A2(_14122_),
    .B(net5828),
    .Y(_14167_));
 OAI21x1_ASAP7_75t_R _22437_ (.A1(_14165_),
    .A2(_14167_),
    .B(net5824),
    .Y(_14168_));
 INVx1_ASAP7_75t_R _22438_ (.A(_13965_),
    .Y(_14169_));
 OA21x2_ASAP7_75t_R _22439_ (.A1(_13796_),
    .A2(_13847_),
    .B(net5468),
    .Y(_14170_));
 OAI21x1_ASAP7_75t_R _22440_ (.A1(_14169_),
    .A2(_14170_),
    .B(net5476),
    .Y(_14171_));
 AND3x1_ASAP7_75t_R _22441_ (.A(_13944_),
    .B(net5841),
    .C(net4573),
    .Y(_14172_));
 OA21x2_ASAP7_75t_R _22442_ (.A1(_13796_),
    .A2(_14010_),
    .B(net5468),
    .Y(_14173_));
 OAI21x1_ASAP7_75t_R _22443_ (.A1(_14172_),
    .A2(_14173_),
    .B(net5832),
    .Y(_14174_));
 AOI21x1_ASAP7_75t_R _22444_ (.A1(_14171_),
    .A2(_14174_),
    .B(net5828),
    .Y(_14175_));
 NOR2x1_ASAP7_75t_R _22445_ (.A(_14168_),
    .B(_14175_),
    .Y(_14176_));
 AOI21x1_ASAP7_75t_R _22446_ (.A1(net5179),
    .A2(_13633_),
    .B(net5835),
    .Y(_14177_));
 AND3x1_ASAP7_75t_R _22447_ (.A(net5835),
    .B(_13780_),
    .C(net4573),
    .Y(_14178_));
 OAI21x1_ASAP7_75t_R _22448_ (.A1(_14177_),
    .A2(_14178_),
    .B(net5477),
    .Y(_14179_));
 AO21x1_ASAP7_75t_R _22449_ (.A1(net4928),
    .A2(_13780_),
    .B(net5835),
    .Y(_14180_));
 AO21x1_ASAP7_75t_R _22450_ (.A1(_13594_),
    .A2(_13593_),
    .B(_01164_),
    .Y(_14181_));
 AO21x1_ASAP7_75t_R _22451_ (.A1(_14180_),
    .A2(_14181_),
    .B(net5476),
    .Y(_14182_));
 AOI21x1_ASAP7_75t_R _22452_ (.A1(_14179_),
    .A2(_14182_),
    .B(net5465),
    .Y(_14183_));
 NOR2x1_ASAP7_75t_R _22453_ (.A(_14022_),
    .B(net5466),
    .Y(_14184_));
 OAI21x1_ASAP7_75t_R _22454_ (.A1(_14184_),
    .A2(_13654_),
    .B(net5463),
    .Y(_14185_));
 AO21x1_ASAP7_75t_R _22455_ (.A1(net6193),
    .A2(net5466),
    .B(net5834),
    .Y(_14186_));
 AOI211x1_ASAP7_75t_R _22456_ (.A1(_13700_),
    .A2(net5171),
    .B(_14186_),
    .C(_14099_),
    .Y(_14187_));
 OAI21x1_ASAP7_75t_R _22457_ (.A1(_14185_),
    .A2(_14187_),
    .B(net6194),
    .Y(_14188_));
 OAI21x1_ASAP7_75t_R _22458_ (.A1(_14183_),
    .A2(_14188_),
    .B(_13725_),
    .Y(_14189_));
 NOR2x1_ASAP7_75t_R _22459_ (.A(net5472),
    .B(net5182),
    .Y(_14190_));
 AO21x1_ASAP7_75t_R _22460_ (.A1(_13795_),
    .A2(net5474),
    .B(net5476),
    .Y(_14191_));
 OAI21x1_ASAP7_75t_R _22461_ (.A1(_14190_),
    .A2(_14191_),
    .B(net5828),
    .Y(_14192_));
 NOR2x1_ASAP7_75t_R _22462_ (.A(_14006_),
    .B(net4471),
    .Y(_14193_));
 NAND2x1_ASAP7_75t_R _22463_ (.A(net5476),
    .B(_14055_),
    .Y(_14194_));
 NOR2x1_ASAP7_75t_R _22464_ (.A(_14194_),
    .B(_14193_),
    .Y(_14195_));
 OAI21x1_ASAP7_75t_R _22465_ (.A1(_14192_),
    .A2(_14195_),
    .B(net6194),
    .Y(_14196_));
 NOR2x1_ASAP7_75t_R _22466_ (.A(net5483),
    .B(net5835),
    .Y(_14197_));
 OA21x2_ASAP7_75t_R _22467_ (.A1(_13802_),
    .A2(net5174),
    .B(net5835),
    .Y(_14198_));
 OAI21x1_ASAP7_75t_R _22468_ (.A1(_14197_),
    .A2(_14198_),
    .B(net5476),
    .Y(_14199_));
 NOR2x1_ASAP7_75t_R _22469_ (.A(_14006_),
    .B(_13737_),
    .Y(_14200_));
 OAI21x1_ASAP7_75t_R _22470_ (.A1(_14041_),
    .A2(_14200_),
    .B(net5830),
    .Y(_14201_));
 AOI21x1_ASAP7_75t_R _22471_ (.A1(_14199_),
    .A2(_14201_),
    .B(net5828),
    .Y(_14202_));
 OAI21x1_ASAP7_75t_R _22472_ (.A1(_14202_),
    .A2(_14196_),
    .B(net6192),
    .Y(_14203_));
 NAND3x1_ASAP7_75t_R _22473_ (.A(_13736_),
    .B(net5483),
    .C(net5466),
    .Y(_14204_));
 NAND3x1_ASAP7_75t_R _22474_ (.A(_13771_),
    .B(net5835),
    .C(net4925),
    .Y(_14205_));
 AOI21x1_ASAP7_75t_R _22475_ (.A1(_14204_),
    .A2(_14205_),
    .B(net5830),
    .Y(_14206_));
 OAI21x1_ASAP7_75t_R _22476_ (.A1(_13847_),
    .A2(_13689_),
    .B(net4915),
    .Y(_14207_));
 OAI21x1_ASAP7_75t_R _22477_ (.A1(net5477),
    .A2(_14207_),
    .B(net5463),
    .Y(_14208_));
 OAI21x1_ASAP7_75t_R _22478_ (.A1(_14206_),
    .A2(_14208_),
    .B(net5824),
    .Y(_14209_));
 NOR2x1_ASAP7_75t_R _22479_ (.A(_13802_),
    .B(_13877_),
    .Y(_14210_));
 OAI21x1_ASAP7_75t_R _22480_ (.A1(_14114_),
    .A2(_14210_),
    .B(net5834),
    .Y(_14211_));
 AND2x2_ASAP7_75t_R _22481_ (.A(_13851_),
    .B(net5839),
    .Y(_14212_));
 OAI21x1_ASAP7_75t_R _22482_ (.A1(_14212_),
    .A2(_13955_),
    .B(net5479),
    .Y(_14213_));
 AOI21x1_ASAP7_75t_R _22483_ (.A1(_14211_),
    .A2(_14213_),
    .B(net5463),
    .Y(_14214_));
 NOR2x1_ASAP7_75t_R _22484_ (.A(_14209_),
    .B(_14214_),
    .Y(_14215_));
 OAI22x1_ASAP7_75t_R _22485_ (.A1(_14176_),
    .A2(_14189_),
    .B1(_14203_),
    .B2(_14215_),
    .Y(_00071_));
 XOR2x2_ASAP7_75t_R _22486_ (.A(_11399_),
    .B(_00584_),
    .Y(_14216_));
 XOR2x2_ASAP7_75t_R _22487_ (.A(_00654_),
    .B(_00647_),
    .Y(_14217_));
 XOR2x1_ASAP7_75t_R _22488_ (.A(net6591),
    .Y(_14218_),
    .B(_00680_));
 XOR2x2_ASAP7_75t_R _22489_ (.A(_14218_),
    .B(_14217_),
    .Y(_14219_));
 OAI21x1_ASAP7_75t_R _22490_ (.A1(_14216_),
    .A2(_14219_),
    .B(net6669),
    .Y(_14220_));
 AND2x2_ASAP7_75t_R _22491_ (.A(_14219_),
    .B(_14216_),
    .Y(_14221_));
 NAND2x1_ASAP7_75t_R _22492_ (.A(_00459_),
    .B(net6464),
    .Y(_14222_));
 OAI21x1_ASAP7_75t_R _22493_ (.A1(_14220_),
    .A2(_14221_),
    .B(_14222_),
    .Y(_14223_));
 XOR2x2_ASAP7_75t_R _22494_ (.A(_14223_),
    .B(net6507),
    .Y(_14224_));
 XOR2x2_ASAP7_75t_R _22496_ (.A(net6642),
    .B(net6614),
    .Y(_14225_));
 NAND2x1_ASAP7_75t_R _22497_ (.A(_11410_),
    .B(_14225_),
    .Y(_14226_));
 XNOR2x2_ASAP7_75t_R _22498_ (.A(net6642),
    .B(net6614),
    .Y(_14227_));
 NAND2x1_ASAP7_75t_R _22499_ (.A(net6559),
    .B(_14227_),
    .Y(_14228_));
 INVx1_ASAP7_75t_R _22500_ (.A(net6415),
    .Y(_14229_));
 AOI21x1_ASAP7_75t_R _22501_ (.A1(_14226_),
    .A2(_14228_),
    .B(_14229_),
    .Y(_14230_));
 XOR2x2_ASAP7_75t_R _22502_ (.A(net6614),
    .B(net6559),
    .Y(_14231_));
 NAND2x1_ASAP7_75t_R _22503_ (.A(net6642),
    .B(_14231_),
    .Y(_14232_));
 INVx1_ASAP7_75t_R _22504_ (.A(_00583_),
    .Y(_14233_));
 XNOR2x2_ASAP7_75t_R _22505_ (.A(net6614),
    .B(net6559),
    .Y(_14234_));
 NAND2x1_ASAP7_75t_R _22506_ (.A(_14233_),
    .B(_14234_),
    .Y(_14235_));
 AOI21x1_ASAP7_75t_R _22507_ (.A1(_14232_),
    .A2(_14235_),
    .B(net6415),
    .Y(_14236_));
 OAI21x1_ASAP7_75t_R _22508_ (.A1(_14230_),
    .A2(_14236_),
    .B(net6669),
    .Y(_14237_));
 NOR2x1_ASAP7_75t_R _22509_ (.A(net6670),
    .B(_00460_),
    .Y(_14238_));
 INVx1_ASAP7_75t_R _22510_ (.A(_14238_),
    .Y(_14239_));
 NAND3x1_ASAP7_75t_R _22511_ (.A(net6358),
    .B(_08764_),
    .C(net6387),
    .Y(_14240_));
 AO21x1_ASAP7_75t_R _22512_ (.A1(net6358),
    .A2(net6387),
    .B(_08764_),
    .Y(_14241_));
 NAND2x1_ASAP7_75t_R _22513_ (.A(_14240_),
    .B(_14241_),
    .Y(_14242_));
 NOR2x1_ASAP7_75t_R _22515_ (.A(net6669),
    .B(_00461_),
    .Y(_14243_));
 INVx1_ASAP7_75t_R _22516_ (.A(_14243_),
    .Y(_14244_));
 XOR2x2_ASAP7_75t_R _22517_ (.A(_11436_),
    .B(_00585_),
    .Y(_14245_));
 NOR2x1_ASAP7_75t_R _22518_ (.A(net6443),
    .B(_14245_),
    .Y(_14246_));
 INVx1_ASAP7_75t_R _22519_ (.A(net6443),
    .Y(_14247_));
 INVx1_ASAP7_75t_R _22520_ (.A(_00585_),
    .Y(_14248_));
 XOR2x2_ASAP7_75t_R _22521_ (.A(_11436_),
    .B(_14248_),
    .Y(_14249_));
 NOR2x1_ASAP7_75t_R _22522_ (.A(_14247_),
    .B(_14249_),
    .Y(_14250_));
 OAI21x1_ASAP7_75t_R _22523_ (.A1(_14246_),
    .A2(_14250_),
    .B(net6669),
    .Y(_14251_));
 AOI21x1_ASAP7_75t_R _22524_ (.A1(_14244_),
    .A2(net6357),
    .B(_08771_),
    .Y(_14252_));
 NAND2x1_ASAP7_75t_R _22525_ (.A(_00461_),
    .B(net6463),
    .Y(_14253_));
 NAND2x1_ASAP7_75t_R _22526_ (.A(_14247_),
    .B(_14249_),
    .Y(_14254_));
 NAND2x1_ASAP7_75t_R _22527_ (.A(_00585_),
    .B(_11432_),
    .Y(_14255_));
 NAND2x1_ASAP7_75t_R _22528_ (.A(_14248_),
    .B(_11436_),
    .Y(_14256_));
 AO21x1_ASAP7_75t_R _22529_ (.A1(_14255_),
    .A2(_14256_),
    .B(_14247_),
    .Y(_14257_));
 NAND3x1_ASAP7_75t_R _22530_ (.A(_14254_),
    .B(_14257_),
    .C(net6669),
    .Y(_14258_));
 AOI21x1_ASAP7_75t_R _22531_ (.A1(_14253_),
    .A2(_14258_),
    .B(net6506),
    .Y(_14259_));
 NOR2x2_ASAP7_75t_R _22532_ (.A(_14252_),
    .B(_14259_),
    .Y(_14260_));
 NAND3x1_ASAP7_75t_R _22534_ (.A(_14237_),
    .B(net6508),
    .C(_14239_),
    .Y(_14261_));
 AO21x1_ASAP7_75t_R _22535_ (.A1(_14237_),
    .A2(_14239_),
    .B(net6508),
    .Y(_14262_));
 NAND2x1p5_ASAP7_75t_R _22536_ (.A(_14261_),
    .B(_14262_),
    .Y(_14263_));
 AOI21x1_ASAP7_75t_R _22538_ (.A1(_14244_),
    .A2(_14251_),
    .B(net6506),
    .Y(_14264_));
 AOI21x1_ASAP7_75t_R _22539_ (.A1(_14253_),
    .A2(_14258_),
    .B(_08771_),
    .Y(_14265_));
 NOR2x1_ASAP7_75t_R _22540_ (.A(_14264_),
    .B(_14265_),
    .Y(_14266_));
 INVx1_ASAP7_75t_R _22543_ (.A(net6187),
    .Y(_14268_));
 NAND3x1_ASAP7_75t_R _22544_ (.A(net6357),
    .B(net6506),
    .C(_14244_),
    .Y(_14269_));
 AOI21x1_ASAP7_75t_R _22545_ (.A1(_14268_),
    .A2(_14269_),
    .B(net5289),
    .Y(_14270_));
 XOR2x2_ASAP7_75t_R _22547_ (.A(_08768_),
    .B(_14223_),
    .Y(_14272_));
 NOR2x1_ASAP7_75t_R _22548_ (.A(net5823),
    .B(net6185),
    .Y(_14273_));
 NOR2x1_ASAP7_75t_R _22549_ (.A(net5821),
    .B(_14273_),
    .Y(_14274_));
 XOR2x2_ASAP7_75t_R _22550_ (.A(_11471_),
    .B(_00586_),
    .Y(_14275_));
 XOR2x2_ASAP7_75t_R _22551_ (.A(net6589),
    .B(net6587),
    .Y(_14276_));
 XNOR2x2_ASAP7_75t_R _22552_ (.A(_14276_),
    .B(_11470_),
    .Y(_14277_));
 NOR2x1_ASAP7_75t_R _22553_ (.A(_14275_),
    .B(_14277_),
    .Y(_14278_));
 XNOR2x2_ASAP7_75t_R _22554_ (.A(_00586_),
    .B(_11471_),
    .Y(_14279_));
 XOR2x2_ASAP7_75t_R _22555_ (.A(_11470_),
    .B(_14276_),
    .Y(_14280_));
 NOR2x1_ASAP7_75t_R _22556_ (.A(_14279_),
    .B(_14280_),
    .Y(_14281_));
 OAI21x1_ASAP7_75t_R _22557_ (.A1(_14278_),
    .A2(_14281_),
    .B(net6669),
    .Y(_14282_));
 NOR2x1_ASAP7_75t_R _22558_ (.A(net6669),
    .B(_00499_),
    .Y(_14283_));
 INVx1_ASAP7_75t_R _22559_ (.A(_14283_),
    .Y(_14284_));
 NAND3x1_ASAP7_75t_R _22560_ (.A(_14282_),
    .B(_00880_),
    .C(_14284_),
    .Y(_14285_));
 AO21x1_ASAP7_75t_R _22561_ (.A1(_14282_),
    .A2(_14284_),
    .B(_00880_),
    .Y(_14286_));
 NAND2x1_ASAP7_75t_R _22562_ (.A(_14285_),
    .B(_14286_),
    .Y(_14287_));
 OAI21x1_ASAP7_75t_R _22565_ (.A1(_14270_),
    .A2(_14274_),
    .B(net5803),
    .Y(_14290_));
 NOR2x1_ASAP7_75t_R _22567_ (.A(net5290),
    .B(_14266_),
    .Y(_14292_));
 NOR2x1_ASAP7_75t_R _22569_ (.A(net6667),
    .B(_00498_),
    .Y(_14294_));
 XOR2x2_ASAP7_75t_R _22571_ (.A(_00587_),
    .B(_00651_),
    .Y(_14296_));
 XOR2x2_ASAP7_75t_R _22572_ (.A(_11482_),
    .B(_14296_),
    .Y(_14297_));
 XOR2x2_ASAP7_75t_R _22573_ (.A(_00650_),
    .B(net6587),
    .Y(_14298_));
 XOR2x2_ASAP7_75t_R _22574_ (.A(_14298_),
    .B(net6556),
    .Y(_14299_));
 XOR2x2_ASAP7_75t_R _22575_ (.A(_14297_),
    .B(_14299_),
    .Y(_14300_));
 NOR2x1_ASAP7_75t_R _22576_ (.A(net6463),
    .B(_14300_),
    .Y(_14301_));
 OAI21x1_ASAP7_75t_R _22577_ (.A1(_14294_),
    .A2(_14301_),
    .B(_00882_),
    .Y(_14302_));
 AND2x2_ASAP7_75t_R _22578_ (.A(net6463),
    .B(_00498_),
    .Y(_14303_));
 XNOR2x2_ASAP7_75t_R _22579_ (.A(_14299_),
    .B(_14297_),
    .Y(_14304_));
 NOR2x1_ASAP7_75t_R _22580_ (.A(net6463),
    .B(_14304_),
    .Y(_14305_));
 OAI21x1_ASAP7_75t_R _22581_ (.A1(_14303_),
    .A2(_14305_),
    .B(_08778_),
    .Y(_14306_));
 NAND2x1_ASAP7_75t_R _22582_ (.A(_14302_),
    .B(_14306_),
    .Y(_14307_));
 AO21x1_ASAP7_75t_R _22584_ (.A1(_14292_),
    .A2(net5803),
    .B(net5799),
    .Y(_14309_));
 NAND2x1_ASAP7_75t_R _22585_ (.A(net5822),
    .B(net5818),
    .Y(_14310_));
 OAI21x1_ASAP7_75t_R _22586_ (.A1(net6189),
    .A2(net6188),
    .B(_01168_),
    .Y(_14311_));
 AO21x1_ASAP7_75t_R _22587_ (.A1(net5462),
    .A2(net5167),
    .B(net5805),
    .Y(_14312_));
 INVx1_ASAP7_75t_R _22588_ (.A(_14312_),
    .Y(_14313_));
 NOR2x1_ASAP7_75t_R _22589_ (.A(_14309_),
    .B(_14313_),
    .Y(_14314_));
 NOR2x1_ASAP7_75t_R _22591_ (.A(_01182_),
    .B(net5804),
    .Y(_14316_));
 INVx1_ASAP7_75t_R _22592_ (.A(_01169_),
    .Y(_14317_));
 OAI21x1_ASAP7_75t_R _22593_ (.A1(net6187),
    .A2(net6186),
    .B(_14317_),
    .Y(_14318_));
 INVx2_ASAP7_75t_R _22594_ (.A(_14318_),
    .Y(_14319_));
 OAI21x1_ASAP7_75t_R _22596_ (.A1(_14294_),
    .A2(_14301_),
    .B(_08778_),
    .Y(_14321_));
 OAI21x1_ASAP7_75t_R _22597_ (.A1(_14303_),
    .A2(_14305_),
    .B(_00882_),
    .Y(_14322_));
 NAND2x1_ASAP7_75t_R _22598_ (.A(_14321_),
    .B(_14322_),
    .Y(_14323_));
 AO21x1_ASAP7_75t_R _22600_ (.A1(_14319_),
    .A2(net5806),
    .B(net5793),
    .Y(_14325_));
 NOR2x1_ASAP7_75t_R _22601_ (.A(net6667),
    .B(_00497_),
    .Y(_14326_));
 INVx1_ASAP7_75t_R _22602_ (.A(_14326_),
    .Y(_14327_));
 XNOR2x2_ASAP7_75t_R _22603_ (.A(_00588_),
    .B(_00619_),
    .Y(_14328_));
 INVx1_ASAP7_75t_R _22604_ (.A(_14328_),
    .Y(_14329_));
 XOR2x2_ASAP7_75t_R _22605_ (.A(_00651_),
    .B(net6588),
    .Y(_14330_));
 XOR2x2_ASAP7_75t_R _22606_ (.A(_14330_),
    .B(net6555),
    .Y(_14331_));
 NOR2x1_ASAP7_75t_R _22607_ (.A(_14329_),
    .B(_14331_),
    .Y(_14332_));
 XOR2x2_ASAP7_75t_R _22608_ (.A(_14330_),
    .B(_11508_),
    .Y(_14333_));
 NOR2x1_ASAP7_75t_R _22609_ (.A(_14328_),
    .B(_14333_),
    .Y(_14334_));
 OAI21x1_ASAP7_75t_R _22610_ (.A1(_14332_),
    .A2(_14334_),
    .B(net6667),
    .Y(_14335_));
 AOI21x1_ASAP7_75t_R _22611_ (.A1(_14327_),
    .A2(_14335_),
    .B(_00883_),
    .Y(_14336_));
 AND3x1_ASAP7_75t_R _22612_ (.A(_14335_),
    .B(_00883_),
    .C(_14327_),
    .Y(_14337_));
 NOR2x1_ASAP7_75t_R _22613_ (.A(_14336_),
    .B(_14337_),
    .Y(_14338_));
 INVx1_ASAP7_75t_R _22614_ (.A(_14338_),
    .Y(_14339_));
 OAI21x1_ASAP7_75t_R _22616_ (.A1(_14316_),
    .A2(_14325_),
    .B(net5461),
    .Y(_14341_));
 AOI21x1_ASAP7_75t_R _22617_ (.A1(_14290_),
    .A2(_14314_),
    .B(_14341_),
    .Y(_14342_));
 INVx1_ASAP7_75t_R _22618_ (.A(net5287),
    .Y(_14343_));
 NAND3x1_ASAP7_75t_R _22619_ (.A(_14282_),
    .B(_08775_),
    .C(_14284_),
    .Y(_14344_));
 AO21x1_ASAP7_75t_R _22620_ (.A1(_14282_),
    .A2(_14284_),
    .B(_08775_),
    .Y(_14345_));
 NAND2x1_ASAP7_75t_R _22621_ (.A(_14344_),
    .B(_14345_),
    .Y(_14346_));
 OAI21x1_ASAP7_75t_R _22622_ (.A1(_14343_),
    .A2(net5816),
    .B(net5791),
    .Y(_14347_));
 NAND2x1_ASAP7_75t_R _22623_ (.A(net5817),
    .B(net6191),
    .Y(_14348_));
 NOR2x1_ASAP7_75t_R _22624_ (.A(net5821),
    .B(_14348_),
    .Y(_14349_));
 NOR2x1_ASAP7_75t_R _22625_ (.A(_14347_),
    .B(_14349_),
    .Y(_14350_));
 NOR2x1_ASAP7_75t_R _22626_ (.A(net5290),
    .B(net5821),
    .Y(_14351_));
 AO21x1_ASAP7_75t_R _22628_ (.A1(_14351_),
    .A2(net5804),
    .B(net5799),
    .Y(_14353_));
 OAI21x1_ASAP7_75t_R _22630_ (.A1(_14350_),
    .A2(_14353_),
    .B(net5792),
    .Y(_14355_));
 OAI21x1_ASAP7_75t_R _22632_ (.A1(net5288),
    .A2(net5812),
    .B(net5808),
    .Y(_14357_));
 NAND2x1_ASAP7_75t_R _22635_ (.A(net5785),
    .B(_14351_),
    .Y(_14360_));
 OAI21x1_ASAP7_75t_R _22636_ (.A1(_14349_),
    .A2(_14357_),
    .B(_14360_),
    .Y(_14361_));
 NOR2x1_ASAP7_75t_R _22637_ (.A(net5793),
    .B(_14361_),
    .Y(_14362_));
 XOR2x2_ASAP7_75t_R _22638_ (.A(_00653_),
    .B(_00685_),
    .Y(_14363_));
 XOR2x2_ASAP7_75t_R _22639_ (.A(_11504_),
    .B(_00589_),
    .Y(_14364_));
 XNOR2x2_ASAP7_75t_R _22640_ (.A(_14363_),
    .B(_14364_),
    .Y(_14365_));
 NOR2x1_ASAP7_75t_R _22641_ (.A(net6667),
    .B(_00496_),
    .Y(_14366_));
 AO21x1_ASAP7_75t_R _22642_ (.A1(_14365_),
    .A2(net6667),
    .B(_14366_),
    .Y(_14367_));
 XOR2x2_ASAP7_75t_R _22643_ (.A(_14367_),
    .B(_00884_),
    .Y(_14368_));
 OAI21x1_ASAP7_75t_R _22645_ (.A1(_14355_),
    .A2(_14362_),
    .B(net6181),
    .Y(_14370_));
 NOR2x1_ASAP7_75t_R _22646_ (.A(_14342_),
    .B(_14370_),
    .Y(_14371_));
 NAND3x1_ASAP7_75t_R _22647_ (.A(net6357),
    .B(_08771_),
    .C(_14244_),
    .Y(_14372_));
 INVx1_ASAP7_75t_R _22648_ (.A(_14252_),
    .Y(_14373_));
 AO21x1_ASAP7_75t_R _22649_ (.A1(_14372_),
    .A2(_14373_),
    .B(net5290),
    .Y(_14374_));
 NAND2x1_ASAP7_75t_R _22650_ (.A(_01168_),
    .B(net5818),
    .Y(_14375_));
 AOI21x1_ASAP7_75t_R _22653_ (.A1(_14374_),
    .A2(_14375_),
    .B(net5791),
    .Y(_14378_));
 INVx1_ASAP7_75t_R _22655_ (.A(_01172_),
    .Y(_14380_));
 NOR2x1_ASAP7_75t_R _22656_ (.A(_14380_),
    .B(net5821),
    .Y(_14381_));
 OAI21x1_ASAP7_75t_R _22658_ (.A1(net5803),
    .A2(_14381_),
    .B(net5799),
    .Y(_14383_));
 OAI21x1_ASAP7_75t_R _22659_ (.A1(_14378_),
    .A2(_14383_),
    .B(net5792),
    .Y(_14384_));
 INVx1_ASAP7_75t_R _22660_ (.A(_01174_),
    .Y(_14385_));
 AO21x1_ASAP7_75t_R _22661_ (.A1(_14269_),
    .A2(_14268_),
    .B(_14385_),
    .Y(_14386_));
 NAND2x1_ASAP7_75t_R _22663_ (.A(net5822),
    .B(net5813),
    .Y(_14388_));
 AOI21x1_ASAP7_75t_R _22664_ (.A1(net4913),
    .A2(net5458),
    .B(net5805),
    .Y(_14389_));
 OAI21x1_ASAP7_75t_R _22666_ (.A1(net6184),
    .A2(net5821),
    .B(net4760),
    .Y(_14390_));
 OAI21x1_ASAP7_75t_R _22667_ (.A1(_14390_),
    .A2(net5785),
    .B(net5793),
    .Y(_14391_));
 NOR2x1_ASAP7_75t_R _22668_ (.A(_14389_),
    .B(_14391_),
    .Y(_14392_));
 INVx1_ASAP7_75t_R _22669_ (.A(_14368_),
    .Y(_14393_));
 OAI21x1_ASAP7_75t_R _22672_ (.A1(_14384_),
    .A2(_14392_),
    .B(net5782),
    .Y(_14396_));
 OAI21x1_ASAP7_75t_R _22673_ (.A1(net6185),
    .A2(net5817),
    .B(net5813),
    .Y(_14397_));
 AOI21x1_ASAP7_75t_R _22674_ (.A1(_14310_),
    .A2(_14397_),
    .B(net5808),
    .Y(_14398_));
 INVx1_ASAP7_75t_R _22675_ (.A(_14398_),
    .Y(_14399_));
 AOI21x1_ASAP7_75t_R _22676_ (.A1(net5806),
    .A2(_14270_),
    .B(net5800),
    .Y(_14400_));
 AO21x1_ASAP7_75t_R _22677_ (.A1(_14270_),
    .A2(net5806),
    .B(net5797),
    .Y(_14401_));
 AOI21x1_ASAP7_75t_R _22679_ (.A1(_14373_),
    .A2(_14372_),
    .B(_14317_),
    .Y(_14403_));
 AOI21x1_ASAP7_75t_R _22680_ (.A1(_14373_),
    .A2(_14372_),
    .B(net5287),
    .Y(_14404_));
 NAND2x1_ASAP7_75t_R _22681_ (.A(net5810),
    .B(net5164),
    .Y(_14405_));
 OAI21x1_ASAP7_75t_R _22682_ (.A1(net5806),
    .A2(net4758),
    .B(net4910),
    .Y(_14406_));
 OAI21x1_ASAP7_75t_R _22683_ (.A1(net4911),
    .A2(_14406_),
    .B(net5461),
    .Y(_14407_));
 AOI21x1_ASAP7_75t_R _22684_ (.A1(net4912),
    .A2(_14400_),
    .B(_14407_),
    .Y(_14408_));
 XOR2x2_ASAP7_75t_R _22685_ (.A(_00653_),
    .B(net6587),
    .Y(_14409_));
 XOR2x2_ASAP7_75t_R _22686_ (.A(_14409_),
    .B(net6440),
    .Y(_14410_));
 XOR2x2_ASAP7_75t_R _22687_ (.A(net6640),
    .B(_00621_),
    .Y(_14411_));
 XOR2x2_ASAP7_75t_R _22688_ (.A(_14410_),
    .B(_14411_),
    .Y(_14412_));
 NOR2x1_ASAP7_75t_R _22689_ (.A(net6667),
    .B(_00495_),
    .Y(_14413_));
 AO21x1_ASAP7_75t_R _22690_ (.A1(_14412_),
    .A2(net6667),
    .B(_14413_),
    .Y(_14414_));
 XOR2x2_ASAP7_75t_R _22691_ (.A(_14414_),
    .B(net6504),
    .Y(_14415_));
 INVx1_ASAP7_75t_R _22692_ (.A(_14415_),
    .Y(_14416_));
 OAI21x1_ASAP7_75t_R _22693_ (.A1(_14396_),
    .A2(_14408_),
    .B(_14416_),
    .Y(_14417_));
 AO21x1_ASAP7_75t_R _22694_ (.A1(_14372_),
    .A2(_14373_),
    .B(net5286),
    .Y(_14418_));
 AOI21x1_ASAP7_75t_R _22695_ (.A1(_14418_),
    .A2(net5462),
    .B(net5809),
    .Y(_14419_));
 NAND2x1_ASAP7_75t_R _22696_ (.A(net6190),
    .B(net5813),
    .Y(_14420_));
 OAI21x1_ASAP7_75t_R _22697_ (.A1(net6185),
    .A2(net5822),
    .B(net5818),
    .Y(_14421_));
 AOI21x1_ASAP7_75t_R _22699_ (.A1(_14420_),
    .A2(_14421_),
    .B(net5783),
    .Y(_14423_));
 OAI21x1_ASAP7_75t_R _22701_ (.A1(_14419_),
    .A2(_14423_),
    .B(net5800),
    .Y(_14425_));
 NAND2x1_ASAP7_75t_R _22702_ (.A(net6185),
    .B(net5818),
    .Y(_14426_));
 AOI21x1_ASAP7_75t_R _22704_ (.A1(_14374_),
    .A2(_14426_),
    .B(net5791),
    .Y(_14428_));
 OAI21x1_ASAP7_75t_R _22707_ (.A1(_14428_),
    .A2(_14398_),
    .B(net5797),
    .Y(_14431_));
 AOI21x1_ASAP7_75t_R _22710_ (.A1(_14425_),
    .A2(_14431_),
    .B(net5792),
    .Y(_14434_));
 NOR2x1_ASAP7_75t_R _22711_ (.A(net5822),
    .B(net5811),
    .Y(_14435_));
 OAI21x1_ASAP7_75t_R _22712_ (.A1(net5784),
    .A2(_14435_),
    .B(net5794),
    .Y(_14436_));
 AO21x1_ASAP7_75t_R _22713_ (.A1(_14372_),
    .A2(_14373_),
    .B(net5289),
    .Y(_14437_));
 AOI21x1_ASAP7_75t_R _22714_ (.A1(_14437_),
    .A2(_14421_),
    .B(net5808),
    .Y(_14438_));
 OAI21x1_ASAP7_75t_R _22715_ (.A1(_14436_),
    .A2(_14438_),
    .B(net5792),
    .Y(_14439_));
 INVx1_ASAP7_75t_R _22716_ (.A(_01177_),
    .Y(_14440_));
 OAI21x1_ASAP7_75t_R _22717_ (.A1(net5162),
    .A2(net5812),
    .B(net5791),
    .Y(_14441_));
 OAI21x1_ASAP7_75t_R _22718_ (.A1(net4758),
    .A2(net4909),
    .B(net5800),
    .Y(_14442_));
 NOR2x1_ASAP7_75t_R _22719_ (.A(net5822),
    .B(net5818),
    .Y(_14443_));
 OAI21x1_ASAP7_75t_R _22720_ (.A1(net5814),
    .A2(_14348_),
    .B(net5802),
    .Y(_14444_));
 NOR2x1_ASAP7_75t_R _22721_ (.A(_14443_),
    .B(_14444_),
    .Y(_14445_));
 NOR2x1_ASAP7_75t_R _22722_ (.A(_14442_),
    .B(_14445_),
    .Y(_14446_));
 OAI21x1_ASAP7_75t_R _22723_ (.A1(_14439_),
    .A2(_14446_),
    .B(net5780),
    .Y(_14447_));
 OAI21x1_ASAP7_75t_R _22724_ (.A1(_14434_),
    .A2(_14447_),
    .B(net6180),
    .Y(_14448_));
 AO21x1_ASAP7_75t_R _22725_ (.A1(_14372_),
    .A2(_14373_),
    .B(net5257),
    .Y(_14449_));
 OAI21x1_ASAP7_75t_R _22726_ (.A1(net6185),
    .A2(net5817),
    .B(net5818),
    .Y(_14450_));
 AOI21x1_ASAP7_75t_R _22728_ (.A1(net5008),
    .A2(_14450_),
    .B(net5783),
    .Y(_14452_));
 NOR2x1_ASAP7_75t_R _22729_ (.A(net5165),
    .B(net5818),
    .Y(_14453_));
 INVx1_ASAP7_75t_R _22730_ (.A(_14453_),
    .Y(_14454_));
 AOI21x1_ASAP7_75t_R _22731_ (.A1(_14375_),
    .A2(net4679),
    .B(net5809),
    .Y(_14455_));
 OAI21x1_ASAP7_75t_R _22734_ (.A1(_14452_),
    .A2(_14455_),
    .B(net5797),
    .Y(_14458_));
 NAND2x1_ASAP7_75t_R _22735_ (.A(net5817),
    .B(net6184),
    .Y(_14459_));
 AOI21x1_ASAP7_75t_R _22736_ (.A1(_14459_),
    .A2(net5457),
    .B(net5805),
    .Y(_14460_));
 NOR2x1_ASAP7_75t_R _22737_ (.A(net5817),
    .B(net5813),
    .Y(_14461_));
 OAI21x1_ASAP7_75t_R _22738_ (.A1(_14273_),
    .A2(_14461_),
    .B(net5809),
    .Y(_14462_));
 INVx1_ASAP7_75t_R _22739_ (.A(_14462_),
    .Y(_14463_));
 OAI21x1_ASAP7_75t_R _22741_ (.A1(_14460_),
    .A2(_14463_),
    .B(net5800),
    .Y(_14465_));
 AOI21x1_ASAP7_75t_R _22743_ (.A1(_14458_),
    .A2(_14465_),
    .B(net5461),
    .Y(_14467_));
 NOR2x1p5_ASAP7_75t_R _22744_ (.A(_14403_),
    .B(net5809),
    .Y(_14468_));
 NOR2x1_ASAP7_75t_R _22745_ (.A(_01168_),
    .B(net5811),
    .Y(_14469_));
 INVx1_ASAP7_75t_R _22746_ (.A(_14469_),
    .Y(_14470_));
 AOI21x1_ASAP7_75t_R _22747_ (.A1(net5167),
    .A2(net4913),
    .B(net5787),
    .Y(_14471_));
 AOI211x1_ASAP7_75t_R _22748_ (.A1(_14470_),
    .A2(_14468_),
    .B(_14471_),
    .C(net5800),
    .Y(_14472_));
 OAI21x1_ASAP7_75t_R _22750_ (.A1(net6189),
    .A2(net6188),
    .B(net5257),
    .Y(_14474_));
 OAI21x1_ASAP7_75t_R _22751_ (.A1(net6190),
    .A2(net5812),
    .B(net5006),
    .Y(_14475_));
 OAI21x1_ASAP7_75t_R _22752_ (.A1(net6187),
    .A2(net6186),
    .B(net5257),
    .Y(_14476_));
 INVx1_ASAP7_75t_R _22753_ (.A(_14476_),
    .Y(_14477_));
 NAND2x1_ASAP7_75t_R _22754_ (.A(net5789),
    .B(_14477_),
    .Y(_14478_));
 OAI21x1_ASAP7_75t_R _22755_ (.A1(net5787),
    .A2(_14475_),
    .B(_14478_),
    .Y(_14479_));
 OAI21x1_ASAP7_75t_R _22756_ (.A1(net5795),
    .A2(_14479_),
    .B(net5461),
    .Y(_14480_));
 OAI21x1_ASAP7_75t_R _22757_ (.A1(_14480_),
    .A2(_14472_),
    .B(net6181),
    .Y(_14481_));
 NOR2x1_ASAP7_75t_R _22758_ (.A(_14467_),
    .B(_14481_),
    .Y(_14482_));
 OAI22x1_ASAP7_75t_R _22759_ (.A1(_14371_),
    .A2(_14417_),
    .B1(_14482_),
    .B2(_14448_),
    .Y(_00072_));
 NOR2x1_ASAP7_75t_R _22760_ (.A(net6191),
    .B(net5814),
    .Y(_14483_));
 AO21x1_ASAP7_75t_R _22761_ (.A1(net5289),
    .A2(net5814),
    .B(net5801),
    .Y(_14484_));
 NOR2x1_ASAP7_75t_R _22762_ (.A(_14483_),
    .B(_14484_),
    .Y(_14485_));
 NAND2x1_ASAP7_75t_R _22764_ (.A(net5817),
    .B(net5814),
    .Y(_14487_));
 AOI21x1_ASAP7_75t_R _22766_ (.A1(_14487_),
    .A2(_14426_),
    .B(net5785),
    .Y(_14489_));
 NOR3x1_ASAP7_75t_R _22767_ (.A(_14485_),
    .B(net5792),
    .C(_14489_),
    .Y(_14490_));
 OAI21x1_ASAP7_75t_R _22768_ (.A1(_01168_),
    .A2(net5811),
    .B(net5807),
    .Y(_14491_));
 OA21x2_ASAP7_75t_R _22769_ (.A1(_14491_),
    .A2(_14443_),
    .B(net5792),
    .Y(_14492_));
 AO21x1_ASAP7_75t_R _22770_ (.A1(_14397_),
    .A2(_14421_),
    .B(net5808),
    .Y(_14493_));
 AO21x1_ASAP7_75t_R _22771_ (.A1(_14492_),
    .A2(_14493_),
    .B(net5780),
    .Y(_14494_));
 NOR2x1_ASAP7_75t_R _22772_ (.A(_14490_),
    .B(_14494_),
    .Y(_14495_));
 AOI21x1_ASAP7_75t_R _22773_ (.A1(net6190),
    .A2(net5823),
    .B(net5816),
    .Y(_14496_));
 OAI21x1_ASAP7_75t_R _22774_ (.A1(net4758),
    .A2(_14496_),
    .B(net5787),
    .Y(_14497_));
 INVx1_ASAP7_75t_R _22775_ (.A(_14497_),
    .Y(_14498_));
 INVx1_ASAP7_75t_R _22776_ (.A(net5290),
    .Y(_14499_));
 NOR2x1_ASAP7_75t_R _22777_ (.A(_14499_),
    .B(net5814),
    .Y(_14500_));
 AO21x1_ASAP7_75t_R _22778_ (.A1(_14372_),
    .A2(_14373_),
    .B(_14440_),
    .Y(_14501_));
 NAND2x1_ASAP7_75t_R _22779_ (.A(net5804),
    .B(_14501_),
    .Y(_14502_));
 OAI21x1_ASAP7_75t_R _22780_ (.A1(_14500_),
    .A2(_14502_),
    .B(net5461),
    .Y(_14503_));
 OAI21x1_ASAP7_75t_R _22781_ (.A1(_14498_),
    .A2(_14503_),
    .B(net5780),
    .Y(_14504_));
 INVx1_ASAP7_75t_R _22782_ (.A(_14311_),
    .Y(_14505_));
 AO21x1_ASAP7_75t_R _22784_ (.A1(_14351_),
    .A2(net5804),
    .B(net5461),
    .Y(_14507_));
 NAND2x1_ASAP7_75t_R _22785_ (.A(net5787),
    .B(_14319_),
    .Y(_14508_));
 OAI21x1_ASAP7_75t_R _22786_ (.A1(net5787),
    .A2(net5462),
    .B(_14508_),
    .Y(_14509_));
 AOI211x1_ASAP7_75t_R _22787_ (.A1(net5789),
    .A2(_14505_),
    .B(_14507_),
    .C(_14509_),
    .Y(_14510_));
 OAI21x1_ASAP7_75t_R _22788_ (.A1(_14504_),
    .A2(_14510_),
    .B(net5800),
    .Y(_14511_));
 NOR2x1_ASAP7_75t_R _22789_ (.A(_14495_),
    .B(_14511_),
    .Y(_14512_));
 AO21x1_ASAP7_75t_R _22790_ (.A1(net5822),
    .A2(net5811),
    .B(net5784),
    .Y(_14513_));
 OAI21x1_ASAP7_75t_R _22791_ (.A1(_14469_),
    .A2(_14513_),
    .B(net5792),
    .Y(_14514_));
 NAND2x1_ASAP7_75t_R _22792_ (.A(net5822),
    .B(net6190),
    .Y(_14515_));
 NOR2x1_ASAP7_75t_R _22793_ (.A(net5819),
    .B(_14515_),
    .Y(_14516_));
 AO21x1_ASAP7_75t_R _22794_ (.A1(net5817),
    .A2(net5820),
    .B(net5791),
    .Y(_14517_));
 AOI21x1_ASAP7_75t_R _22795_ (.A1(net5786),
    .A2(net5007),
    .B(net5792),
    .Y(_14518_));
 OAI21x1_ASAP7_75t_R _22796_ (.A1(_14516_),
    .A2(net5455),
    .B(_14518_),
    .Y(_14519_));
 OAI21x1_ASAP7_75t_R _22797_ (.A1(_14485_),
    .A2(_14514_),
    .B(_14519_),
    .Y(_14520_));
 NAND2x1_ASAP7_75t_R _22798_ (.A(_14386_),
    .B(_14397_),
    .Y(_14521_));
 INVx1_ASAP7_75t_R _22799_ (.A(_01184_),
    .Y(_14522_));
 NOR2x1_ASAP7_75t_R _22800_ (.A(_14522_),
    .B(net5792),
    .Y(_14523_));
 AO21x1_ASAP7_75t_R _22801_ (.A1(_14523_),
    .A2(net5784),
    .B(net5780),
    .Y(_14524_));
 AOI21x1_ASAP7_75t_R _22802_ (.A1(net5801),
    .A2(net4678),
    .B(_14524_),
    .Y(_14525_));
 AOI21x1_ASAP7_75t_R _22803_ (.A1(net5780),
    .A2(_14520_),
    .B(_14525_),
    .Y(_14526_));
 OAI21x1_ASAP7_75t_R _22804_ (.A1(net5798),
    .A2(_14526_),
    .B(net6180),
    .Y(_14527_));
 OAI21x1_ASAP7_75t_R _22805_ (.A1(net6187),
    .A2(net6186),
    .B(_14380_),
    .Y(_14528_));
 AO21x1_ASAP7_75t_R _22806_ (.A1(_14528_),
    .A2(net5006),
    .B(net5805),
    .Y(_14529_));
 OAI21x1_ASAP7_75t_R _22807_ (.A1(_14505_),
    .A2(_14461_),
    .B(net5805),
    .Y(_14530_));
 AOI21x1_ASAP7_75t_R _22808_ (.A1(_14529_),
    .A2(_14530_),
    .B(net5795),
    .Y(_14531_));
 NOR2x1_ASAP7_75t_R _22809_ (.A(net5817),
    .B(net6185),
    .Y(_14532_));
 OAI21x1_ASAP7_75t_R _22811_ (.A1(_14532_),
    .A2(_14443_),
    .B(net5784),
    .Y(_14534_));
 NOR2x1_ASAP7_75t_R _22812_ (.A(net5817),
    .B(net5818),
    .Y(_14535_));
 OAI21x1_ASAP7_75t_R _22813_ (.A1(_14477_),
    .A2(_14535_),
    .B(net5805),
    .Y(_14536_));
 AOI21x1_ASAP7_75t_R _22814_ (.A1(_14534_),
    .A2(_14536_),
    .B(net5800),
    .Y(_14537_));
 OAI21x1_ASAP7_75t_R _22815_ (.A1(_14531_),
    .A2(_14537_),
    .B(net5461),
    .Y(_14538_));
 AOI21x1_ASAP7_75t_R _22816_ (.A1(net6190),
    .A2(net5823),
    .B(net5818),
    .Y(_14539_));
 NAND2x1_ASAP7_75t_R _22817_ (.A(net5809),
    .B(_14539_),
    .Y(_14540_));
 NAND2x1_ASAP7_75t_R _22818_ (.A(net6184),
    .B(_14266_),
    .Y(_14541_));
 INVx1_ASAP7_75t_R _22820_ (.A(_14441_),
    .Y(_14543_));
 AOI21x1_ASAP7_75t_R _22821_ (.A1(net5453),
    .A2(_14543_),
    .B(net5797),
    .Y(_14544_));
 NAND2x1_ASAP7_75t_R _22822_ (.A(_14540_),
    .B(_14544_),
    .Y(_14545_));
 OA21x2_ASAP7_75t_R _22823_ (.A1(_14437_),
    .A2(net5791),
    .B(net5797),
    .Y(_14546_));
 AOI21x1_ASAP7_75t_R _22824_ (.A1(_14497_),
    .A2(_14546_),
    .B(net5461),
    .Y(_14547_));
 AOI21x1_ASAP7_75t_R _22825_ (.A1(_14545_),
    .A2(_14547_),
    .B(net6181),
    .Y(_14548_));
 NAND2x1_ASAP7_75t_R _22826_ (.A(_14538_),
    .B(_14548_),
    .Y(_14549_));
 NAND2x1_ASAP7_75t_R _22827_ (.A(net6191),
    .B(net5818),
    .Y(_14550_));
 AOI21x1_ASAP7_75t_R _22828_ (.A1(net5785),
    .A2(_14550_),
    .B(net5793),
    .Y(_14551_));
 OA21x2_ASAP7_75t_R _22829_ (.A1(net5788),
    .A2(_14528_),
    .B(_14541_),
    .Y(_14552_));
 AOI21x1_ASAP7_75t_R _22830_ (.A1(_14551_),
    .A2(_14552_),
    .B(net5792),
    .Y(_14553_));
 NAND2x1_ASAP7_75t_R _22831_ (.A(net5790),
    .B(_14476_),
    .Y(_14554_));
 INVx1_ASAP7_75t_R _22832_ (.A(_14501_),
    .Y(_14555_));
 OA21x2_ASAP7_75t_R _22833_ (.A1(_14554_),
    .A2(_14555_),
    .B(net5793),
    .Y(_14556_));
 NAND2x1_ASAP7_75t_R _22834_ (.A(_14290_),
    .B(_14556_),
    .Y(_14557_));
 NAND2x1_ASAP7_75t_R _22835_ (.A(_14553_),
    .B(_14557_),
    .Y(_14558_));
 NAND2x1_ASAP7_75t_R _22836_ (.A(net5817),
    .B(net5819),
    .Y(_14559_));
 AOI21x1_ASAP7_75t_R _22837_ (.A1(_14559_),
    .A2(_14468_),
    .B(net5797),
    .Y(_14560_));
 AO21x1_ASAP7_75t_R _22838_ (.A1(_14559_),
    .A2(_14437_),
    .B(net5791),
    .Y(_14561_));
 NAND2x1_ASAP7_75t_R _22839_ (.A(_14561_),
    .B(_14560_),
    .Y(_14562_));
 NOR2x1_ASAP7_75t_R _22840_ (.A(net5817),
    .B(net6190),
    .Y(_14563_));
 NOR2x1_ASAP7_75t_R _22841_ (.A(net6184),
    .B(net5815),
    .Y(_14564_));
 OAI21x1_ASAP7_75t_R _22842_ (.A1(_14563_),
    .A2(_14564_),
    .B(net5803),
    .Y(_14565_));
 NOR2x1_ASAP7_75t_R _22843_ (.A(net5814),
    .B(net5801),
    .Y(_14566_));
 AOI21x1_ASAP7_75t_R _22844_ (.A1(net5459),
    .A2(_14566_),
    .B(net5799),
    .Y(_14567_));
 AOI21x1_ASAP7_75t_R _22845_ (.A1(_14565_),
    .A2(_14567_),
    .B(net5461),
    .Y(_14568_));
 AOI21x1_ASAP7_75t_R _22846_ (.A1(_14562_),
    .A2(_14568_),
    .B(net5780),
    .Y(_14569_));
 AOI21x1_ASAP7_75t_R _22847_ (.A1(_14558_),
    .A2(_14569_),
    .B(net6180),
    .Y(_14570_));
 NAND2x1_ASAP7_75t_R _22848_ (.A(_14549_),
    .B(_14570_),
    .Y(_14571_));
 OAI21x1_ASAP7_75t_R _22849_ (.A1(_14512_),
    .A2(_14527_),
    .B(_14571_),
    .Y(_00073_));
 OAI21x1_ASAP7_75t_R _22850_ (.A1(net4758),
    .A2(_14564_),
    .B(net5806),
    .Y(_14572_));
 AO21x1_ASAP7_75t_R _22851_ (.A1(_14269_),
    .A2(_14268_),
    .B(net5290),
    .Y(_14573_));
 NAND3x1_ASAP7_75t_R _22852_ (.A(net5457),
    .B(_14573_),
    .C(net5787),
    .Y(_14574_));
 AOI21x1_ASAP7_75t_R _22853_ (.A1(_14572_),
    .A2(_14574_),
    .B(net5795),
    .Y(_14575_));
 AOI21x1_ASAP7_75t_R _22854_ (.A1(_14418_),
    .A2(_14450_),
    .B(net5809),
    .Y(_14576_));
 NAND2x1_ASAP7_75t_R _22855_ (.A(net5794),
    .B(_14444_),
    .Y(_14577_));
 OAI21x1_ASAP7_75t_R _22856_ (.A1(_14576_),
    .A2(_14577_),
    .B(net5792),
    .Y(_14578_));
 OAI21x1_ASAP7_75t_R _22857_ (.A1(_14575_),
    .A2(_14578_),
    .B(net6181),
    .Y(_14579_));
 AO21x1_ASAP7_75t_R _22858_ (.A1(_14269_),
    .A2(_14268_),
    .B(net5286),
    .Y(_14580_));
 AOI21x1_ASAP7_75t_R _22859_ (.A1(_14580_),
    .A2(_14437_),
    .B(net5788),
    .Y(_14581_));
 AOI21x1_ASAP7_75t_R _22860_ (.A1(net5454),
    .A2(_14421_),
    .B(net5803),
    .Y(_14582_));
 OAI21x1_ASAP7_75t_R _22861_ (.A1(_14581_),
    .A2(_14582_),
    .B(net5799),
    .Y(_14583_));
 NAND2x1_ASAP7_75t_R _22862_ (.A(net5791),
    .B(_14528_),
    .Y(_14584_));
 NOR2x1_ASAP7_75t_R _22863_ (.A(_14584_),
    .B(_14274_),
    .Y(_14585_));
 OR2x2_ASAP7_75t_R _22864_ (.A(_14391_),
    .B(_14585_),
    .Y(_14586_));
 AOI21x1_ASAP7_75t_R _22865_ (.A1(_14583_),
    .A2(_14586_),
    .B(net5792),
    .Y(_14587_));
 NOR2x1_ASAP7_75t_R _22866_ (.A(_14579_),
    .B(_14587_),
    .Y(_14588_));
 INVx1_ASAP7_75t_R _22867_ (.A(_14404_),
    .Y(_14589_));
 AOI21x1_ASAP7_75t_R _22868_ (.A1(net4905),
    .A2(_14426_),
    .B(net5805),
    .Y(_14590_));
 AOI21x1_ASAP7_75t_R _22869_ (.A1(net5161),
    .A2(net5458),
    .B(net5790),
    .Y(_14591_));
 OAI21x1_ASAP7_75t_R _22870_ (.A1(_14590_),
    .A2(_14591_),
    .B(net5799),
    .Y(_14592_));
 AO21x1_ASAP7_75t_R _22871_ (.A1(_14269_),
    .A2(_14268_),
    .B(net5287),
    .Y(_14593_));
 AOI21x1_ASAP7_75t_R _22872_ (.A1(_14593_),
    .A2(net5457),
    .B(net5787),
    .Y(_14594_));
 AND3x1_ASAP7_75t_R _22873_ (.A(net4760),
    .B(net5006),
    .C(net5790),
    .Y(_14595_));
 OAI21x1_ASAP7_75t_R _22874_ (.A1(_14594_),
    .A2(_14595_),
    .B(net5796),
    .Y(_14596_));
 AOI21x1_ASAP7_75t_R _22875_ (.A1(_14592_),
    .A2(_14596_),
    .B(net5461),
    .Y(_14597_));
 AOI21x1_ASAP7_75t_R _22876_ (.A1(net4906),
    .A2(_14420_),
    .B(net5810),
    .Y(_14598_));
 NAND2x1_ASAP7_75t_R _22877_ (.A(_14405_),
    .B(_14400_),
    .Y(_14599_));
 OAI21x1_ASAP7_75t_R _22878_ (.A1(_14598_),
    .A2(_14599_),
    .B(net5461),
    .Y(_14600_));
 OA21x2_ASAP7_75t_R _22879_ (.A1(_14535_),
    .A2(_14270_),
    .B(net5789),
    .Y(_14601_));
 AOI21x1_ASAP7_75t_R _22880_ (.A1(net5806),
    .A2(net5163),
    .B(net5797),
    .Y(_14602_));
 OAI21x1_ASAP7_75t_R _22881_ (.A1(net5789),
    .A2(net5161),
    .B(_14602_),
    .Y(_14603_));
 NOR2x1_ASAP7_75t_R _22882_ (.A(_14601_),
    .B(_14603_),
    .Y(_14604_));
 OAI21x1_ASAP7_75t_R _22883_ (.A1(_14600_),
    .A2(_14604_),
    .B(net5782),
    .Y(_14605_));
 OAI21x1_ASAP7_75t_R _22884_ (.A1(_14597_),
    .A2(_14605_),
    .B(net6180),
    .Y(_14606_));
 OAI21x1_ASAP7_75t_R _22885_ (.A1(net5785),
    .A2(_14390_),
    .B(net5799),
    .Y(_14607_));
 OA21x2_ASAP7_75t_R _22886_ (.A1(_14535_),
    .A2(_14564_),
    .B(net5785),
    .Y(_14608_));
 NOR2x1_ASAP7_75t_R _22887_ (.A(_14607_),
    .B(_14608_),
    .Y(_14609_));
 OAI21x1_ASAP7_75t_R _22888_ (.A1(_01182_),
    .A2(net5785),
    .B(net5793),
    .Y(_14610_));
 NOR2x1_ASAP7_75t_R _22889_ (.A(net4756),
    .B(_14349_),
    .Y(_14611_));
 OAI21x1_ASAP7_75t_R _22890_ (.A1(_14610_),
    .A2(_14611_),
    .B(net5792),
    .Y(_14612_));
 OAI21x1_ASAP7_75t_R _22891_ (.A1(_14609_),
    .A2(_14612_),
    .B(_14393_),
    .Y(_14613_));
 NOR2x1_ASAP7_75t_R _22892_ (.A(_14522_),
    .B(net5784),
    .Y(_14614_));
 NOR2x1_ASAP7_75t_R _22893_ (.A(net5822),
    .B(net6190),
    .Y(_14615_));
 AOI211x1_ASAP7_75t_R _22894_ (.A1(net6190),
    .A2(net5811),
    .B(_14615_),
    .C(net5807),
    .Y(_14616_));
 OAI21x1_ASAP7_75t_R _22895_ (.A1(_14614_),
    .A2(_14616_),
    .B(net5794),
    .Y(_14617_));
 AOI21x1_ASAP7_75t_R _22896_ (.A1(_14375_),
    .A2(_14420_),
    .B(net5783),
    .Y(_14618_));
 OA21x2_ASAP7_75t_R _22897_ (.A1(net4908),
    .A2(net4572),
    .B(net5787),
    .Y(_14619_));
 OAI21x1_ASAP7_75t_R _22898_ (.A1(_14618_),
    .A2(_14619_),
    .B(net5800),
    .Y(_14620_));
 AOI21x1_ASAP7_75t_R _22899_ (.A1(_14617_),
    .A2(_14620_),
    .B(net5792),
    .Y(_14621_));
 NOR2x1_ASAP7_75t_R _22900_ (.A(_14613_),
    .B(_14621_),
    .Y(_14622_));
 AND3x1_ASAP7_75t_R _22901_ (.A(net6182),
    .B(net6183),
    .C(_01181_),
    .Y(_14623_));
 INVx1_ASAP7_75t_R _22902_ (.A(_14444_),
    .Y(_14624_));
 NOR2x1_ASAP7_75t_R _22903_ (.A(_14623_),
    .B(_14624_),
    .Y(_14625_));
 OAI21x1_ASAP7_75t_R _22904_ (.A1(net5786),
    .A2(net5167),
    .B(net5792),
    .Y(_14626_));
 AOI21x1_ASAP7_75t_R _22905_ (.A1(net4906),
    .A2(net5008),
    .B(net5802),
    .Y(_14627_));
 OAI21x1_ASAP7_75t_R _22906_ (.A1(_14626_),
    .A2(_14627_),
    .B(net5793),
    .Y(_14628_));
 AOI21x1_ASAP7_75t_R _22907_ (.A1(net5460),
    .A2(_14625_),
    .B(_14628_),
    .Y(_14629_));
 OAI21x1_ASAP7_75t_R _22908_ (.A1(_01186_),
    .A2(net5785),
    .B(net5460),
    .Y(_14630_));
 OAI21x1_ASAP7_75t_R _22909_ (.A1(_14630_),
    .A2(_14582_),
    .B(net5799),
    .Y(_14631_));
 NAND2x1_ASAP7_75t_R _22910_ (.A(_01170_),
    .B(net5289),
    .Y(_14632_));
 OA21x2_ASAP7_75t_R _22911_ (.A1(net6188),
    .A2(net6189),
    .B(_14632_),
    .Y(_14633_));
 INVx1_ASAP7_75t_R _22912_ (.A(_14633_),
    .Y(_14634_));
 AOI21x1_ASAP7_75t_R _22913_ (.A1(_14450_),
    .A2(_14634_),
    .B(net5807),
    .Y(_14635_));
 OAI21x1_ASAP7_75t_R _22914_ (.A1(_14357_),
    .A2(_14516_),
    .B(net5792),
    .Y(_14636_));
 NOR2x1_ASAP7_75t_R _22915_ (.A(_14635_),
    .B(_14636_),
    .Y(_14637_));
 OAI21x1_ASAP7_75t_R _22916_ (.A1(_14631_),
    .A2(_14637_),
    .B(net6181),
    .Y(_14638_));
 OAI21x1_ASAP7_75t_R _22917_ (.A1(_14629_),
    .A2(_14638_),
    .B(_14416_),
    .Y(_14639_));
 OAI22x1_ASAP7_75t_R _22918_ (.A1(_14588_),
    .A2(_14606_),
    .B1(_14622_),
    .B2(_14639_),
    .Y(_00074_));
 NOR2x1_ASAP7_75t_R _22919_ (.A(net5786),
    .B(_14474_),
    .Y(_14640_));
 INVx1_ASAP7_75t_R _22920_ (.A(_14640_),
    .Y(_14641_));
 OA21x2_ASAP7_75t_R _22921_ (.A1(_14641_),
    .A2(net5461),
    .B(_14360_),
    .Y(_14642_));
 AO21x1_ASAP7_75t_R _22922_ (.A1(net5453),
    .A2(net4913),
    .B(net5789),
    .Y(_14643_));
 AO21x1_ASAP7_75t_R _22923_ (.A1(_14643_),
    .A2(_14478_),
    .B(net5792),
    .Y(_14644_));
 AOI21x1_ASAP7_75t_R _22924_ (.A1(_14642_),
    .A2(_14644_),
    .B(net5796),
    .Y(_14645_));
 AO21x1_ASAP7_75t_R _22925_ (.A1(net5789),
    .A2(net5163),
    .B(net5461),
    .Y(_14646_));
 OAI21x1_ASAP7_75t_R _22926_ (.A1(_14594_),
    .A2(_14646_),
    .B(net5796),
    .Y(_14647_));
 NOR2x1p5_ASAP7_75t_R _22927_ (.A(net4758),
    .B(_14517_),
    .Y(_14648_));
 NOR2x1_ASAP7_75t_R _22928_ (.A(net5286),
    .B(net5813),
    .Y(_14649_));
 OA21x2_ASAP7_75t_R _22929_ (.A1(_14649_),
    .A2(_14633_),
    .B(net5790),
    .Y(_14650_));
 NOR3x1_ASAP7_75t_R _22930_ (.A(net4571),
    .B(_14650_),
    .C(net5792),
    .Y(_14651_));
 OAI21x1_ASAP7_75t_R _22931_ (.A1(_14647_),
    .A2(_14651_),
    .B(net6181),
    .Y(_14652_));
 NOR2x1_ASAP7_75t_R _22932_ (.A(_14645_),
    .B(_14652_),
    .Y(_14653_));
 AO21x1_ASAP7_75t_R _22933_ (.A1(_14559_),
    .A2(net4905),
    .B(net5805),
    .Y(_14654_));
 AO21x1_ASAP7_75t_R _22934_ (.A1(_14580_),
    .A2(net5008),
    .B(net5788),
    .Y(_14655_));
 AO21x1_ASAP7_75t_R _22935_ (.A1(_14654_),
    .A2(_14655_),
    .B(net5796),
    .Y(_14656_));
 AO21x1_ASAP7_75t_R _22936_ (.A1(_14312_),
    .A2(_14565_),
    .B(net5799),
    .Y(_14657_));
 AOI21x1_ASAP7_75t_R _22937_ (.A1(_14656_),
    .A2(_14657_),
    .B(net5461),
    .Y(_14658_));
 OA21x2_ASAP7_75t_R _22938_ (.A1(net6186),
    .A2(net6187),
    .B(_14343_),
    .Y(_14659_));
 OAI21x1_ASAP7_75t_R _22939_ (.A1(_14659_),
    .A2(_14633_),
    .B(net5788),
    .Y(_14660_));
 OAI21x1_ASAP7_75t_R _22940_ (.A1(_14357_),
    .A2(_14516_),
    .B(_14660_),
    .Y(_14661_));
 NOR2x1_ASAP7_75t_R _22941_ (.A(net5790),
    .B(_14649_),
    .Y(_14662_));
 AOI21x1_ASAP7_75t_R _22942_ (.A1(net5458),
    .A2(_14662_),
    .B(net5796),
    .Y(_14663_));
 AOI21x1_ASAP7_75t_R _22943_ (.A1(net5796),
    .A2(_14661_),
    .B(_14663_),
    .Y(_14664_));
 OAI21x1_ASAP7_75t_R _22944_ (.A1(net5792),
    .A2(_14664_),
    .B(_14393_),
    .Y(_14665_));
 OAI21x1_ASAP7_75t_R _22945_ (.A1(_14658_),
    .A2(_14665_),
    .B(net6180),
    .Y(_14666_));
 NAND2x1_ASAP7_75t_R _22946_ (.A(net5811),
    .B(net5784),
    .Y(_14667_));
 OAI21x1_ASAP7_75t_R _22947_ (.A1(net5817),
    .A2(net5811),
    .B(net5797),
    .Y(_14668_));
 NOR2x1_ASAP7_75t_R _22948_ (.A(_14615_),
    .B(_14668_),
    .Y(_14669_));
 AOI21x1_ASAP7_75t_R _22949_ (.A1(_14667_),
    .A2(_14669_),
    .B(net5792),
    .Y(_14670_));
 AO21x1_ASAP7_75t_R _22950_ (.A1(_14593_),
    .A2(net5006),
    .B(net5787),
    .Y(_14671_));
 NAND2x1_ASAP7_75t_R _22951_ (.A(_14671_),
    .B(_14544_),
    .Y(_14672_));
 AOI21x1_ASAP7_75t_R _22952_ (.A1(_14670_),
    .A2(_14672_),
    .B(net6181),
    .Y(_14673_));
 OAI21x1_ASAP7_75t_R _22953_ (.A1(_14273_),
    .A2(_14461_),
    .B(net5783),
    .Y(_14674_));
 AO21x1_ASAP7_75t_R _22954_ (.A1(_14386_),
    .A2(net5006),
    .B(net5783),
    .Y(_14675_));
 AOI21x1_ASAP7_75t_R _22955_ (.A1(_14674_),
    .A2(_14675_),
    .B(net5797),
    .Y(_14676_));
 AND2x2_ASAP7_75t_R _22956_ (.A(_14454_),
    .B(_14421_),
    .Y(_14677_));
 NAND2x1_ASAP7_75t_R _22957_ (.A(net5808),
    .B(_14318_),
    .Y(_14678_));
 OAI21x1_ASAP7_75t_R _22958_ (.A1(_14678_),
    .A2(_14539_),
    .B(net5797),
    .Y(_14679_));
 AOI21x1_ASAP7_75t_R _22959_ (.A1(net5783),
    .A2(_14677_),
    .B(_14679_),
    .Y(_14680_));
 OAI21x1_ASAP7_75t_R _22960_ (.A1(_14676_),
    .A2(_14680_),
    .B(net5792),
    .Y(_14681_));
 NAND2x1_ASAP7_75t_R _22961_ (.A(_14673_),
    .B(_14681_),
    .Y(_14682_));
 AOI21x1_ASAP7_75t_R _22962_ (.A1(net5789),
    .A2(net5005),
    .B(net5795),
    .Y(_14683_));
 OAI21x1_ASAP7_75t_R _22963_ (.A1(_14535_),
    .A2(_14564_),
    .B(net5806),
    .Y(_14684_));
 AOI21x1_ASAP7_75t_R _22964_ (.A1(_14683_),
    .A2(_14684_),
    .B(net5792),
    .Y(_14685_));
 AOI21x1_ASAP7_75t_R _22965_ (.A1(_14426_),
    .A2(_14468_),
    .B(net5800),
    .Y(_14686_));
 AO21x1_ASAP7_75t_R _22966_ (.A1(net5462),
    .A2(_14459_),
    .B(net5787),
    .Y(_14687_));
 NAND2x1_ASAP7_75t_R _22967_ (.A(_14686_),
    .B(_14687_),
    .Y(_14688_));
 AOI21x1_ASAP7_75t_R _22968_ (.A1(_14685_),
    .A2(_14688_),
    .B(net5782),
    .Y(_14689_));
 NOR2x1_ASAP7_75t_R _22969_ (.A(net5286),
    .B(net5820),
    .Y(_14690_));
 OAI21x1_ASAP7_75t_R _22970_ (.A1(net5168),
    .A2(_14690_),
    .B(net5789),
    .Y(_14691_));
 AOI21x1_ASAP7_75t_R _22971_ (.A1(_14572_),
    .A2(_14691_),
    .B(net5800),
    .Y(_14692_));
 AO21x1_ASAP7_75t_R _22972_ (.A1(net5167),
    .A2(net5005),
    .B(net5806),
    .Y(_14693_));
 OAI21x1_ASAP7_75t_R _22973_ (.A1(_14461_),
    .A2(net4908),
    .B(net5806),
    .Y(_14694_));
 AOI21x1_ASAP7_75t_R _22974_ (.A1(_14693_),
    .A2(_14694_),
    .B(net5795),
    .Y(_14695_));
 OAI21x1_ASAP7_75t_R _22975_ (.A1(_14692_),
    .A2(_14695_),
    .B(net5792),
    .Y(_14696_));
 AOI21x1_ASAP7_75t_R _22976_ (.A1(_14689_),
    .A2(_14696_),
    .B(net6180),
    .Y(_14697_));
 NAND2x1_ASAP7_75t_R _22977_ (.A(_14682_),
    .B(_14697_),
    .Y(_14698_));
 OAI21x1_ASAP7_75t_R _22978_ (.A1(_14653_),
    .A2(_14666_),
    .B(_14698_),
    .Y(_00075_));
 NOR2x1_ASAP7_75t_R _22979_ (.A(net5785),
    .B(_14381_),
    .Y(_14699_));
 AOI21x1_ASAP7_75t_R _22980_ (.A1(net4760),
    .A2(_14699_),
    .B(net5799),
    .Y(_14700_));
 OAI21x1_ASAP7_75t_R _22981_ (.A1(net5785),
    .A2(_14500_),
    .B(net5799),
    .Y(_14701_));
 NOR2x1_ASAP7_75t_R _22982_ (.A(net5814),
    .B(_14515_),
    .Y(_14702_));
 NOR2x1_ASAP7_75t_R _22983_ (.A(net5810),
    .B(_14702_),
    .Y(_14703_));
 OAI21x1_ASAP7_75t_R _22984_ (.A1(_14701_),
    .A2(_14703_),
    .B(net5792),
    .Y(_14704_));
 AOI21x1_ASAP7_75t_R _22985_ (.A1(net4912),
    .A2(_14700_),
    .B(_14704_),
    .Y(_14705_));
 AO21x1_ASAP7_75t_R _22986_ (.A1(net5785),
    .A2(net5821),
    .B(net5799),
    .Y(_14706_));
 OA21x2_ASAP7_75t_R _22987_ (.A1(_14443_),
    .A2(_14649_),
    .B(net5805),
    .Y(_14707_));
 OAI21x1_ASAP7_75t_R _22988_ (.A1(_14706_),
    .A2(_14707_),
    .B(net5461),
    .Y(_14708_));
 NOR2x1_ASAP7_75t_R _22989_ (.A(net5804),
    .B(_14381_),
    .Y(_14709_));
 AO21x1_ASAP7_75t_R _22990_ (.A1(_14505_),
    .A2(net5804),
    .B(net5793),
    .Y(_14710_));
 NOR2x1_ASAP7_75t_R _22991_ (.A(net5785),
    .B(_14426_),
    .Y(_14711_));
 AOI211x1_ASAP7_75t_R _22992_ (.A1(_14709_),
    .A2(_14426_),
    .B(_14710_),
    .C(_14711_),
    .Y(_14712_));
 OAI21x1_ASAP7_75t_R _22993_ (.A1(_14708_),
    .A2(_14712_),
    .B(net5781),
    .Y(_14713_));
 NOR2x1_ASAP7_75t_R _22994_ (.A(_14705_),
    .B(_14713_),
    .Y(_14714_));
 OAI21x1_ASAP7_75t_R _22995_ (.A1(_14378_),
    .A2(_14460_),
    .B(net5796),
    .Y(_14715_));
 AOI21x1_ASAP7_75t_R _22996_ (.A1(net5456),
    .A2(net5454),
    .B(net5785),
    .Y(_14716_));
 NOR2x1_ASAP7_75t_R _22997_ (.A(_14535_),
    .B(_14347_),
    .Y(_14717_));
 OAI21x1_ASAP7_75t_R _22998_ (.A1(_14716_),
    .A2(_14717_),
    .B(net5799),
    .Y(_14718_));
 AOI21x1_ASAP7_75t_R _22999_ (.A1(_14715_),
    .A2(_14718_),
    .B(net5792),
    .Y(_14719_));
 NAND2x1_ASAP7_75t_R _23000_ (.A(net5814),
    .B(net5459),
    .Y(_14720_));
 NOR2x1_ASAP7_75t_R _23001_ (.A(net5785),
    .B(_14720_),
    .Y(_14721_));
 INVx1_ASAP7_75t_R _23002_ (.A(_14541_),
    .Y(_14722_));
 OAI21x1_ASAP7_75t_R _23003_ (.A1(_14722_),
    .A2(net4914),
    .B(net5799),
    .Y(_14723_));
 NOR2x1_ASAP7_75t_R _23004_ (.A(_14721_),
    .B(_14723_),
    .Y(_14724_));
 AO21x1_ASAP7_75t_R _23005_ (.A1(net6182),
    .A2(net6183),
    .B(_01176_),
    .Y(_14725_));
 OA21x2_ASAP7_75t_R _23006_ (.A1(net5801),
    .A2(net4759),
    .B(_14725_),
    .Y(_14726_));
 OAI21x1_ASAP7_75t_R _23007_ (.A1(net5798),
    .A2(_14726_),
    .B(net5792),
    .Y(_14727_));
 OAI21x1_ASAP7_75t_R _23008_ (.A1(_14724_),
    .A2(_14727_),
    .B(net6181),
    .Y(_14728_));
 OAI21x1_ASAP7_75t_R _23009_ (.A1(_14719_),
    .A2(_14728_),
    .B(net6180),
    .Y(_14729_));
 AO21x1_ASAP7_75t_R _23010_ (.A1(_14319_),
    .A2(net5790),
    .B(net5163),
    .Y(_14730_));
 OAI21x1_ASAP7_75t_R _23011_ (.A1(net4911),
    .A2(_14730_),
    .B(net5792),
    .Y(_14731_));
 OAI21x1_ASAP7_75t_R _23012_ (.A1(net4757),
    .A2(_14502_),
    .B(net5793),
    .Y(_14732_));
 NOR2x1_ASAP7_75t_R _23013_ (.A(_14350_),
    .B(_14732_),
    .Y(_14733_));
 OAI21x1_ASAP7_75t_R _23014_ (.A1(_14733_),
    .A2(_14731_),
    .B(net6181),
    .Y(_14734_));
 OAI21x1_ASAP7_75t_R _23015_ (.A1(net5818),
    .A2(net5459),
    .B(net5785),
    .Y(_14735_));
 NOR2x1_ASAP7_75t_R _23016_ (.A(_14483_),
    .B(_14735_),
    .Y(_14736_));
 OAI21x1_ASAP7_75t_R _23017_ (.A1(_14581_),
    .A2(_14736_),
    .B(net5799),
    .Y(_14737_));
 OA21x2_ASAP7_75t_R _23018_ (.A1(_14564_),
    .A2(_14505_),
    .B(net5785),
    .Y(_14738_));
 AOI21x1_ASAP7_75t_R _23019_ (.A1(net4906),
    .A2(_14720_),
    .B(net5785),
    .Y(_14739_));
 OAI21x1_ASAP7_75t_R _23020_ (.A1(_14738_),
    .A2(_14739_),
    .B(net5793),
    .Y(_14740_));
 AOI21x1_ASAP7_75t_R _23021_ (.A1(_14737_),
    .A2(_14740_),
    .B(net5792),
    .Y(_14741_));
 NOR2x1_ASAP7_75t_R _23022_ (.A(_14741_),
    .B(_14734_),
    .Y(_14742_));
 NOR2x1_ASAP7_75t_R _23023_ (.A(net5793),
    .B(_14351_),
    .Y(_14743_));
 AO21x1_ASAP7_75t_R _23024_ (.A1(_14743_),
    .A2(net4914),
    .B(net5460),
    .Y(_14744_));
 OAI21x1_ASAP7_75t_R _23025_ (.A1(_14443_),
    .A2(_14491_),
    .B(net5794),
    .Y(_14745_));
 OA21x2_ASAP7_75t_R _23026_ (.A1(_14535_),
    .A2(_14483_),
    .B(net5785),
    .Y(_14746_));
 NOR2x1_ASAP7_75t_R _23027_ (.A(_14745_),
    .B(_14746_),
    .Y(_14747_));
 OAI21x1_ASAP7_75t_R _23028_ (.A1(_14744_),
    .A2(_14747_),
    .B(net5781),
    .Y(_14748_));
 AOI21x1_ASAP7_75t_R _23029_ (.A1(net5459),
    .A2(_14426_),
    .B(net5785),
    .Y(_14749_));
 AOI21x1_ASAP7_75t_R _23030_ (.A1(_14375_),
    .A2(_14420_),
    .B(net5802),
    .Y(_14750_));
 OAI21x1_ASAP7_75t_R _23031_ (.A1(_14749_),
    .A2(_14750_),
    .B(net5799),
    .Y(_14751_));
 OAI21x1_ASAP7_75t_R _23032_ (.A1(_14489_),
    .A2(_14616_),
    .B(net5793),
    .Y(_14752_));
 AOI21x1_ASAP7_75t_R _23033_ (.A1(_14751_),
    .A2(_14752_),
    .B(net5792),
    .Y(_14753_));
 OAI21x1_ASAP7_75t_R _23034_ (.A1(_14748_),
    .A2(_14753_),
    .B(_14416_),
    .Y(_14754_));
 OAI22x1_ASAP7_75t_R _23035_ (.A1(_14714_),
    .A2(_14729_),
    .B1(_14742_),
    .B2(_14754_),
    .Y(_00076_));
 AO21x1_ASAP7_75t_R _23036_ (.A1(_14580_),
    .A2(net5809),
    .B(net5800),
    .Y(_14755_));
 AO21x1_ASAP7_75t_R _23037_ (.A1(_14468_),
    .A2(_14375_),
    .B(_14755_),
    .Y(_14756_));
 AO21x1_ASAP7_75t_R _23038_ (.A1(net5453),
    .A2(_14573_),
    .B(net5787),
    .Y(_14757_));
 AO21x1_ASAP7_75t_R _23039_ (.A1(_14757_),
    .A2(_14508_),
    .B(net5795),
    .Y(_14758_));
 AOI21x1_ASAP7_75t_R _23040_ (.A1(_14756_),
    .A2(_14758_),
    .B(net5792),
    .Y(_14759_));
 AO21x1_ASAP7_75t_R _23041_ (.A1(net5785),
    .A2(net6191),
    .B(net5798),
    .Y(_14760_));
 OAI21x1_ASAP7_75t_R _23042_ (.A1(_14760_),
    .A2(_14749_),
    .B(net5792),
    .Y(_14761_));
 OA21x2_ASAP7_75t_R _23043_ (.A1(_14435_),
    .A2(_14532_),
    .B(net5807),
    .Y(_14762_));
 AOI211x1_ASAP7_75t_R _23044_ (.A1(net5784),
    .A2(_14521_),
    .B(_14762_),
    .C(net5794),
    .Y(_14763_));
 OAI21x1_ASAP7_75t_R _23045_ (.A1(_14761_),
    .A2(_14763_),
    .B(net6181),
    .Y(_14764_));
 NOR2x1_ASAP7_75t_R _23046_ (.A(_14759_),
    .B(_14764_),
    .Y(_14765_));
 AOI211x1_ASAP7_75t_R _23047_ (.A1(net5459),
    .A2(_14566_),
    .B(_14699_),
    .C(net5793),
    .Y(_14766_));
 NAND2x1_ASAP7_75t_R _23048_ (.A(net5788),
    .B(_14589_),
    .Y(_14767_));
 NAND2x1_ASAP7_75t_R _23049_ (.A(_14641_),
    .B(_14767_),
    .Y(_14768_));
 AOI21x1_ASAP7_75t_R _23050_ (.A1(net5817),
    .A2(_14566_),
    .B(net5799),
    .Y(_14769_));
 AO21x1_ASAP7_75t_R _23051_ (.A1(_14768_),
    .A2(_14769_),
    .B(net5792),
    .Y(_14770_));
 OAI21x1_ASAP7_75t_R _23052_ (.A1(_14766_),
    .A2(_14770_),
    .B(net5781),
    .Y(_14771_));
 NOR2x1_ASAP7_75t_R _23053_ (.A(_14381_),
    .B(net4909),
    .Y(_14772_));
 NOR3x1_ASAP7_75t_R _23054_ (.A(_14772_),
    .B(_14428_),
    .C(net5800),
    .Y(_14773_));
 AOI21x1_ASAP7_75t_R _23055_ (.A1(net5287),
    .A2(_14260_),
    .B(net5791),
    .Y(_14774_));
 OA21x2_ASAP7_75t_R _23056_ (.A1(net5821),
    .A2(net5459),
    .B(net5159),
    .Y(_14775_));
 AO21x1_ASAP7_75t_R _23057_ (.A1(net5814),
    .A2(_14499_),
    .B(net5166),
    .Y(_14776_));
 AO21x1_ASAP7_75t_R _23058_ (.A1(_14776_),
    .A2(net5785),
    .B(net5793),
    .Y(_14777_));
 OAI21x1_ASAP7_75t_R _23059_ (.A1(_14775_),
    .A2(_14777_),
    .B(net5792),
    .Y(_14778_));
 NOR2x1_ASAP7_75t_R _23060_ (.A(_14773_),
    .B(_14778_),
    .Y(_14779_));
 OAI21x1_ASAP7_75t_R _23061_ (.A1(_14771_),
    .A2(_14779_),
    .B(_14416_),
    .Y(_14780_));
 NAND2x1_ASAP7_75t_R _23062_ (.A(_14400_),
    .B(_14399_),
    .Y(_14781_));
 NOR2x1_ASAP7_75t_R _23063_ (.A(net5789),
    .B(_14388_),
    .Y(_14782_));
 OAI21x1_ASAP7_75t_R _23064_ (.A1(_14649_),
    .A2(_14539_),
    .B(net5809),
    .Y(_14783_));
 OA21x2_ASAP7_75t_R _23065_ (.A1(_14386_),
    .A2(net5809),
    .B(net5800),
    .Y(_14784_));
 AOI21x1_ASAP7_75t_R _23066_ (.A1(_14783_),
    .A2(_14784_),
    .B(net5792),
    .Y(_14785_));
 OAI21x1_ASAP7_75t_R _23067_ (.A1(_14781_),
    .A2(_14782_),
    .B(_14785_),
    .Y(_14786_));
 OA21x2_ASAP7_75t_R _23068_ (.A1(net5809),
    .A2(net5817),
    .B(net5797),
    .Y(_14787_));
 AOI21x1_ASAP7_75t_R _23069_ (.A1(_14787_),
    .A2(_14462_),
    .B(net5461),
    .Y(_14788_));
 AOI21x1_ASAP7_75t_R _23070_ (.A1(net5453),
    .A2(_14774_),
    .B(net5795),
    .Y(_14789_));
 AO21x1_ASAP7_75t_R _23071_ (.A1(_14421_),
    .A2(net5008),
    .B(net5809),
    .Y(_14790_));
 NAND2x1_ASAP7_75t_R _23072_ (.A(_14789_),
    .B(_14790_),
    .Y(_14791_));
 AOI21x1_ASAP7_75t_R _23073_ (.A1(_14788_),
    .A2(_14791_),
    .B(net6181),
    .Y(_14792_));
 NAND2x1_ASAP7_75t_R _23074_ (.A(_14786_),
    .B(_14792_),
    .Y(_14793_));
 NOR2x1_ASAP7_75t_R _23075_ (.A(_14516_),
    .B(_14444_),
    .Y(_14794_));
 NOR2x1_ASAP7_75t_R _23076_ (.A(_14632_),
    .B(net5819),
    .Y(_14795_));
 OAI21x1_ASAP7_75t_R _23077_ (.A1(net5805),
    .A2(_14795_),
    .B(net5797),
    .Y(_14796_));
 INVx1_ASAP7_75t_R _23078_ (.A(_14401_),
    .Y(_14797_));
 AOI21x1_ASAP7_75t_R _23079_ (.A1(net4909),
    .A2(_14797_),
    .B(net5461),
    .Y(_14798_));
 OAI21x1_ASAP7_75t_R _23080_ (.A1(_14794_),
    .A2(_14796_),
    .B(_14798_),
    .Y(_14799_));
 AO21x1_ASAP7_75t_R _23081_ (.A1(_14580_),
    .A2(net5006),
    .B(net5783),
    .Y(_14800_));
 AO21x1_ASAP7_75t_R _23082_ (.A1(_14269_),
    .A2(_14268_),
    .B(net5288),
    .Y(_14801_));
 AOI21x1_ASAP7_75t_R _23083_ (.A1(_14801_),
    .A2(_14468_),
    .B(net5797),
    .Y(_14802_));
 NAND2x1_ASAP7_75t_R _23084_ (.A(_14800_),
    .B(_14802_),
    .Y(_14803_));
 OA21x2_ASAP7_75t_R _23085_ (.A1(net5808),
    .A2(net5165),
    .B(net5797),
    .Y(_14804_));
 AO21x1_ASAP7_75t_R _23086_ (.A1(_14532_),
    .A2(net5813),
    .B(net5784),
    .Y(_14805_));
 AOI21x1_ASAP7_75t_R _23087_ (.A1(_14804_),
    .A2(_14805_),
    .B(net5792),
    .Y(_14806_));
 AOI21x1_ASAP7_75t_R _23088_ (.A1(_14803_),
    .A2(_14806_),
    .B(net5780),
    .Y(_14807_));
 AOI21x1_ASAP7_75t_R _23089_ (.A1(_14799_),
    .A2(_14807_),
    .B(_14416_),
    .Y(_14808_));
 NAND2x1_ASAP7_75t_R _23090_ (.A(_14793_),
    .B(_14808_),
    .Y(_14809_));
 OAI21x1_ASAP7_75t_R _23091_ (.A1(_14765_),
    .A2(_14780_),
    .B(_14809_),
    .Y(_00077_));
 NAND2x1_ASAP7_75t_R _23092_ (.A(_14374_),
    .B(_14450_),
    .Y(_14810_));
 AND2x2_ASAP7_75t_R _23093_ (.A(_14774_),
    .B(_14501_),
    .Y(_14811_));
 AOI21x1_ASAP7_75t_R _23094_ (.A1(net5785),
    .A2(_14810_),
    .B(_14811_),
    .Y(_14812_));
 AO21x1_ASAP7_75t_R _23095_ (.A1(net5821),
    .A2(net5160),
    .B(_14767_),
    .Y(_14813_));
 NOR2x1_ASAP7_75t_R _23096_ (.A(_14782_),
    .B(_14325_),
    .Y(_14814_));
 NAND2x1_ASAP7_75t_R _23097_ (.A(_14813_),
    .B(_14814_),
    .Y(_14815_));
 OAI21x1_ASAP7_75t_R _23098_ (.A1(net5799),
    .A2(_14812_),
    .B(_14815_),
    .Y(_14816_));
 OA21x2_ASAP7_75t_R _23099_ (.A1(_14292_),
    .A2(net5163),
    .B(net5785),
    .Y(_14817_));
 OAI21x1_ASAP7_75t_R _23100_ (.A1(_14710_),
    .A2(_14817_),
    .B(net5792),
    .Y(_14818_));
 NAND2x1_ASAP7_75t_R _23101_ (.A(_01179_),
    .B(_01185_),
    .Y(_14819_));
 AOI21x1_ASAP7_75t_R _23102_ (.A1(net5456),
    .A2(net5454),
    .B(net5810),
    .Y(_14820_));
 AOI211x1_ASAP7_75t_R _23103_ (.A1(net5804),
    .A2(_14819_),
    .B(_14820_),
    .C(net5799),
    .Y(_14821_));
 OAI21x1_ASAP7_75t_R _23104_ (.A1(_14818_),
    .A2(_14821_),
    .B(net5781),
    .Y(_14822_));
 AOI21x1_ASAP7_75t_R _23105_ (.A1(net5461),
    .A2(_14816_),
    .B(_14822_),
    .Y(_14823_));
 NOR2x1_ASAP7_75t_R _23106_ (.A(net5797),
    .B(_14640_),
    .Y(_14824_));
 OAI21x1_ASAP7_75t_R _23107_ (.A1(_14623_),
    .A2(_14624_),
    .B(_14824_),
    .Y(_14825_));
 AOI21x1_ASAP7_75t_R _23108_ (.A1(_14420_),
    .A2(_14421_),
    .B(net5802),
    .Y(_14826_));
 NAND2x1_ASAP7_75t_R _23109_ (.A(net5810),
    .B(_14449_),
    .Y(_14827_));
 NOR2x1_ASAP7_75t_R _23110_ (.A(_14500_),
    .B(_14827_),
    .Y(_14828_));
 OAI21x1_ASAP7_75t_R _23111_ (.A1(_14826_),
    .A2(_14828_),
    .B(net5793),
    .Y(_14829_));
 AOI21x1_ASAP7_75t_R _23112_ (.A1(_14825_),
    .A2(_14829_),
    .B(net5460),
    .Y(_14830_));
 AO21x1_ASAP7_75t_R _23113_ (.A1(_14388_),
    .A2(net6190),
    .B(net5807),
    .Y(_14831_));
 OA21x2_ASAP7_75t_R _23114_ (.A1(_14386_),
    .A2(net5783),
    .B(net5800),
    .Y(_14832_));
 AO21x1_ASAP7_75t_R _23115_ (.A1(_14831_),
    .A2(_14832_),
    .B(net5792),
    .Y(_14833_));
 AOI21x1_ASAP7_75t_R _23116_ (.A1(_14559_),
    .A2(_14720_),
    .B(net5805),
    .Y(_14834_));
 NOR2x1_ASAP7_75t_R _23117_ (.A(_14795_),
    .B(_14678_),
    .Y(_14835_));
 NOR3x1_ASAP7_75t_R _23118_ (.A(_14834_),
    .B(net5800),
    .C(_14835_),
    .Y(_14836_));
 OAI21x1_ASAP7_75t_R _23119_ (.A1(_14833_),
    .A2(_14836_),
    .B(net6181),
    .Y(_14837_));
 OAI21x1_ASAP7_75t_R _23120_ (.A1(_14830_),
    .A2(_14837_),
    .B(_14416_),
    .Y(_14838_));
 OAI21x1_ASAP7_75t_R _23121_ (.A1(_14443_),
    .A2(_14444_),
    .B(_14551_),
    .Y(_14839_));
 NAND2x1_ASAP7_75t_R _23122_ (.A(_14767_),
    .B(_14827_),
    .Y(_14840_));
 AOI21x1_ASAP7_75t_R _23123_ (.A1(_14769_),
    .A2(_14840_),
    .B(net6181),
    .Y(_14841_));
 NAND2x1_ASAP7_75t_R _23124_ (.A(_14839_),
    .B(_14841_),
    .Y(_14842_));
 AOI21x1_ASAP7_75t_R _23125_ (.A1(net5796),
    .A2(_14585_),
    .B(_14393_),
    .Y(_14843_));
 INVx1_ASAP7_75t_R _23126_ (.A(_14347_),
    .Y(_14844_));
 AOI21x1_ASAP7_75t_R _23127_ (.A1(net5454),
    .A2(_14844_),
    .B(net5793),
    .Y(_14845_));
 NAND2x1_ASAP7_75t_R _23128_ (.A(_14357_),
    .B(_14845_),
    .Y(_14846_));
 AOI21x1_ASAP7_75t_R _23129_ (.A1(_14843_),
    .A2(_14846_),
    .B(net5792),
    .Y(_14847_));
 NAND2x1_ASAP7_75t_R _23130_ (.A(_14842_),
    .B(_14847_),
    .Y(_14848_));
 NAND2x1_ASAP7_75t_R _23131_ (.A(net5787),
    .B(_14459_),
    .Y(_14849_));
 AOI21x1_ASAP7_75t_R _23132_ (.A1(_14849_),
    .A2(_14502_),
    .B(_14461_),
    .Y(_14850_));
 NAND2x1_ASAP7_75t_R _23133_ (.A(net6185),
    .B(net5807),
    .Y(_14851_));
 AOI21x1_ASAP7_75t_R _23134_ (.A1(_14851_),
    .A2(_14669_),
    .B(net6181),
    .Y(_14852_));
 OAI21x1_ASAP7_75t_R _23135_ (.A1(net5796),
    .A2(_14850_),
    .B(_14852_),
    .Y(_14853_));
 AOI21x1_ASAP7_75t_R _23136_ (.A1(net5806),
    .A2(_14461_),
    .B(net5795),
    .Y(_14854_));
 OAI21x1_ASAP7_75t_R _23137_ (.A1(net4758),
    .A2(_14649_),
    .B(net5789),
    .Y(_14855_));
 AOI21x1_ASAP7_75t_R _23138_ (.A1(_14854_),
    .A2(_14855_),
    .B(net5782),
    .Y(_14856_));
 AO21x1_ASAP7_75t_R _23139_ (.A1(net5790),
    .A2(_01180_),
    .B(net5799),
    .Y(_14857_));
 AO21x1_ASAP7_75t_R _23140_ (.A1(net5453),
    .A2(_14774_),
    .B(_14857_),
    .Y(_14858_));
 AOI21x1_ASAP7_75t_R _23141_ (.A1(_14856_),
    .A2(_14858_),
    .B(net5461),
    .Y(_14859_));
 AOI21x1_ASAP7_75t_R _23142_ (.A1(_14853_),
    .A2(_14859_),
    .B(_14416_),
    .Y(_14860_));
 NAND2x1_ASAP7_75t_R _23143_ (.A(_14848_),
    .B(_14860_),
    .Y(_14861_));
 OAI21x1_ASAP7_75t_R _23144_ (.A1(_14823_),
    .A2(_14838_),
    .B(_14861_),
    .Y(_00078_));
 NOR2x1_ASAP7_75t_R _23145_ (.A(_14722_),
    .B(_14347_),
    .Y(_14862_));
 AO21x1_ASAP7_75t_R _23146_ (.A1(net4907),
    .A2(net5804),
    .B(net5799),
    .Y(_14863_));
 OAI21x1_ASAP7_75t_R _23147_ (.A1(_14862_),
    .A2(_14863_),
    .B(net5792),
    .Y(_14864_));
 OAI21x1_ASAP7_75t_R _23148_ (.A1(_14349_),
    .A2(_14517_),
    .B(net5799),
    .Y(_14865_));
 OA21x2_ASAP7_75t_R _23149_ (.A1(_14496_),
    .A2(_14505_),
    .B(net5785),
    .Y(_14866_));
 NOR2x1_ASAP7_75t_R _23150_ (.A(_14865_),
    .B(_14866_),
    .Y(_14867_));
 OAI21x1_ASAP7_75t_R _23151_ (.A1(_14864_),
    .A2(_14867_),
    .B(net5781),
    .Y(_14868_));
 OA21x2_ASAP7_75t_R _23152_ (.A1(_14690_),
    .A2(_14319_),
    .B(net5789),
    .Y(_14869_));
 OAI21x1_ASAP7_75t_R _23153_ (.A1(_14869_),
    .A2(_14648_),
    .B(net5799),
    .Y(_14870_));
 OAI21x1_ASAP7_75t_R _23154_ (.A1(_14608_),
    .A2(_14811_),
    .B(net5793),
    .Y(_14871_));
 AOI21x1_ASAP7_75t_R _23155_ (.A1(_14870_),
    .A2(_14871_),
    .B(net5792),
    .Y(_14872_));
 NOR2x1_ASAP7_75t_R _23156_ (.A(_14868_),
    .B(_14872_),
    .Y(_14873_));
 AO21x1_ASAP7_75t_R _23157_ (.A1(net4758),
    .A2(net5807),
    .B(net5800),
    .Y(_14874_));
 NOR2x1_ASAP7_75t_R _23158_ (.A(_14532_),
    .B(_14667_),
    .Y(_14875_));
 OAI21x1_ASAP7_75t_R _23159_ (.A1(_14874_),
    .A2(_14875_),
    .B(net5460),
    .Y(_14876_));
 NOR2x1_ASAP7_75t_R _23160_ (.A(_14702_),
    .B(_14827_),
    .Y(_14877_));
 NAND2x1_ASAP7_75t_R _23161_ (.A(net5799),
    .B(_14735_),
    .Y(_14878_));
 NOR2x1_ASAP7_75t_R _23162_ (.A(_14877_),
    .B(_14878_),
    .Y(_14879_));
 OAI21x1_ASAP7_75t_R _23163_ (.A1(_14876_),
    .A2(_14879_),
    .B(net6181),
    .Y(_14880_));
 NOR2x1_ASAP7_75t_R _23164_ (.A(net5817),
    .B(net5785),
    .Y(_14881_));
 AOI21x1_ASAP7_75t_R _23165_ (.A1(_14487_),
    .A2(_14550_),
    .B(net5801),
    .Y(_14882_));
 OAI21x1_ASAP7_75t_R _23166_ (.A1(_14881_),
    .A2(_14882_),
    .B(net5798),
    .Y(_14883_));
 AOI21x1_ASAP7_75t_R _23167_ (.A1(_14420_),
    .A2(_14450_),
    .B(net5786),
    .Y(_14884_));
 OAI21x1_ASAP7_75t_R _23168_ (.A1(_14884_),
    .A2(_14616_),
    .B(net5797),
    .Y(_14885_));
 AOI21x1_ASAP7_75t_R _23169_ (.A1(_14883_),
    .A2(_14885_),
    .B(net5460),
    .Y(_14886_));
 OAI21x1_ASAP7_75t_R _23170_ (.A1(_14880_),
    .A2(_14886_),
    .B(net6180),
    .Y(_14887_));
 INVx1_ASAP7_75t_R _23171_ (.A(_14485_),
    .Y(_14888_));
 OA211x2_ASAP7_75t_R _23172_ (.A1(net5786),
    .A2(_14388_),
    .B(_14851_),
    .C(net5800),
    .Y(_14889_));
 AND3x1_ASAP7_75t_R _23173_ (.A(net6182),
    .B(net6183),
    .C(_01176_),
    .Y(_14890_));
 OAI21x1_ASAP7_75t_R _23174_ (.A1(_14890_),
    .A2(_14309_),
    .B(net5792),
    .Y(_14891_));
 AOI21x1_ASAP7_75t_R _23175_ (.A1(_14888_),
    .A2(_14889_),
    .B(_14891_),
    .Y(_14892_));
 OA21x2_ASAP7_75t_R _23176_ (.A1(net5804),
    .A2(_01185_),
    .B(net5793),
    .Y(_14893_));
 NAND2x1_ASAP7_75t_R _23177_ (.A(net5804),
    .B(_14477_),
    .Y(_14894_));
 AND3x1_ASAP7_75t_R _23178_ (.A(_14893_),
    .B(_14405_),
    .C(_14894_),
    .Y(_14895_));
 NOR2x1_ASAP7_75t_R _23179_ (.A(net5256),
    .B(net5820),
    .Y(_14896_));
 OAI21x1_ASAP7_75t_R _23180_ (.A1(_14896_),
    .A2(net4756),
    .B(net5799),
    .Y(_14897_));
 NOR2x1_ASAP7_75t_R _23181_ (.A(_14722_),
    .B(_14517_),
    .Y(_14898_));
 OAI21x1_ASAP7_75t_R _23182_ (.A1(_14897_),
    .A2(_14898_),
    .B(net5461),
    .Y(_14899_));
 OAI21x1_ASAP7_75t_R _23183_ (.A1(_14895_),
    .A2(_14899_),
    .B(net6181),
    .Y(_14900_));
 NOR2x1_ASAP7_75t_R _23184_ (.A(_14892_),
    .B(_14900_),
    .Y(_14901_));
 NOR2x1_ASAP7_75t_R _23185_ (.A(_14795_),
    .B(_14347_),
    .Y(_14902_));
 AOI21x1_ASAP7_75t_R _23186_ (.A1(net5454),
    .A2(_14450_),
    .B(net5788),
    .Y(_14903_));
 OAI21x1_ASAP7_75t_R _23187_ (.A1(_14902_),
    .A2(_14903_),
    .B(net5800),
    .Y(_14904_));
 AOI21x1_ASAP7_75t_R _23188_ (.A1(net5006),
    .A2(_14386_),
    .B(net5808),
    .Y(_14905_));
 AOI21x1_ASAP7_75t_R _23189_ (.A1(net5167),
    .A2(_14450_),
    .B(net5784),
    .Y(_14906_));
 OAI21x1_ASAP7_75t_R _23190_ (.A1(_14905_),
    .A2(_14906_),
    .B(net5794),
    .Y(_14907_));
 AOI21x1_ASAP7_75t_R _23191_ (.A1(_14904_),
    .A2(_14907_),
    .B(net5460),
    .Y(_14908_));
 AO21x1_ASAP7_75t_R _23192_ (.A1(net5802),
    .A2(net5166),
    .B(net5793),
    .Y(_14909_));
 OAI21x1_ASAP7_75t_R _23193_ (.A1(_14909_),
    .A2(_14820_),
    .B(net5460),
    .Y(_14910_));
 AO21x1_ASAP7_75t_R _23194_ (.A1(_14483_),
    .A2(net5785),
    .B(_14505_),
    .Y(_14911_));
 NOR2x1_ASAP7_75t_R _23195_ (.A(_14309_),
    .B(_14911_),
    .Y(_14912_));
 OAI21x1_ASAP7_75t_R _23196_ (.A1(_14910_),
    .A2(_14912_),
    .B(net5781),
    .Y(_14913_));
 OAI21x1_ASAP7_75t_R _23197_ (.A1(_14908_),
    .A2(_14913_),
    .B(_14416_),
    .Y(_14914_));
 OAI22x1_ASAP7_75t_R _23198_ (.A1(_14873_),
    .A2(_14887_),
    .B1(_14901_),
    .B2(_14914_),
    .Y(_00079_));
 INVx1_ASAP7_75t_R _23199_ (.A(_00592_),
    .Y(_14915_));
 XOR2x2_ASAP7_75t_R _23200_ (.A(_12121_),
    .B(_14915_),
    .Y(_14916_));
 XNOR2x2_ASAP7_75t_R _23201_ (.A(_00655_),
    .B(_00662_),
    .Y(_14917_));
 XOR2x2_ASAP7_75t_R _23202_ (.A(_00688_),
    .B(_00656_),
    .Y(_14918_));
 XOR2x2_ASAP7_75t_R _23203_ (.A(_14918_),
    .B(_14917_),
    .Y(_14919_));
 NOR2x1_ASAP7_75t_R _23204_ (.A(_14916_),
    .B(_14919_),
    .Y(_14920_));
 XOR2x2_ASAP7_75t_R _23205_ (.A(_12121_),
    .B(net6636),
    .Y(_14921_));
 XOR2x2_ASAP7_75t_R _23206_ (.A(_00655_),
    .B(_00662_),
    .Y(_14922_));
 XOR2x2_ASAP7_75t_R _23207_ (.A(_14918_),
    .B(_14922_),
    .Y(_14923_));
 OAI21x1_ASAP7_75t_R _23208_ (.A1(_14921_),
    .A2(_14923_),
    .B(net6664),
    .Y(_14924_));
 NAND2x1_ASAP7_75t_R _23209_ (.A(_00462_),
    .B(net6455),
    .Y(_14925_));
 OAI21x1_ASAP7_75t_R _23210_ (.A1(_14924_),
    .A2(_14920_),
    .B(_14925_),
    .Y(_14926_));
 XOR2x2_ASAP7_75t_R _23211_ (.A(net6356),
    .B(net6488),
    .Y(_14927_));
 NOR2x1_ASAP7_75t_R _23213_ (.A(net6673),
    .B(_00463_),
    .Y(_14928_));
 XOR2x2_ASAP7_75t_R _23214_ (.A(net6606),
    .B(net6639),
    .Y(_14929_));
 NAND2x1_ASAP7_75t_R _23215_ (.A(_12140_),
    .B(_14929_),
    .Y(_14930_));
 XNOR2x2_ASAP7_75t_R _23216_ (.A(net6639),
    .B(net6606),
    .Y(_14931_));
 NAND2x1_ASAP7_75t_R _23217_ (.A(net6553),
    .B(_14931_),
    .Y(_14932_));
 AOI21x1_ASAP7_75t_R _23218_ (.A1(_14930_),
    .A2(_14932_),
    .B(net6412),
    .Y(_14933_));
 XOR2x2_ASAP7_75t_R _23219_ (.A(net6606),
    .B(_00687_),
    .Y(_14934_));
 NAND2x1_ASAP7_75t_R _23220_ (.A(net6638),
    .B(_14934_),
    .Y(_14935_));
 INVx1_ASAP7_75t_R _23221_ (.A(net6638),
    .Y(_14936_));
 XNOR2x2_ASAP7_75t_R _23222_ (.A(net6606),
    .B(_00687_),
    .Y(_14937_));
 NAND2x1_ASAP7_75t_R _23223_ (.A(_14936_),
    .B(_14937_),
    .Y(_14938_));
 AOI21x1_ASAP7_75t_R _23224_ (.A1(_14935_),
    .A2(_14938_),
    .B(net6410),
    .Y(_14939_));
 OAI21x1_ASAP7_75t_R _23225_ (.A1(_14939_),
    .A2(_14933_),
    .B(net6664),
    .Y(_14940_));
 INVx1_ASAP7_75t_R _23226_ (.A(net6355),
    .Y(_14941_));
 OAI21x1_ASAP7_75t_R _23227_ (.A1(net6409),
    .A2(_14941_),
    .B(net6489),
    .Y(_14942_));
 INVx1_ASAP7_75t_R _23228_ (.A(net6489),
    .Y(_14943_));
 INVx1_ASAP7_75t_R _23229_ (.A(_14928_),
    .Y(_14944_));
 NAND3x1_ASAP7_75t_R _23230_ (.A(net6355),
    .B(_14943_),
    .C(_14944_),
    .Y(_14945_));
 NAND2x1_ASAP7_75t_R _23231_ (.A(_14942_),
    .B(_14945_),
    .Y(_01194_));
 NOR2x1_ASAP7_75t_R _23232_ (.A(net6661),
    .B(_00464_),
    .Y(_14946_));
 INVx1_ASAP7_75t_R _23233_ (.A(_14946_),
    .Y(_14947_));
 INVx1_ASAP7_75t_R _23234_ (.A(net6634),
    .Y(_14948_));
 NOR2x1_ASAP7_75t_R _23235_ (.A(_14948_),
    .B(_12168_),
    .Y(_14949_));
 NOR2x1_ASAP7_75t_R _23236_ (.A(net6634),
    .B(_12164_),
    .Y(_14950_));
 OAI21x1_ASAP7_75t_R _23237_ (.A1(_14949_),
    .A2(_14950_),
    .B(net6437),
    .Y(_14951_));
 INVx1_ASAP7_75t_R _23238_ (.A(_14951_),
    .Y(_14952_));
 NOR3x1_ASAP7_75t_R _23239_ (.A(_14950_),
    .B(_14949_),
    .C(net6437),
    .Y(_14953_));
 OAI21x1_ASAP7_75t_R _23240_ (.A1(_14952_),
    .A2(_14953_),
    .B(net6656),
    .Y(_14954_));
 INVx1_ASAP7_75t_R _23241_ (.A(_00911_),
    .Y(_14955_));
 AOI21x1_ASAP7_75t_R _23242_ (.A1(_14947_),
    .A2(_14954_),
    .B(_14955_),
    .Y(_14956_));
 AND2x2_ASAP7_75t_R _23243_ (.A(net6456),
    .B(_00464_),
    .Y(_14957_));
 INVx1_ASAP7_75t_R _23244_ (.A(_14957_),
    .Y(_14958_));
 NAND2x1_ASAP7_75t_R _23245_ (.A(_14948_),
    .B(_12168_),
    .Y(_14959_));
 INVx1_ASAP7_75t_R _23246_ (.A(net6437),
    .Y(_14960_));
 NOR2x1_ASAP7_75t_R _23247_ (.A(_00657_),
    .B(net6551),
    .Y(_14961_));
 AND2x2_ASAP7_75t_R _23248_ (.A(_00657_),
    .B(net6551),
    .Y(_14962_));
 OAI21x1_ASAP7_75t_R _23249_ (.A1(_14961_),
    .A2(_14962_),
    .B(net6634),
    .Y(_14963_));
 NAND3x1_ASAP7_75t_R _23250_ (.A(_14959_),
    .B(_14960_),
    .C(_14963_),
    .Y(_14964_));
 NAND3x1_ASAP7_75t_R _23251_ (.A(_14964_),
    .B(net6656),
    .C(_14951_),
    .Y(_14965_));
 AOI21x1_ASAP7_75t_R _23252_ (.A1(_14958_),
    .A2(_14965_),
    .B(_00911_),
    .Y(_14966_));
 NOR2x2_ASAP7_75t_R _23253_ (.A(_14956_),
    .B(_14966_),
    .Y(_14967_));
 NAND3x1_ASAP7_75t_R _23256_ (.A(_14944_),
    .B(net6489),
    .C(_14940_),
    .Y(_14969_));
 AO21x1_ASAP7_75t_R _23257_ (.A1(_14944_),
    .A2(_14940_),
    .B(net6489),
    .Y(_14970_));
 NAND2x1p5_ASAP7_75t_R _23258_ (.A(_14970_),
    .B(_14969_),
    .Y(_14971_));
 AOI21x1_ASAP7_75t_R _23260_ (.A1(_14947_),
    .A2(_14954_),
    .B(_00911_),
    .Y(_14972_));
 AOI21x1_ASAP7_75t_R _23261_ (.A1(_14958_),
    .A2(_14965_),
    .B(_14955_),
    .Y(_14973_));
 NOR2x2_ASAP7_75t_R _23262_ (.A(_14972_),
    .B(_14973_),
    .Y(_14974_));
 NOR2x1_ASAP7_75t_R _23264_ (.A(_01193_),
    .B(_14974_),
    .Y(_14975_));
 AOI21x1_ASAP7_75t_R _23265_ (.A1(net6178),
    .A2(net5778),
    .B(net5448),
    .Y(_14976_));
 XOR2x2_ASAP7_75t_R _23266_ (.A(_12192_),
    .B(net6633),
    .Y(_14977_));
 XOR2x2_ASAP7_75t_R _23267_ (.A(_00657_),
    .B(net6579),
    .Y(_14978_));
 XOR2x2_ASAP7_75t_R _23268_ (.A(_12196_),
    .B(_14978_),
    .Y(_14979_));
 NOR2x1_ASAP7_75t_R _23269_ (.A(_14977_),
    .B(_14979_),
    .Y(_14980_));
 XNOR2x2_ASAP7_75t_R _23270_ (.A(net6633),
    .B(_12192_),
    .Y(_14981_));
 XOR2x2_ASAP7_75t_R _23271_ (.A(_12191_),
    .B(_14978_),
    .Y(_14982_));
 NOR2x1_ASAP7_75t_R _23272_ (.A(_14981_),
    .B(_14982_),
    .Y(_14983_));
 OAI21x1_ASAP7_75t_R _23273_ (.A1(_14980_),
    .A2(_14983_),
    .B(net6657),
    .Y(_14984_));
 NOR2x1_ASAP7_75t_R _23274_ (.A(net6669),
    .B(_00522_),
    .Y(_14985_));
 INVx1_ASAP7_75t_R _23275_ (.A(_14985_),
    .Y(_14986_));
 NAND3x1_ASAP7_75t_R _23276_ (.A(_14984_),
    .B(_00912_),
    .C(_14986_),
    .Y(_14987_));
 AO21x1_ASAP7_75t_R _23277_ (.A1(_14984_),
    .A2(_14986_),
    .B(_00912_),
    .Y(_14988_));
 NAND2x1_ASAP7_75t_R _23278_ (.A(_14987_),
    .B(_14988_),
    .Y(_14989_));
 OAI21x1_ASAP7_75t_R _23280_ (.A1(net5158),
    .A2(_14976_),
    .B(net5776),
    .Y(_14991_));
 OAI21x1_ASAP7_75t_R _23281_ (.A1(net5779),
    .A2(net6177),
    .B(_01189_),
    .Y(_14992_));
 INVx1_ASAP7_75t_R _23282_ (.A(_14992_),
    .Y(_14993_));
 NOR2x2_ASAP7_75t_R _23284_ (.A(net5778),
    .B(net5446),
    .Y(_14995_));
 INVx1_ASAP7_75t_R _23285_ (.A(_00912_),
    .Y(_14996_));
 NAND3x1_ASAP7_75t_R _23286_ (.A(_14984_),
    .B(_14996_),
    .C(_14986_),
    .Y(_14997_));
 AO21x1_ASAP7_75t_R _23287_ (.A1(_14984_),
    .A2(_14986_),
    .B(_14996_),
    .Y(_14998_));
 NAND2x1_ASAP7_75t_R _23288_ (.A(_14997_),
    .B(_14998_),
    .Y(_14999_));
 OAI21x1_ASAP7_75t_R _23291_ (.A1(net4904),
    .A2(_14995_),
    .B(net5760),
    .Y(_15002_));
 INVx1_ASAP7_75t_R _23292_ (.A(net5285),
    .Y(_15003_));
 OAI21x1_ASAP7_75t_R _23293_ (.A1(net5777),
    .A2(net6176),
    .B(_15003_),
    .Y(_15004_));
 INVx1_ASAP7_75t_R _23294_ (.A(_15004_),
    .Y(_15005_));
 NAND2x1_ASAP7_75t_R _23295_ (.A(net5776),
    .B(_15005_),
    .Y(_15006_));
 AND2x2_ASAP7_75t_R _23296_ (.A(net6455),
    .B(_00521_),
    .Y(_15007_));
 XOR2x2_ASAP7_75t_R _23297_ (.A(net6581),
    .B(net6579),
    .Y(_15008_));
 INVx1_ASAP7_75t_R _23298_ (.A(_00691_),
    .Y(_15009_));
 XOR2x2_ASAP7_75t_R _23299_ (.A(_15008_),
    .B(_15009_),
    .Y(_15010_));
 XOR2x2_ASAP7_75t_R _23300_ (.A(net6609),
    .B(net6604),
    .Y(_15011_));
 XOR2x2_ASAP7_75t_R _23301_ (.A(_00595_),
    .B(_00659_),
    .Y(_15012_));
 XOR2x2_ASAP7_75t_R _23302_ (.A(_15011_),
    .B(_15012_),
    .Y(_15013_));
 NAND2x1_ASAP7_75t_R _23303_ (.A(_15010_),
    .B(_15013_),
    .Y(_15014_));
 INVx1_ASAP7_75t_R _23304_ (.A(_15010_),
    .Y(_15015_));
 INVx1_ASAP7_75t_R _23305_ (.A(_15013_),
    .Y(_15016_));
 NAND2x1_ASAP7_75t_R _23306_ (.A(_15015_),
    .B(_15016_),
    .Y(_15017_));
 AOI21x1_ASAP7_75t_R _23307_ (.A1(_15014_),
    .A2(_15017_),
    .B(net6455),
    .Y(_15018_));
 OAI21x1_ASAP7_75t_R _23308_ (.A1(_15007_),
    .A2(_15018_),
    .B(net6486),
    .Y(_15019_));
 NOR2x1_ASAP7_75t_R _23309_ (.A(net6664),
    .B(_00521_),
    .Y(_15020_));
 XOR2x2_ASAP7_75t_R _23310_ (.A(_15011_),
    .B(_00595_),
    .Y(_15021_));
 XOR2x2_ASAP7_75t_R _23311_ (.A(_12213_),
    .B(_15008_),
    .Y(_15022_));
 NAND2x1_ASAP7_75t_R _23312_ (.A(_15021_),
    .B(_15022_),
    .Y(_15023_));
 INVx1_ASAP7_75t_R _23313_ (.A(_15021_),
    .Y(_15024_));
 INVx1_ASAP7_75t_R _23314_ (.A(_15022_),
    .Y(_15025_));
 NAND2x1_ASAP7_75t_R _23315_ (.A(_15024_),
    .B(_15025_),
    .Y(_15026_));
 AOI21x1_ASAP7_75t_R _23316_ (.A1(_15023_),
    .A2(_15026_),
    .B(net6455),
    .Y(_15027_));
 INVx1_ASAP7_75t_R _23317_ (.A(net6486),
    .Y(_15028_));
 OAI21x1_ASAP7_75t_R _23318_ (.A1(_15020_),
    .A2(_15027_),
    .B(_15028_),
    .Y(_15029_));
 NAND2x1_ASAP7_75t_R _23319_ (.A(_15019_),
    .B(_15029_),
    .Y(_15030_));
 AND3x1_ASAP7_75t_R _23321_ (.A(_15002_),
    .B(_15006_),
    .C(net5443),
    .Y(_15032_));
 INVx1_ASAP7_75t_R _23323_ (.A(_01190_),
    .Y(_15034_));
 OAI21x1_ASAP7_75t_R _23324_ (.A1(net5777),
    .A2(net6176),
    .B(_15034_),
    .Y(_15035_));
 INVx2_ASAP7_75t_R _23326_ (.A(_15030_),
    .Y(_15037_));
 OA21x2_ASAP7_75t_R _23328_ (.A1(net5760),
    .A2(net4755),
    .B(net5151),
    .Y(_15039_));
 AO21x1_ASAP7_75t_R _23329_ (.A1(_14998_),
    .A2(net6175),
    .B(_01203_),
    .Y(_15040_));
 NOR2x1_ASAP7_75t_R _23330_ (.A(net6668),
    .B(_00520_),
    .Y(_15041_));
 XNOR2x2_ASAP7_75t_R _23331_ (.A(net6632),
    .B(net6608),
    .Y(_15042_));
 INVx1_ASAP7_75t_R _23332_ (.A(_15042_),
    .Y(_15043_));
 XOR2x2_ASAP7_75t_R _23333_ (.A(_00659_),
    .B(_00660_),
    .Y(_15044_));
 XOR2x2_ASAP7_75t_R _23334_ (.A(_15044_),
    .B(_00692_),
    .Y(_15045_));
 NOR2x1_ASAP7_75t_R _23335_ (.A(_15043_),
    .B(_15045_),
    .Y(_15046_));
 XOR2x2_ASAP7_75t_R _23336_ (.A(_15044_),
    .B(_12236_),
    .Y(_15047_));
 NOR2x1_ASAP7_75t_R _23337_ (.A(_15042_),
    .B(_15047_),
    .Y(_15048_));
 OA21x2_ASAP7_75t_R _23338_ (.A1(_15046_),
    .A2(_15048_),
    .B(net6653),
    .Y(_15049_));
 NOR2x1_ASAP7_75t_R _23339_ (.A(_15041_),
    .B(_15049_),
    .Y(_15050_));
 XOR2x2_ASAP7_75t_R _23340_ (.A(_15050_),
    .B(_00915_),
    .Y(_15051_));
 AO21x1_ASAP7_75t_R _23342_ (.A1(_15040_),
    .A2(_15039_),
    .B(net5751),
    .Y(_15053_));
 AOI21x1_ASAP7_75t_R _23343_ (.A1(_14991_),
    .A2(_15032_),
    .B(_15053_),
    .Y(_15054_));
 NOR2x1_ASAP7_75t_R _23344_ (.A(_01191_),
    .B(net5449),
    .Y(_15055_));
 AO21x1_ASAP7_75t_R _23348_ (.A1(_15055_),
    .A2(net5769),
    .B(net5154),
    .Y(_15059_));
 NAND2x1_ASAP7_75t_R _23349_ (.A(net5778),
    .B(net6179),
    .Y(_15060_));
 NOR2x1_ASAP7_75t_R _23350_ (.A(net5450),
    .B(_15060_),
    .Y(_15061_));
 AO21x1_ASAP7_75t_R _23352_ (.A1(net5062),
    .A2(net5451),
    .B(net5776),
    .Y(_15063_));
 NOR2x1_ASAP7_75t_R _23353_ (.A(net5147),
    .B(_15063_),
    .Y(_15064_));
 OAI21x1_ASAP7_75t_R _23355_ (.A1(_15059_),
    .A2(_15064_),
    .B(net5751),
    .Y(_15066_));
 INVx1_ASAP7_75t_R _23356_ (.A(net5147),
    .Y(_15067_));
 INVx1_ASAP7_75t_R _23357_ (.A(_01195_),
    .Y(_15068_));
 AOI21x1_ASAP7_75t_R _23358_ (.A1(_15068_),
    .A2(net5451),
    .B(net5763),
    .Y(_15069_));
 INVx1_ASAP7_75t_R _23359_ (.A(_15055_),
    .Y(_15070_));
 NOR2x1_ASAP7_75t_R _23360_ (.A(net5776),
    .B(_15070_),
    .Y(_15071_));
 AOI211x1_ASAP7_75t_R _23362_ (.A1(_15067_),
    .A2(net4676),
    .B(net4675),
    .C(net5443),
    .Y(_15073_));
 XOR2x2_ASAP7_75t_R _23363_ (.A(_00661_),
    .B(_00693_),
    .Y(_15074_));
 XOR2x2_ASAP7_75t_R _23364_ (.A(_12238_),
    .B(_00597_),
    .Y(_15075_));
 XNOR2x2_ASAP7_75t_R _23365_ (.A(_15074_),
    .B(_15075_),
    .Y(_15076_));
 NOR2x1_ASAP7_75t_R _23366_ (.A(net6654),
    .B(_00519_),
    .Y(_15077_));
 AO21x1_ASAP7_75t_R _23367_ (.A1(_15076_),
    .A2(net6653),
    .B(_15077_),
    .Y(_15078_));
 XNOR2x2_ASAP7_75t_R _23368_ (.A(_00916_),
    .B(_15078_),
    .Y(_15079_));
 INVx1_ASAP7_75t_R _23369_ (.A(_15079_),
    .Y(_15080_));
 OAI21x1_ASAP7_75t_R _23371_ (.A1(_15066_),
    .A2(_15073_),
    .B(net5750),
    .Y(_15082_));
 NOR2x1_ASAP7_75t_R _23372_ (.A(_15082_),
    .B(_15054_),
    .Y(_15083_));
 NAND2x2_ASAP7_75t_R _23373_ (.A(net5778),
    .B(net5451),
    .Y(_15084_));
 NAND2x1_ASAP7_75t_R _23374_ (.A(net5763),
    .B(_15084_),
    .Y(_15085_));
 NAND2x1_ASAP7_75t_R _23375_ (.A(net5452),
    .B(net6179),
    .Y(_15086_));
 NOR2x1_ASAP7_75t_R _23376_ (.A(net5450),
    .B(_15086_),
    .Y(_15087_));
 AOI21x1_ASAP7_75t_R _23379_ (.A1(net5769),
    .A2(net5158),
    .B(net5154),
    .Y(_15090_));
 OAI21x1_ASAP7_75t_R _23380_ (.A1(_15085_),
    .A2(_15087_),
    .B(_15090_),
    .Y(_15091_));
 INVx1_ASAP7_75t_R _23381_ (.A(_15091_),
    .Y(_15092_));
 INVx1_ASAP7_75t_R _23382_ (.A(_01196_),
    .Y(_15093_));
 OAI21x1_ASAP7_75t_R _23383_ (.A1(net5779),
    .A2(net6177),
    .B(_15093_),
    .Y(_15094_));
 INVx1_ASAP7_75t_R _23384_ (.A(_15094_),
    .Y(_15095_));
 OAI21x1_ASAP7_75t_R _23386_ (.A1(_15095_),
    .A2(net5158),
    .B(net5772),
    .Y(_15097_));
 INVx1_ASAP7_75t_R _23387_ (.A(_15097_),
    .Y(_15098_));
 NAND2x1_ASAP7_75t_R _23388_ (.A(net5255),
    .B(_14974_),
    .Y(_15099_));
 AO21x1_ASAP7_75t_R _23390_ (.A1(net5003),
    .A2(net5760),
    .B(net5443),
    .Y(_15101_));
 XNOR2x2_ASAP7_75t_R _23391_ (.A(_00915_),
    .B(_15050_),
    .Y(_15102_));
 OAI21x1_ASAP7_75t_R _23393_ (.A1(_15098_),
    .A2(_15101_),
    .B(net5748),
    .Y(_15104_));
 OAI21x1_ASAP7_75t_R _23395_ (.A1(_15092_),
    .A2(_15104_),
    .B(net6174),
    .Y(_15106_));
 INVx1_ASAP7_75t_R _23396_ (.A(net5283),
    .Y(_15107_));
 OAI21x1_ASAP7_75t_R _23398_ (.A1(_15107_),
    .A2(net5450),
    .B(net5763),
    .Y(_15109_));
 INVx1_ASAP7_75t_R _23399_ (.A(_15109_),
    .Y(_15110_));
 OAI21x1_ASAP7_75t_R _23400_ (.A1(net5777),
    .A2(net6176),
    .B(_01189_),
    .Y(_15111_));
 INVx1_ASAP7_75t_R _23401_ (.A(_15111_),
    .Y(_15112_));
 OA21x2_ASAP7_75t_R _23403_ (.A1(_15055_),
    .A2(_15112_),
    .B(net5769),
    .Y(_15114_));
 OAI21x1_ASAP7_75t_R _23405_ (.A1(_15110_),
    .A2(_15114_),
    .B(net5154),
    .Y(_15116_));
 NOR2x1_ASAP7_75t_R _23406_ (.A(net6178),
    .B(net5451),
    .Y(_15117_));
 NOR2x1_ASAP7_75t_R _23407_ (.A(net5004),
    .B(net5444),
    .Y(_15118_));
 OA21x2_ASAP7_75t_R _23409_ (.A1(_15117_),
    .A2(_15118_),
    .B(net5776),
    .Y(_15120_));
 NOR2x1_ASAP7_75t_R _23410_ (.A(net5778),
    .B(_14967_),
    .Y(_15121_));
 NOR2x1_ASAP7_75t_R _23412_ (.A(_15068_),
    .B(net5444),
    .Y(_15123_));
 OA21x2_ASAP7_75t_R _23413_ (.A1(net5145),
    .A2(_15123_),
    .B(net5759),
    .Y(_15124_));
 OAI21x1_ASAP7_75t_R _23416_ (.A1(_15120_),
    .A2(_15124_),
    .B(net5443),
    .Y(_15127_));
 AOI21x1_ASAP7_75t_R _23419_ (.A1(_15116_),
    .A2(_15127_),
    .B(net5749),
    .Y(_15130_));
 XOR2x2_ASAP7_75t_R _23420_ (.A(_00661_),
    .B(net6580),
    .Y(_15131_));
 XOR2x2_ASAP7_75t_R _23421_ (.A(_15131_),
    .B(net6427),
    .Y(_15132_));
 XOR2x2_ASAP7_75t_R _23422_ (.A(net6631),
    .B(net6607),
    .Y(_15133_));
 XOR2x2_ASAP7_75t_R _23423_ (.A(_15132_),
    .B(_15133_),
    .Y(_15134_));
 NOR2x1_ASAP7_75t_R _23424_ (.A(net6668),
    .B(_00518_),
    .Y(_15135_));
 AO21x1_ASAP7_75t_R _23425_ (.A1(_15134_),
    .A2(net6660),
    .B(_15135_),
    .Y(_15136_));
 XOR2x2_ASAP7_75t_R _23426_ (.A(_15136_),
    .B(net6485),
    .Y(_15137_));
 INVx1_ASAP7_75t_R _23427_ (.A(_15137_),
    .Y(_15138_));
 OAI21x1_ASAP7_75t_R _23428_ (.A1(_15106_),
    .A2(_15130_),
    .B(_15138_),
    .Y(_15139_));
 INVx1_ASAP7_75t_R _23430_ (.A(_01198_),
    .Y(_15141_));
 NOR2x1_ASAP7_75t_R _23431_ (.A(_15141_),
    .B(_14974_),
    .Y(_15142_));
 NAND2x1_ASAP7_75t_R _23432_ (.A(net5761),
    .B(_15099_),
    .Y(_15143_));
 NOR2x1_ASAP7_75t_R _23433_ (.A(net4673),
    .B(_15143_),
    .Y(_15144_));
 OAI21x1_ASAP7_75t_R _23434_ (.A1(net6179),
    .A2(net5447),
    .B(net5778),
    .Y(_15145_));
 AO21x1_ASAP7_75t_R _23435_ (.A1(_15145_),
    .A2(net5767),
    .B(net5443),
    .Y(_15146_));
 NOR2x1_ASAP7_75t_R _23436_ (.A(_15144_),
    .B(_15146_),
    .Y(_15147_));
 AO21x1_ASAP7_75t_R _23438_ (.A1(_15084_),
    .A2(net5766),
    .B(net5155),
    .Y(_15149_));
 NOR2x1_ASAP7_75t_R _23439_ (.A(net5447),
    .B(net5440),
    .Y(_15150_));
 NOR2x1_ASAP7_75t_R _23440_ (.A(_15109_),
    .B(_15150_),
    .Y(_15151_));
 OAI21x1_ASAP7_75t_R _23442_ (.A1(_15149_),
    .A2(_15151_),
    .B(net5752),
    .Y(_15153_));
 OAI21x1_ASAP7_75t_R _23443_ (.A1(_15147_),
    .A2(_15153_),
    .B(net6174),
    .Y(_15154_));
 NOR2x1_ASAP7_75t_R _23444_ (.A(net6179),
    .B(net5447),
    .Y(_15155_));
 OA21x2_ASAP7_75t_R _23445_ (.A1(_15055_),
    .A2(_15155_),
    .B(net5776),
    .Y(_15156_));
 OAI21x1_ASAP7_75t_R _23446_ (.A1(_15087_),
    .A2(_15085_),
    .B(net5442),
    .Y(_15157_));
 OAI21x1_ASAP7_75t_R _23447_ (.A1(_15156_),
    .A2(_15157_),
    .B(net5749),
    .Y(_15158_));
 XNOR2x2_ASAP7_75t_R _23450_ (.A(_14926_),
    .B(net6488),
    .Y(_15161_));
 NOR2x1_ASAP7_75t_R _23452_ (.A(net6172),
    .B(net5448),
    .Y(_15162_));
 AO21x1_ASAP7_75t_R _23453_ (.A1(net5450),
    .A2(net5440),
    .B(net5143),
    .Y(_15163_));
 NAND2x1_ASAP7_75t_R _23454_ (.A(net5061),
    .B(net5445),
    .Y(_15164_));
 INVx1_ASAP7_75t_R _23455_ (.A(_15164_),
    .Y(_15165_));
 OAI21x1_ASAP7_75t_R _23457_ (.A1(_15165_),
    .A2(_15085_),
    .B(net5152),
    .Y(_15167_));
 AOI21x1_ASAP7_75t_R _23458_ (.A1(net5766),
    .A2(_15163_),
    .B(_15167_),
    .Y(_15168_));
 NOR2x1_ASAP7_75t_R _23459_ (.A(_15158_),
    .B(_15168_),
    .Y(_15169_));
 OAI21x1_ASAP7_75t_R _23460_ (.A1(_15154_),
    .A2(_15169_),
    .B(net6173),
    .Y(_15170_));
 NAND2x1_ASAP7_75t_R _23461_ (.A(net5778),
    .B(net6172),
    .Y(_15171_));
 INVx1_ASAP7_75t_R _23462_ (.A(_15171_),
    .Y(_15172_));
 NAND2x1_ASAP7_75t_R _23463_ (.A(net5452),
    .B(net5447),
    .Y(_15173_));
 NAND2x1_ASAP7_75t_R _23464_ (.A(net5767),
    .B(_15173_),
    .Y(_15174_));
 NOR2x1_ASAP7_75t_R _23465_ (.A(_15172_),
    .B(_15174_),
    .Y(_15175_));
 INVx1_ASAP7_75t_R _23466_ (.A(_15175_),
    .Y(_15176_));
 OAI21x1_ASAP7_75t_R _23467_ (.A1(net6172),
    .A2(net5452),
    .B(net5763),
    .Y(_15177_));
 OA21x2_ASAP7_75t_R _23469_ (.A1(_15177_),
    .A2(_14995_),
    .B(net5148),
    .Y(_15179_));
 NAND2x1_ASAP7_75t_R _23470_ (.A(_15176_),
    .B(_15179_),
    .Y(_15180_));
 OAI21x1_ASAP7_75t_R _23472_ (.A1(net5779),
    .A2(net6177),
    .B(_01195_),
    .Y(_15182_));
 NAND2x1_ASAP7_75t_R _23473_ (.A(_15111_),
    .B(_15182_),
    .Y(_15183_));
 AOI21x1_ASAP7_75t_R _23474_ (.A1(net5763),
    .A2(_15183_),
    .B(net5148),
    .Y(_15184_));
 OAI21x1_ASAP7_75t_R _23475_ (.A1(net5779),
    .A2(net6177),
    .B(_15034_),
    .Y(_15185_));
 INVx2_ASAP7_75t_R _23476_ (.A(_15185_),
    .Y(_15186_));
 AOI21x1_ASAP7_75t_R _23477_ (.A1(net6178),
    .A2(net5452),
    .B(net5445),
    .Y(_15187_));
 OAI21x1_ASAP7_75t_R _23478_ (.A1(_15186_),
    .A2(net5140),
    .B(net5764),
    .Y(_15188_));
 AOI21x1_ASAP7_75t_R _23479_ (.A1(_15184_),
    .A2(_15188_),
    .B(net5748),
    .Y(_15189_));
 NOR2x1_ASAP7_75t_R _23480_ (.A(net6172),
    .B(_14974_),
    .Y(_15190_));
 NAND2x1p5_ASAP7_75t_R _23481_ (.A(net5764),
    .B(_15185_),
    .Y(_15191_));
 NAND2x1_ASAP7_75t_R _23482_ (.A(net5255),
    .B(net5448),
    .Y(_15192_));
 AOI21x1_ASAP7_75t_R _23484_ (.A1(net5756),
    .A2(_15192_),
    .B(net5443),
    .Y(_15194_));
 OAI21x1_ASAP7_75t_R _23485_ (.A1(net5138),
    .A2(net4570),
    .B(_15194_),
    .Y(_15195_));
 AOI21x1_ASAP7_75t_R _23486_ (.A1(_15111_),
    .A2(net4750),
    .B(net5764),
    .Y(_15196_));
 NAND2x1_ASAP7_75t_R _23487_ (.A(net5063),
    .B(net5448),
    .Y(_15197_));
 AOI21x1_ASAP7_75t_R _23488_ (.A1(net5156),
    .A2(net4899),
    .B(net5756),
    .Y(_15198_));
 OAI21x1_ASAP7_75t_R _23489_ (.A1(_15196_),
    .A2(_15198_),
    .B(net5443),
    .Y(_15199_));
 AOI21x1_ASAP7_75t_R _23490_ (.A1(_15195_),
    .A2(_15199_),
    .B(_15051_),
    .Y(_15200_));
 AOI211x1_ASAP7_75t_R _23491_ (.A1(_15180_),
    .A2(_15189_),
    .B(_15200_),
    .C(net6174),
    .Y(_15201_));
 OAI22x1_ASAP7_75t_R _23492_ (.A1(_15083_),
    .A2(_15139_),
    .B1(_15170_),
    .B2(_15201_),
    .Y(_00080_));
 NAND2x1_ASAP7_75t_R _23494_ (.A(_01205_),
    .B(net5757),
    .Y(_15203_));
 AO21x1_ASAP7_75t_R _23495_ (.A1(_15203_),
    .A2(net5443),
    .B(net5752),
    .Y(_15204_));
 NOR2x1_ASAP7_75t_R _23496_ (.A(net5452),
    .B(net5449),
    .Y(_15205_));
 OAI21x1_ASAP7_75t_R _23497_ (.A1(_01189_),
    .A2(net5445),
    .B(net5764),
    .Y(_15206_));
 NOR2x1_ASAP7_75t_R _23498_ (.A(net5137),
    .B(_15206_),
    .Y(_15207_));
 AOI21x1_ASAP7_75t_R _23499_ (.A1(net6178),
    .A2(net5452),
    .B(net5449),
    .Y(_15208_));
 NAND2x1_ASAP7_75t_R _23500_ (.A(net5761),
    .B(_15208_),
    .Y(_15209_));
 NOR2x1_ASAP7_75t_R _23501_ (.A(net5447),
    .B(net5767),
    .Y(_15210_));
 AOI21x1_ASAP7_75t_R _23502_ (.A1(net5440),
    .A2(net5136),
    .B(net5443),
    .Y(_15211_));
 NAND2x1_ASAP7_75t_R _23503_ (.A(_15209_),
    .B(_15211_),
    .Y(_15212_));
 NOR2x1_ASAP7_75t_R _23504_ (.A(net5778),
    .B(net6172),
    .Y(_15213_));
 NAND2x1_ASAP7_75t_R _23505_ (.A(net5444),
    .B(_15213_),
    .Y(_15214_));
 AOI21x1_ASAP7_75t_R _23506_ (.A1(_15069_),
    .A2(_15214_),
    .B(net5151),
    .Y(_15215_));
 INVx1_ASAP7_75t_R _23507_ (.A(_15215_),
    .Y(_15216_));
 OAI21x1_ASAP7_75t_R _23508_ (.A1(_15207_),
    .A2(_15212_),
    .B(_15216_),
    .Y(_15217_));
 NOR2x1_ASAP7_75t_R _23509_ (.A(net5139),
    .B(net4900),
    .Y(_15218_));
 NOR2x1_ASAP7_75t_R _23510_ (.A(net5443),
    .B(_15051_),
    .Y(_15219_));
 NOR2x1_ASAP7_75t_R _23511_ (.A(net5283),
    .B(net5451),
    .Y(_15220_));
 OAI21x1_ASAP7_75t_R _23512_ (.A1(_15190_),
    .A2(_15220_),
    .B(net5763),
    .Y(_15221_));
 NAND2x1_ASAP7_75t_R _23513_ (.A(_15219_),
    .B(_15221_),
    .Y(_15222_));
 OAI21x1_ASAP7_75t_R _23514_ (.A1(_15218_),
    .A2(_15222_),
    .B(_15080_),
    .Y(_15223_));
 AOI21x1_ASAP7_75t_R _23515_ (.A1(_15204_),
    .A2(_15217_),
    .B(_15223_),
    .Y(_15224_));
 AO21x1_ASAP7_75t_R _23516_ (.A1(net5156),
    .A2(net4753),
    .B(net5766),
    .Y(_15225_));
 OAI21x1_ASAP7_75t_R _23517_ (.A1(_14995_),
    .A2(_15055_),
    .B(net5766),
    .Y(_15226_));
 AOI21x1_ASAP7_75t_R _23518_ (.A1(_15225_),
    .A2(_15226_),
    .B(net5443),
    .Y(_15227_));
 OAI21x1_ASAP7_75t_R _23519_ (.A1(_15112_),
    .A2(net5137),
    .B(net5766),
    .Y(_15228_));
 AOI21x1_ASAP7_75t_R _23520_ (.A1(_15228_),
    .A2(_15221_),
    .B(_15037_),
    .Y(_15229_));
 OAI21x1_ASAP7_75t_R _23521_ (.A1(_15227_),
    .A2(_15229_),
    .B(net5752),
    .Y(_15230_));
 OA21x2_ASAP7_75t_R _23522_ (.A1(net6177),
    .A2(net5779),
    .B(net5255),
    .Y(_15231_));
 OAI21x1_ASAP7_75t_R _23524_ (.A1(_15231_),
    .A2(_15187_),
    .B(net5758),
    .Y(_15233_));
 OAI21x1_ASAP7_75t_R _23525_ (.A1(net5061),
    .A2(net5451),
    .B(_15004_),
    .Y(_15234_));
 AOI21x1_ASAP7_75t_R _23526_ (.A1(net5770),
    .A2(_15234_),
    .B(net5443),
    .Y(_15235_));
 NAND2x1_ASAP7_75t_R _23527_ (.A(_15233_),
    .B(_15235_),
    .Y(_15236_));
 OAI21x1_ASAP7_75t_R _23528_ (.A1(_14995_),
    .A2(_15208_),
    .B(net5768),
    .Y(_15237_));
 NOR2x1p5_ASAP7_75t_R _23529_ (.A(net5776),
    .B(_15231_),
    .Y(_15238_));
 NOR2x1_ASAP7_75t_R _23530_ (.A(net5154),
    .B(_15238_),
    .Y(_15239_));
 AOI21x1_ASAP7_75t_R _23531_ (.A1(_15237_),
    .A2(_15239_),
    .B(net5752),
    .Y(_15240_));
 NAND2x1_ASAP7_75t_R _23532_ (.A(_15236_),
    .B(_15240_),
    .Y(_15241_));
 AOI21x1_ASAP7_75t_R _23533_ (.A1(_15230_),
    .A2(_15241_),
    .B(net5750),
    .Y(_15242_));
 OAI21x1_ASAP7_75t_R _23534_ (.A1(_15224_),
    .A2(_15242_),
    .B(net6173),
    .Y(_15243_));
 OAI21x1_ASAP7_75t_R _23536_ (.A1(net5002),
    .A2(net5158),
    .B(net5755),
    .Y(_15245_));
 OAI21x1_ASAP7_75t_R _23537_ (.A1(net4904),
    .A2(_14995_),
    .B(net5775),
    .Y(_15246_));
 AOI21x1_ASAP7_75t_R _23538_ (.A1(_15245_),
    .A2(_15246_),
    .B(net5443),
    .Y(_15247_));
 OAI21x1_ASAP7_75t_R _23539_ (.A1(net5438),
    .A2(net5137),
    .B(net5755),
    .Y(_15248_));
 OAI21x1_ASAP7_75t_R _23540_ (.A1(net5145),
    .A2(_15118_),
    .B(net5772),
    .Y(_15249_));
 AOI21x1_ASAP7_75t_R _23541_ (.A1(_15248_),
    .A2(_15249_),
    .B(net5150),
    .Y(_15250_));
 OAI21x1_ASAP7_75t_R _23542_ (.A1(_15247_),
    .A2(_15250_),
    .B(net5748),
    .Y(_15251_));
 AOI21x1_ASAP7_75t_R _23543_ (.A1(net5771),
    .A2(_15220_),
    .B(net5151),
    .Y(_15252_));
 AOI21x1_ASAP7_75t_R _23544_ (.A1(_15252_),
    .A2(_15233_),
    .B(net5748),
    .Y(_15253_));
 NAND2x1_ASAP7_75t_R _23545_ (.A(net5764),
    .B(_15208_),
    .Y(_15254_));
 NAND2x1_ASAP7_75t_R _23546_ (.A(net6172),
    .B(net5445),
    .Y(_15255_));
 NOR2x1_ASAP7_75t_R _23547_ (.A(net5764),
    .B(_15142_),
    .Y(_15256_));
 AOI21x1_ASAP7_75t_R _23548_ (.A1(net5134),
    .A2(_15256_),
    .B(net5443),
    .Y(_15257_));
 NAND2x1_ASAP7_75t_R _23549_ (.A(_15254_),
    .B(_15257_),
    .Y(_15258_));
 NAND2x1_ASAP7_75t_R _23550_ (.A(_15253_),
    .B(_15258_),
    .Y(_15259_));
 AOI21x1_ASAP7_75t_R _23551_ (.A1(_15251_),
    .A2(_15259_),
    .B(net5750),
    .Y(_15260_));
 OAI21x1_ASAP7_75t_R _23552_ (.A1(net5061),
    .A2(net5451),
    .B(net4755),
    .Y(_15261_));
 AOI21x1_ASAP7_75t_R _23553_ (.A1(net5759),
    .A2(_15261_),
    .B(net5154),
    .Y(_15262_));
 NAND2x1_ASAP7_75t_R _23554_ (.A(_14991_),
    .B(_15262_),
    .Y(_15263_));
 AOI21x1_ASAP7_75t_R _23555_ (.A1(net5774),
    .A2(net5158),
    .B(net5443),
    .Y(_15264_));
 OA21x2_ASAP7_75t_R _23556_ (.A1(_15190_),
    .A2(net5774),
    .B(net5134),
    .Y(_15265_));
 AOI21x1_ASAP7_75t_R _23557_ (.A1(_15264_),
    .A2(_15265_),
    .B(net5751),
    .Y(_15266_));
 NAND2x1_ASAP7_75t_R _23558_ (.A(_15263_),
    .B(_15266_),
    .Y(_15267_));
 NOR2x1_ASAP7_75t_R _23559_ (.A(net5001),
    .B(_15085_),
    .Y(_15268_));
 OA21x2_ASAP7_75t_R _23560_ (.A1(_15107_),
    .A2(net5450),
    .B(net5776),
    .Y(_15269_));
 NAND2x1_ASAP7_75t_R _23561_ (.A(net5452),
    .B(net5449),
    .Y(_15270_));
 AO21x1_ASAP7_75t_R _23562_ (.A1(_15269_),
    .A2(_15270_),
    .B(net5442),
    .Y(_15271_));
 NAND2x1_ASAP7_75t_R _23563_ (.A(net6179),
    .B(net5446),
    .Y(_15272_));
 NAND3x1_ASAP7_75t_R _23564_ (.A(_15272_),
    .B(net5439),
    .C(net5765),
    .Y(_15273_));
 AOI21x1_ASAP7_75t_R _23565_ (.A1(net5440),
    .A2(net5136),
    .B(net5154),
    .Y(_15274_));
 AOI21x1_ASAP7_75t_R _23566_ (.A1(_15273_),
    .A2(_15274_),
    .B(net5749),
    .Y(_15275_));
 OAI21x1_ASAP7_75t_R _23567_ (.A1(_15268_),
    .A2(_15271_),
    .B(_15275_),
    .Y(_15276_));
 AOI21x1_ASAP7_75t_R _23568_ (.A1(_15267_),
    .A2(_15276_),
    .B(net6174),
    .Y(_15277_));
 OAI21x1_ASAP7_75t_R _23569_ (.A1(_15260_),
    .A2(_15277_),
    .B(_15138_),
    .Y(_15278_));
 NAND2x1_ASAP7_75t_R _23570_ (.A(_15243_),
    .B(_15278_),
    .Y(_00081_));
 NAND2x1_ASAP7_75t_R _23571_ (.A(net5753),
    .B(_15192_),
    .Y(_15279_));
 OA21x2_ASAP7_75t_R _23572_ (.A1(_01203_),
    .A2(net5753),
    .B(_15051_),
    .Y(_15280_));
 OA21x2_ASAP7_75t_R _23573_ (.A1(net5146),
    .A2(_15279_),
    .B(_15280_),
    .Y(_15281_));
 AO21x1_ASAP7_75t_R _23574_ (.A1(_01205_),
    .A2(net5765),
    .B(_15051_),
    .Y(_15282_));
 NAND2x1_ASAP7_75t_R _23575_ (.A(net5763),
    .B(_15171_),
    .Y(_15283_));
 NOR2x1_ASAP7_75t_R _23576_ (.A(net5143),
    .B(_15283_),
    .Y(_15284_));
 OAI21x1_ASAP7_75t_R _23578_ (.A1(_15282_),
    .A2(_15284_),
    .B(net6174),
    .Y(_15286_));
 OAI21x1_ASAP7_75t_R _23579_ (.A1(net5444),
    .A2(net5441),
    .B(net5776),
    .Y(_15287_));
 NAND2x1_ASAP7_75t_R _23580_ (.A(_01202_),
    .B(net5753),
    .Y(_15288_));
 NAND3x1_ASAP7_75t_R _23581_ (.A(_15287_),
    .B(_15102_),
    .C(_15288_),
    .Y(_15289_));
 OAI21x1_ASAP7_75t_R _23582_ (.A1(_15186_),
    .A2(net5158),
    .B(net5753),
    .Y(_15290_));
 NAND2x1_ASAP7_75t_R _23583_ (.A(net5764),
    .B(_14993_),
    .Y(_15291_));
 AND2x2_ASAP7_75t_R _23584_ (.A(_15291_),
    .B(_15051_),
    .Y(_15292_));
 AOI21x1_ASAP7_75t_R _23585_ (.A1(_15290_),
    .A2(_15292_),
    .B(net6174),
    .Y(_15293_));
 AOI21x1_ASAP7_75t_R _23586_ (.A1(_15289_),
    .A2(_15293_),
    .B(net5149),
    .Y(_15294_));
 OAI21x1_ASAP7_75t_R _23587_ (.A1(_15281_),
    .A2(_15286_),
    .B(_15294_),
    .Y(_15295_));
 OAI21x1_ASAP7_75t_R _23588_ (.A1(net5778),
    .A2(net5444),
    .B(net6178),
    .Y(_15296_));
 NAND2x1_ASAP7_75t_R _23589_ (.A(net5753),
    .B(_15296_),
    .Y(_15297_));
 OA21x2_ASAP7_75t_R _23590_ (.A1(_01207_),
    .A2(net5753),
    .B(_15102_),
    .Y(_15298_));
 AOI21x1_ASAP7_75t_R _23591_ (.A1(_15297_),
    .A2(_15298_),
    .B(net6174),
    .Y(_15299_));
 AND2x2_ASAP7_75t_R _23592_ (.A(net5285),
    .B(_01193_),
    .Y(_15300_));
 NOR2x1_ASAP7_75t_R _23593_ (.A(_15300_),
    .B(net5448),
    .Y(_15301_));
 OAI21x1_ASAP7_75t_R _23594_ (.A1(_15301_),
    .A2(net5140),
    .B(net5753),
    .Y(_15302_));
 AOI21x1_ASAP7_75t_R _23595_ (.A1(_15069_),
    .A2(_15214_),
    .B(net5748),
    .Y(_15303_));
 NAND2x1_ASAP7_75t_R _23596_ (.A(_15302_),
    .B(_15303_),
    .Y(_15304_));
 AOI21x1_ASAP7_75t_R _23597_ (.A1(_15299_),
    .A2(_15304_),
    .B(net5443),
    .Y(_15305_));
 NAND2x1_ASAP7_75t_R _23598_ (.A(net6172),
    .B(net5451),
    .Y(_15306_));
 NAND2x1_ASAP7_75t_R _23599_ (.A(net5763),
    .B(_15306_),
    .Y(_15307_));
 NOR2x1_ASAP7_75t_R _23600_ (.A(net5753),
    .B(net5143),
    .Y(_15308_));
 AOI21x1_ASAP7_75t_R _23601_ (.A1(net4754),
    .A2(_15308_),
    .B(_15102_),
    .Y(_15309_));
 OAI21x1_ASAP7_75t_R _23602_ (.A1(net5137),
    .A2(net4898),
    .B(_15309_),
    .Y(_15310_));
 NAND2x1_ASAP7_75t_R _23603_ (.A(_15111_),
    .B(_15272_),
    .Y(_15311_));
 AOI21x1_ASAP7_75t_R _23604_ (.A1(net4753),
    .A2(_15182_),
    .B(net5764),
    .Y(_15312_));
 AOI21x1_ASAP7_75t_R _23605_ (.A1(net5764),
    .A2(_15311_),
    .B(_15312_),
    .Y(_15313_));
 AOI21x1_ASAP7_75t_R _23606_ (.A1(_15102_),
    .A2(_15313_),
    .B(_15080_),
    .Y(_15314_));
 NAND2x1_ASAP7_75t_R _23607_ (.A(_15310_),
    .B(_15314_),
    .Y(_15315_));
 AOI21x1_ASAP7_75t_R _23608_ (.A1(_15305_),
    .A2(_15315_),
    .B(net6173),
    .Y(_15316_));
 NAND2x1_ASAP7_75t_R _23609_ (.A(_15295_),
    .B(_15316_),
    .Y(_15317_));
 OAI21x1_ASAP7_75t_R _23610_ (.A1(net5777),
    .A2(net6176),
    .B(_15141_),
    .Y(_15318_));
 AO21x1_ASAP7_75t_R _23611_ (.A1(net4674),
    .A2(_15318_),
    .B(net5754),
    .Y(_15319_));
 OAI21x1_ASAP7_75t_R _23612_ (.A1(net5144),
    .A2(net5157),
    .B(net5754),
    .Y(_15320_));
 AOI21x1_ASAP7_75t_R _23613_ (.A1(_15319_),
    .A2(_15320_),
    .B(net5443),
    .Y(_15321_));
 OAI21x1_ASAP7_75t_R _23614_ (.A1(net5143),
    .A2(net5157),
    .B(net5754),
    .Y(_15322_));
 AOI21x1_ASAP7_75t_R _23615_ (.A1(_15097_),
    .A2(_15322_),
    .B(net5150),
    .Y(_15323_));
 OAI21x1_ASAP7_75t_R _23616_ (.A1(_15321_),
    .A2(_15323_),
    .B(net5748),
    .Y(_15324_));
 OAI21x1_ASAP7_75t_R _23617_ (.A1(_15186_),
    .A2(_15118_),
    .B(net5754),
    .Y(_15325_));
 NOR2x1_ASAP7_75t_R _23618_ (.A(net5062),
    .B(net5444),
    .Y(_15326_));
 OAI21x1_ASAP7_75t_R _23619_ (.A1(_15121_),
    .A2(_15326_),
    .B(net5773),
    .Y(_15327_));
 AOI21x1_ASAP7_75t_R _23620_ (.A1(_15325_),
    .A2(_15327_),
    .B(net5151),
    .Y(_15328_));
 AOI211x1_ASAP7_75t_R _23621_ (.A1(net6172),
    .A2(net5448),
    .B(_15095_),
    .C(net5773),
    .Y(_15329_));
 NAND2x1_ASAP7_75t_R _23622_ (.A(_15318_),
    .B(net5776),
    .Y(_15330_));
 OAI21x1_ASAP7_75t_R _23623_ (.A1(net5144),
    .A2(_15330_),
    .B(net5151),
    .Y(_15331_));
 NOR2x1_ASAP7_75t_R _23624_ (.A(_15329_),
    .B(_15331_),
    .Y(_15332_));
 OAI21x1_ASAP7_75t_R _23625_ (.A1(_15328_),
    .A2(_15332_),
    .B(net5751),
    .Y(_15333_));
 AOI21x1_ASAP7_75t_R _23626_ (.A1(_15324_),
    .A2(_15333_),
    .B(_15080_),
    .Y(_15334_));
 OAI21x1_ASAP7_75t_R _23627_ (.A1(net4677),
    .A2(net5145),
    .B(net5755),
    .Y(_15335_));
 OAI21x1_ASAP7_75t_R _23628_ (.A1(_15186_),
    .A2(_15155_),
    .B(net5773),
    .Y(_15336_));
 AOI21x1_ASAP7_75t_R _23629_ (.A1(_15335_),
    .A2(_15336_),
    .B(net5443),
    .Y(_15337_));
 NOR2x1_ASAP7_75t_R _23630_ (.A(net5061),
    .B(net5448),
    .Y(_15338_));
 OAI21x1_ASAP7_75t_R _23631_ (.A1(_15338_),
    .A2(net5140),
    .B(net5753),
    .Y(_15339_));
 AOI21x1_ASAP7_75t_R _23632_ (.A1(_15287_),
    .A2(_15339_),
    .B(net5151),
    .Y(_15340_));
 OAI21x1_ASAP7_75t_R _23633_ (.A1(_15337_),
    .A2(_15340_),
    .B(net5751),
    .Y(_15341_));
 INVx1_ASAP7_75t_R _23634_ (.A(_15318_),
    .Y(_15342_));
 OAI21x1_ASAP7_75t_R _23635_ (.A1(_15342_),
    .A2(_15220_),
    .B(net5771),
    .Y(_15343_));
 AOI21x1_ASAP7_75t_R _23636_ (.A1(_15297_),
    .A2(_15343_),
    .B(net5443),
    .Y(_15344_));
 INVx2_ASAP7_75t_R _23637_ (.A(net4755),
    .Y(_15345_));
 OAI21x1_ASAP7_75t_R _23638_ (.A1(_15345_),
    .A2(net5143),
    .B(net5772),
    .Y(_15346_));
 OAI21x1_ASAP7_75t_R _23639_ (.A1(net5157),
    .A2(_14976_),
    .B(net5754),
    .Y(_15347_));
 AOI21x1_ASAP7_75t_R _23640_ (.A1(_15346_),
    .A2(_15347_),
    .B(net5150),
    .Y(_15348_));
 OAI21x1_ASAP7_75t_R _23641_ (.A1(_15344_),
    .A2(_15348_),
    .B(net5748),
    .Y(_15349_));
 AOI21x1_ASAP7_75t_R _23642_ (.A1(_15341_),
    .A2(_15349_),
    .B(net6174),
    .Y(_15350_));
 OAI21x1_ASAP7_75t_R _23643_ (.A1(_15334_),
    .A2(_15350_),
    .B(net6173),
    .Y(_15351_));
 NAND2x1_ASAP7_75t_R _23644_ (.A(_15317_),
    .B(_15351_),
    .Y(_00082_));
 NAND2x1_ASAP7_75t_R _23645_ (.A(net5754),
    .B(_15118_),
    .Y(_15352_));
 AO21x1_ASAP7_75t_R _23646_ (.A1(net5134),
    .A2(_15197_),
    .B(net5754),
    .Y(_15353_));
 AOI21x1_ASAP7_75t_R _23647_ (.A1(_15352_),
    .A2(_15353_),
    .B(net5751),
    .Y(_15354_));
 NOR2x1_ASAP7_75t_R _23648_ (.A(net5763),
    .B(_15099_),
    .Y(_15355_));
 AO21x1_ASAP7_75t_R _23649_ (.A1(net5751),
    .A2(_15355_),
    .B(_15071_),
    .Y(_15356_));
 OAI21x1_ASAP7_75t_R _23650_ (.A1(_15354_),
    .A2(_15356_),
    .B(net5151),
    .Y(_15357_));
 NOR2x1_ASAP7_75t_R _23651_ (.A(_15094_),
    .B(net5764),
    .Y(_15358_));
 NOR2x1_ASAP7_75t_R _23652_ (.A(_15102_),
    .B(_15358_),
    .Y(_15359_));
 AOI21x1_ASAP7_75t_R _23653_ (.A1(_15327_),
    .A2(_15359_),
    .B(net5151),
    .Y(_15360_));
 NAND2x1_ASAP7_75t_R _23654_ (.A(_15300_),
    .B(net5444),
    .Y(_15361_));
 NAND2x1_ASAP7_75t_R _23655_ (.A(net5754),
    .B(_15361_),
    .Y(_15362_));
 NAND2x1_ASAP7_75t_R _23656_ (.A(_15185_),
    .B(_15270_),
    .Y(_15363_));
 AOI21x1_ASAP7_75t_R _23657_ (.A1(net5764),
    .A2(_15363_),
    .B(_15051_),
    .Y(_15364_));
 OAI21x1_ASAP7_75t_R _23658_ (.A1(net4673),
    .A2(_15362_),
    .B(_15364_),
    .Y(_15365_));
 AOI21x1_ASAP7_75t_R _23659_ (.A1(_15360_),
    .A2(_15365_),
    .B(net6174),
    .Y(_15366_));
 NAND2x1_ASAP7_75t_R _23660_ (.A(_15357_),
    .B(_15366_),
    .Y(_15367_));
 AO21x1_ASAP7_75t_R _23661_ (.A1(net4751),
    .A2(_15318_),
    .B(net5758),
    .Y(_15368_));
 AOI21x1_ASAP7_75t_R _23662_ (.A1(net4674),
    .A2(_15084_),
    .B(net5768),
    .Y(_15369_));
 INVx1_ASAP7_75t_R _23663_ (.A(_15369_),
    .Y(_15370_));
 AOI21x1_ASAP7_75t_R _23664_ (.A1(_15368_),
    .A2(_15370_),
    .B(net5443),
    .Y(_15371_));
 AOI21x1_ASAP7_75t_R _23665_ (.A1(_15002_),
    .A2(_15273_),
    .B(net5154),
    .Y(_15372_));
 OAI21x1_ASAP7_75t_R _23666_ (.A1(_15371_),
    .A2(_15372_),
    .B(net5751),
    .Y(_15373_));
 NOR2x1_ASAP7_75t_R _23667_ (.A(_15121_),
    .B(_15330_),
    .Y(_15374_));
 AOI21x1_ASAP7_75t_R _23668_ (.A1(net5151),
    .A2(_15374_),
    .B(net5751),
    .Y(_15375_));
 OAI21x1_ASAP7_75t_R _23669_ (.A1(_15326_),
    .A2(_15301_),
    .B(net5754),
    .Y(_15376_));
 NAND2x1_ASAP7_75t_R _23670_ (.A(_15376_),
    .B(_15215_),
    .Y(_15377_));
 AOI21x1_ASAP7_75t_R _23671_ (.A1(_15375_),
    .A2(_15377_),
    .B(_15080_),
    .Y(_15378_));
 AOI21x1_ASAP7_75t_R _23672_ (.A1(_15373_),
    .A2(_15378_),
    .B(_15138_),
    .Y(_15379_));
 NAND2x1_ASAP7_75t_R _23673_ (.A(_15367_),
    .B(_15379_),
    .Y(_15380_));
 NAND2x1_ASAP7_75t_R _23674_ (.A(_15182_),
    .B(_15270_),
    .Y(_15381_));
 OAI22x1_ASAP7_75t_R _23675_ (.A1(_15279_),
    .A2(net4904),
    .B1(net4671),
    .B2(net5753),
    .Y(_15382_));
 OA21x2_ASAP7_75t_R _23676_ (.A1(_15191_),
    .A2(_15155_),
    .B(net5443),
    .Y(_15383_));
 OAI21x1_ASAP7_75t_R _23677_ (.A1(net5158),
    .A2(_15338_),
    .B(net5753),
    .Y(_15384_));
 AO21x1_ASAP7_75t_R _23678_ (.A1(_15383_),
    .A2(_15384_),
    .B(net6174),
    .Y(_15385_));
 AOI21x1_ASAP7_75t_R _23679_ (.A1(net5149),
    .A2(_15382_),
    .B(_15385_),
    .Y(_15386_));
 NAND2x1_ASAP7_75t_R _23680_ (.A(_15035_),
    .B(net5764),
    .Y(_15387_));
 OAI21x1_ASAP7_75t_R _23681_ (.A1(_15208_),
    .A2(_15387_),
    .B(net5443),
    .Y(_15388_));
 NOR2x1_ASAP7_75t_R _23682_ (.A(_15307_),
    .B(_15381_),
    .Y(_15389_));
 NOR2x1_ASAP7_75t_R _23683_ (.A(_15388_),
    .B(_15389_),
    .Y(_15390_));
 NOR2x1_ASAP7_75t_R _23684_ (.A(net5002),
    .B(_15123_),
    .Y(_15391_));
 OAI21x1_ASAP7_75t_R _23685_ (.A1(_14995_),
    .A2(_15177_),
    .B(net5154),
    .Y(_15392_));
 AOI21x1_ASAP7_75t_R _23686_ (.A1(net5776),
    .A2(_15391_),
    .B(_15392_),
    .Y(_15393_));
 OAI21x1_ASAP7_75t_R _23687_ (.A1(_15390_),
    .A2(_15393_),
    .B(net6174),
    .Y(_15394_));
 NAND2x1_ASAP7_75t_R _23688_ (.A(net5751),
    .B(_15394_),
    .Y(_15395_));
 NAND2x1_ASAP7_75t_R _23689_ (.A(net5447),
    .B(net5757),
    .Y(_15396_));
 OAI21x1_ASAP7_75t_R _23690_ (.A1(net5778),
    .A2(net5447),
    .B(net5443),
    .Y(_15397_));
 NOR2x1_ASAP7_75t_R _23691_ (.A(_15172_),
    .B(_15397_),
    .Y(_15398_));
 AOI21x1_ASAP7_75t_R _23692_ (.A1(_15396_),
    .A2(_15398_),
    .B(_15080_),
    .Y(_15399_));
 AO21x1_ASAP7_75t_R _23693_ (.A1(net5062),
    .A2(net5448),
    .B(_15191_),
    .Y(_15400_));
 NAND2x1_ASAP7_75t_R _23694_ (.A(_15257_),
    .B(_15400_),
    .Y(_15401_));
 NAND2x1_ASAP7_75t_R _23695_ (.A(_15401_),
    .B(_15399_),
    .Y(_15402_));
 OAI21x1_ASAP7_75t_R _23696_ (.A1(_15121_),
    .A2(_15190_),
    .B(net5767),
    .Y(_15403_));
 AOI21x1_ASAP7_75t_R _23697_ (.A1(_15194_),
    .A2(_15403_),
    .B(net6174),
    .Y(_15404_));
 AO21x1_ASAP7_75t_R _23698_ (.A1(_15270_),
    .A2(net5439),
    .B(net5757),
    .Y(_15405_));
 AOI21x1_ASAP7_75t_R _23699_ (.A1(net5133),
    .A2(_15238_),
    .B(_15037_),
    .Y(_15406_));
 NAND2x1_ASAP7_75t_R _23700_ (.A(_15405_),
    .B(_15406_),
    .Y(_15407_));
 AOI21x1_ASAP7_75t_R _23701_ (.A1(_15404_),
    .A2(_15407_),
    .B(_15051_),
    .Y(_15408_));
 AOI21x1_ASAP7_75t_R _23702_ (.A1(_15408_),
    .A2(_15402_),
    .B(net6173),
    .Y(_15409_));
 OAI21x1_ASAP7_75t_R _23703_ (.A1(_15395_),
    .A2(_15386_),
    .B(_15409_),
    .Y(_15410_));
 NAND2x1_ASAP7_75t_R _23704_ (.A(_15380_),
    .B(_15410_),
    .Y(_00083_));
 AO21x1_ASAP7_75t_R _23705_ (.A1(_15345_),
    .A2(net5755),
    .B(_15095_),
    .Y(_15411_));
 INVx1_ASAP7_75t_R _23706_ (.A(_15264_),
    .Y(_15412_));
 OAI21x1_ASAP7_75t_R _23707_ (.A1(_15411_),
    .A2(_15412_),
    .B(net5751),
    .Y(_15413_));
 AO21x1_ASAP7_75t_R _23708_ (.A1(_15261_),
    .A2(net5774),
    .B(net5154),
    .Y(_15414_));
 NOR2x1_ASAP7_75t_R _23709_ (.A(_15064_),
    .B(_15414_),
    .Y(_15415_));
 OAI21x1_ASAP7_75t_R _23710_ (.A1(_15413_),
    .A2(_15415_),
    .B(net5750),
    .Y(_15416_));
 INVx1_ASAP7_75t_R _23711_ (.A(_15343_),
    .Y(_15417_));
 NOR2x1_ASAP7_75t_R _23712_ (.A(net5147),
    .B(net4898),
    .Y(_15418_));
 OAI21x1_ASAP7_75t_R _23713_ (.A1(_15417_),
    .A2(_15418_),
    .B(net5153),
    .Y(_15419_));
 OA21x2_ASAP7_75t_R _23714_ (.A1(_15190_),
    .A2(net4904),
    .B(net5759),
    .Y(_15420_));
 INVx1_ASAP7_75t_R _23715_ (.A(_14991_),
    .Y(_15421_));
 OAI21x1_ASAP7_75t_R _23716_ (.A1(_15420_),
    .A2(_15421_),
    .B(net5443),
    .Y(_15422_));
 AOI21x1_ASAP7_75t_R _23717_ (.A1(_15419_),
    .A2(_15422_),
    .B(net5751),
    .Y(_15423_));
 OAI21x1_ASAP7_75t_R _23718_ (.A1(_15416_),
    .A2(_15423_),
    .B(_15138_),
    .Y(_15424_));
 OAI21x1_ASAP7_75t_R _23719_ (.A1(net5139),
    .A2(net4900),
    .B(net5749),
    .Y(_15425_));
 NOR2x1_ASAP7_75t_R _23720_ (.A(_15284_),
    .B(_15425_),
    .Y(_15426_));
 OA21x2_ASAP7_75t_R _23721_ (.A1(_15121_),
    .A2(_15155_),
    .B(net5757),
    .Y(_15427_));
 OAI21x1_ASAP7_75t_R _23722_ (.A1(net5137),
    .A2(_15206_),
    .B(net5752),
    .Y(_15428_));
 OAI21x1_ASAP7_75t_R _23723_ (.A1(_15427_),
    .A2(_15428_),
    .B(net5443),
    .Y(_15429_));
 OAI21x1_ASAP7_75t_R _23724_ (.A1(_15426_),
    .A2(_15429_),
    .B(net6174),
    .Y(_15430_));
 AO21x1_ASAP7_75t_R _23725_ (.A1(_15063_),
    .A2(_15070_),
    .B(net5749),
    .Y(_15431_));
 NAND2x1_ASAP7_75t_R _23726_ (.A(_15086_),
    .B(net5134),
    .Y(_15432_));
 AOI21x1_ASAP7_75t_R _23727_ (.A1(net5769),
    .A2(_15432_),
    .B(net5751),
    .Y(_15433_));
 OR3x1_ASAP7_75t_R _23728_ (.A(net5143),
    .B(_15112_),
    .C(net5769),
    .Y(_15434_));
 NAND2x1_ASAP7_75t_R _23729_ (.A(_15433_),
    .B(_15434_),
    .Y(_15435_));
 AOI21x1_ASAP7_75t_R _23730_ (.A1(_15431_),
    .A2(_15435_),
    .B(net5442),
    .Y(_15436_));
 NOR2x1_ASAP7_75t_R _23731_ (.A(_15430_),
    .B(_15436_),
    .Y(_15437_));
 NOR2x1_ASAP7_75t_R _23732_ (.A(_14995_),
    .B(_15177_),
    .Y(_15438_));
 OAI21x1_ASAP7_75t_R _23733_ (.A1(_15438_),
    .A2(_15114_),
    .B(net5442),
    .Y(_15439_));
 AO21x1_ASAP7_75t_R _23734_ (.A1(net5134),
    .A2(_15086_),
    .B(net5763),
    .Y(_15440_));
 INVx1_ASAP7_75t_R _23735_ (.A(_15440_),
    .Y(_15441_));
 NOR2x1_ASAP7_75t_R _23736_ (.A(net5145),
    .B(_15063_),
    .Y(_15442_));
 OAI21x1_ASAP7_75t_R _23737_ (.A1(_15441_),
    .A2(_15442_),
    .B(net5154),
    .Y(_15443_));
 AOI21x1_ASAP7_75t_R _23738_ (.A1(_15439_),
    .A2(_15443_),
    .B(net5751),
    .Y(_15444_));
 INVx1_ASAP7_75t_R _23739_ (.A(_01197_),
    .Y(_15445_));
 NOR2x1_ASAP7_75t_R _23740_ (.A(net4753),
    .B(net5776),
    .Y(_15446_));
 AOI21x1_ASAP7_75t_R _23741_ (.A1(_15445_),
    .A2(net5766),
    .B(_15446_),
    .Y(_15447_));
 OAI21x1_ASAP7_75t_R _23742_ (.A1(net5155),
    .A2(_15447_),
    .B(net5752),
    .Y(_15448_));
 OAI21x1_ASAP7_75t_R _23743_ (.A1(net5143),
    .A2(_15326_),
    .B(net5755),
    .Y(_15449_));
 INVx1_ASAP7_75t_R _23744_ (.A(_15449_),
    .Y(_15450_));
 NOR2x1_ASAP7_75t_R _23745_ (.A(net5762),
    .B(net5134),
    .Y(_15451_));
 OAI21x1_ASAP7_75t_R _23746_ (.A1(net5762),
    .A2(net5142),
    .B(net5155),
    .Y(_15452_));
 NOR3x1_ASAP7_75t_R _23747_ (.A(_15450_),
    .B(_15451_),
    .C(_15452_),
    .Y(_15453_));
 OAI21x1_ASAP7_75t_R _23748_ (.A1(_15448_),
    .A2(_15453_),
    .B(net5750),
    .Y(_15454_));
 NOR2x1_ASAP7_75t_R _23749_ (.A(_15444_),
    .B(_15454_),
    .Y(_15455_));
 AO21x1_ASAP7_75t_R _23750_ (.A1(net5445),
    .A2(net5438),
    .B(_15085_),
    .Y(_15456_));
 AOI21x1_ASAP7_75t_R _23751_ (.A1(net4752),
    .A2(_15269_),
    .B(net5152),
    .Y(_15457_));
 OA21x2_ASAP7_75t_R _23752_ (.A1(_15086_),
    .A2(net5445),
    .B(net5762),
    .Y(_15458_));
 NAND2x1_ASAP7_75t_R _23753_ (.A(net5284),
    .B(net5449),
    .Y(_15459_));
 AO21x1_ASAP7_75t_R _23754_ (.A1(_15459_),
    .A2(net5776),
    .B(net5442),
    .Y(_15460_));
 OAI21x1_ASAP7_75t_R _23755_ (.A1(_15458_),
    .A2(_15460_),
    .B(net5752),
    .Y(_15461_));
 AOI21x1_ASAP7_75t_R _23756_ (.A1(_15456_),
    .A2(_15457_),
    .B(_15461_),
    .Y(_15462_));
 AO21x1_ASAP7_75t_R _23757_ (.A1(_15155_),
    .A2(net5766),
    .B(net5443),
    .Y(_15463_));
 OAI21x1_ASAP7_75t_R _23758_ (.A1(_15155_),
    .A2(_15109_),
    .B(net4672),
    .Y(_15464_));
 NOR2x1_ASAP7_75t_R _23759_ (.A(_15463_),
    .B(_15464_),
    .Y(_15465_));
 AO21x1_ASAP7_75t_R _23760_ (.A1(net5761),
    .A2(net5450),
    .B(net5155),
    .Y(_15466_));
 NOR2x1_ASAP7_75t_R _23761_ (.A(net4673),
    .B(net4900),
    .Y(_15467_));
 OAI21x1_ASAP7_75t_R _23762_ (.A1(_15466_),
    .A2(_15467_),
    .B(net5749),
    .Y(_15468_));
 OAI21x1_ASAP7_75t_R _23763_ (.A1(_15465_),
    .A2(_15468_),
    .B(net6174),
    .Y(_15469_));
 OAI21x1_ASAP7_75t_R _23764_ (.A1(_15462_),
    .A2(_15469_),
    .B(net6173),
    .Y(_15470_));
 OAI22x1_ASAP7_75t_R _23765_ (.A1(_15424_),
    .A2(_15437_),
    .B1(_15455_),
    .B2(_15470_),
    .Y(_00084_));
 NOR2x1_ASAP7_75t_R _23766_ (.A(_15150_),
    .B(_15143_),
    .Y(_15471_));
 OAI21x1_ASAP7_75t_R _23767_ (.A1(net4902),
    .A2(_14974_),
    .B(net5764),
    .Y(_15472_));
 OAI21x1_ASAP7_75t_R _23768_ (.A1(_15117_),
    .A2(_15472_),
    .B(net5154),
    .Y(_15473_));
 NOR2x1_ASAP7_75t_R _23769_ (.A(_15471_),
    .B(_15473_),
    .Y(_15474_));
 AO21x1_ASAP7_75t_R _23770_ (.A1(net5761),
    .A2(net5452),
    .B(net5155),
    .Y(_15475_));
 OAI21x1_ASAP7_75t_R _23771_ (.A1(_15475_),
    .A2(_15175_),
    .B(net5752),
    .Y(_15476_));
 OAI21x1_ASAP7_75t_R _23772_ (.A1(_15474_),
    .A2(_15476_),
    .B(net6174),
    .Y(_15477_));
 NAND2x1_ASAP7_75t_R _23773_ (.A(net5776),
    .B(_15121_),
    .Y(_15478_));
 INVx1_ASAP7_75t_R _23774_ (.A(_15478_),
    .Y(_15479_));
 NOR2x1_ASAP7_75t_R _23775_ (.A(_15479_),
    .B(_15091_),
    .Y(_15480_));
 AO21x1_ASAP7_75t_R _23776_ (.A1(_15123_),
    .A2(net5759),
    .B(net5443),
    .Y(_15481_));
 OA21x2_ASAP7_75t_R _23777_ (.A1(_15208_),
    .A2(_15342_),
    .B(net5771),
    .Y(_15482_));
 OAI21x1_ASAP7_75t_R _23778_ (.A1(_15481_),
    .A2(_15482_),
    .B(net5748),
    .Y(_15483_));
 NOR2x1_ASAP7_75t_R _23779_ (.A(_15480_),
    .B(_15483_),
    .Y(_15484_));
 OAI21x1_ASAP7_75t_R _23780_ (.A1(_15477_),
    .A2(_15484_),
    .B(net6173),
    .Y(_15485_));
 NAND2x1_ASAP7_75t_R _23781_ (.A(net4903),
    .B(net5451),
    .Y(_15486_));
 OAI21x1_ASAP7_75t_R _23782_ (.A1(net4569),
    .A2(net4673),
    .B(net5151),
    .Y(_15487_));
 AO21x1_ASAP7_75t_R _23783_ (.A1(_15486_),
    .A2(net4749),
    .B(_15487_),
    .Y(_15488_));
 AO21x1_ASAP7_75t_R _23784_ (.A1(net5755),
    .A2(net5063),
    .B(net5151),
    .Y(_15489_));
 AO21x1_ASAP7_75t_R _23785_ (.A1(net5772),
    .A2(net5135),
    .B(_15489_),
    .Y(_15490_));
 AND2x2_ASAP7_75t_R _23786_ (.A(_15490_),
    .B(net5748),
    .Y(_15491_));
 OAI21x1_ASAP7_75t_R _23787_ (.A1(net4518),
    .A2(_15412_),
    .B(net5751),
    .Y(_15492_));
 INVx1_ASAP7_75t_R _23788_ (.A(_15287_),
    .Y(_15493_));
 AO21x1_ASAP7_75t_R _23789_ (.A1(_15361_),
    .A2(net5754),
    .B(net5151),
    .Y(_15494_));
 AOI21x1_ASAP7_75t_R _23790_ (.A1(_15214_),
    .A2(_15493_),
    .B(_15494_),
    .Y(_15495_));
 OAI21x1_ASAP7_75t_R _23791_ (.A1(_15492_),
    .A2(_15495_),
    .B(net5750),
    .Y(_15496_));
 AOI21x1_ASAP7_75t_R _23792_ (.A1(_15491_),
    .A2(_15488_),
    .B(_15496_),
    .Y(_15497_));
 AO21x1_ASAP7_75t_R _23793_ (.A1(net5003),
    .A2(net5776),
    .B(net5154),
    .Y(_15498_));
 OAI21x1_ASAP7_75t_R _23794_ (.A1(net4517),
    .A2(_15498_),
    .B(net5749),
    .Y(_15499_));
 AOI211x1_ASAP7_75t_R _23795_ (.A1(net5136),
    .A2(net5440),
    .B(_15269_),
    .C(net5442),
    .Y(_15500_));
 OAI21x1_ASAP7_75t_R _23796_ (.A1(_15499_),
    .A2(_15500_),
    .B(net6174),
    .Y(_15501_));
 NOR2x1_ASAP7_75t_R _23797_ (.A(net4673),
    .B(_15109_),
    .Y(_15502_));
 OAI21x1_ASAP7_75t_R _23798_ (.A1(_15502_),
    .A2(_15156_),
    .B(net5442),
    .Y(_15503_));
 OA21x2_ASAP7_75t_R _23799_ (.A1(_15055_),
    .A2(_15107_),
    .B(net5762),
    .Y(_15504_));
 NOR2x1_ASAP7_75t_R _23800_ (.A(_15472_),
    .B(net5146),
    .Y(_15505_));
 OAI21x1_ASAP7_75t_R _23801_ (.A1(_15504_),
    .A2(_15505_),
    .B(net5152),
    .Y(_15506_));
 AOI21x1_ASAP7_75t_R _23802_ (.A1(_15503_),
    .A2(_15506_),
    .B(net5749),
    .Y(_15507_));
 OAI21x1_ASAP7_75t_R _23803_ (.A1(_15501_),
    .A2(_15507_),
    .B(_15138_),
    .Y(_15508_));
 AOI21x1_ASAP7_75t_R _23804_ (.A1(_15486_),
    .A2(net5135),
    .B(net5775),
    .Y(_15509_));
 NAND2x1_ASAP7_75t_R _23805_ (.A(net5776),
    .B(_15084_),
    .Y(_15510_));
 OAI21x1_ASAP7_75t_R _23806_ (.A1(net5438),
    .A2(_15510_),
    .B(net5154),
    .Y(_15511_));
 OA21x2_ASAP7_75t_R _23807_ (.A1(net5769),
    .A2(net6179),
    .B(net5443),
    .Y(_15512_));
 AOI21x1_ASAP7_75t_R _23808_ (.A1(_15512_),
    .A2(_15440_),
    .B(net5749),
    .Y(_15513_));
 OAI21x1_ASAP7_75t_R _23809_ (.A1(_15509_),
    .A2(_15511_),
    .B(_15513_),
    .Y(_15514_));
 AND2x2_ASAP7_75t_R _23810_ (.A(_15330_),
    .B(net5443),
    .Y(_15515_));
 NAND2x1_ASAP7_75t_R _23811_ (.A(_15111_),
    .B(net4749),
    .Y(_15516_));
 AOI21x1_ASAP7_75t_R _23812_ (.A1(_15515_),
    .A2(_15516_),
    .B(net5751),
    .Y(_15517_));
 AND3x1_ASAP7_75t_R _23813_ (.A(_15272_),
    .B(_15459_),
    .C(net5776),
    .Y(_15518_));
 OAI21x1_ASAP7_75t_R _23814_ (.A1(_15446_),
    .A2(_15518_),
    .B(net5154),
    .Y(_15519_));
 NAND2x1_ASAP7_75t_R _23815_ (.A(_15517_),
    .B(_15519_),
    .Y(_15520_));
 AOI21x1_ASAP7_75t_R _23816_ (.A1(_15514_),
    .A2(_15520_),
    .B(net6174),
    .Y(_15521_));
 OAI22x1_ASAP7_75t_R _23817_ (.A1(_15497_),
    .A2(_15485_),
    .B1(_15508_),
    .B2(_15521_),
    .Y(_00085_));
 NOR2x1_ASAP7_75t_R _23818_ (.A(_15165_),
    .B(_15472_),
    .Y(_15522_));
 AOI211x1_ASAP7_75t_R _23819_ (.A1(net5759),
    .A2(net5141),
    .B(_15522_),
    .C(net4675),
    .Y(_15523_));
 NOR2x1_ASAP7_75t_R _23820_ (.A(_15095_),
    .B(net5158),
    .Y(_15524_));
 NOR2x1_ASAP7_75t_R _23821_ (.A(net5771),
    .B(net4677),
    .Y(_15525_));
 NAND2x1_ASAP7_75t_R _23822_ (.A(_15478_),
    .B(_15039_),
    .Y(_15526_));
 AO21x1_ASAP7_75t_R _23823_ (.A1(_15524_),
    .A2(_15525_),
    .B(_15526_),
    .Y(_15527_));
 OAI21x1_ASAP7_75t_R _23824_ (.A1(net5154),
    .A2(_15523_),
    .B(_15527_),
    .Y(_15528_));
 AO21x1_ASAP7_75t_R _23825_ (.A1(_15004_),
    .A2(net4674),
    .B(net5770),
    .Y(_15529_));
 AND3x1_ASAP7_75t_R _23826_ (.A(_15529_),
    .B(_15037_),
    .C(net4672),
    .Y(_15530_));
 NAND2x1_ASAP7_75t_R _23827_ (.A(_01200_),
    .B(_01206_),
    .Y(_15531_));
 AO21x1_ASAP7_75t_R _23828_ (.A1(net5764),
    .A2(_15531_),
    .B(net5148),
    .Y(_15532_));
 AND3x1_ASAP7_75t_R _23829_ (.A(net5133),
    .B(net5761),
    .C(net5440),
    .Y(_15533_));
 OAI21x1_ASAP7_75t_R _23830_ (.A1(_15532_),
    .A2(_15533_),
    .B(net5752),
    .Y(_15534_));
 OAI21x1_ASAP7_75t_R _23831_ (.A1(_15530_),
    .A2(_15534_),
    .B(net6174),
    .Y(_15535_));
 AOI21x1_ASAP7_75t_R _23832_ (.A1(net5749),
    .A2(_15528_),
    .B(_15535_),
    .Y(_15536_));
 AO21x1_ASAP7_75t_R _23833_ (.A1(net5002),
    .A2(net5772),
    .B(net5443),
    .Y(_15537_));
 AO21x1_ASAP7_75t_R _23834_ (.A1(_15287_),
    .A2(_15288_),
    .B(_15537_),
    .Y(_15538_));
 AND3x1_ASAP7_75t_R _23835_ (.A(_15459_),
    .B(net5776),
    .C(net4750),
    .Y(_15539_));
 AOI211x1_ASAP7_75t_R _23836_ (.A1(net5138),
    .A2(net5778),
    .B(_15117_),
    .C(net5768),
    .Y(_15540_));
 OAI21x1_ASAP7_75t_R _23837_ (.A1(_15539_),
    .A2(_15540_),
    .B(net5443),
    .Y(_15541_));
 AOI21x1_ASAP7_75t_R _23838_ (.A1(_15538_),
    .A2(_15541_),
    .B(net5749),
    .Y(_15542_));
 OA21x2_ASAP7_75t_R _23839_ (.A1(_15197_),
    .A2(net5763),
    .B(_15037_),
    .Y(_15543_));
 AO21x1_ASAP7_75t_R _23840_ (.A1(net5142),
    .A2(net6179),
    .B(net5766),
    .Y(_15544_));
 AO21x1_ASAP7_75t_R _23841_ (.A1(_15543_),
    .A2(_15544_),
    .B(net5752),
    .Y(_15545_));
 AND3x1_ASAP7_75t_R _23842_ (.A(_15361_),
    .B(net5768),
    .C(net4753),
    .Y(_15546_));
 AOI21x1_ASAP7_75t_R _23843_ (.A1(net5778),
    .A2(_15210_),
    .B(net5155),
    .Y(_15547_));
 OAI21x1_ASAP7_75t_R _23844_ (.A1(_14995_),
    .A2(_15177_),
    .B(_15547_),
    .Y(_15548_));
 NOR2x1_ASAP7_75t_R _23845_ (.A(_15546_),
    .B(_15548_),
    .Y(_15549_));
 OAI21x1_ASAP7_75t_R _23846_ (.A1(_15545_),
    .A2(_15549_),
    .B(net5750),
    .Y(_15550_));
 OAI21x1_ASAP7_75t_R _23847_ (.A1(_15542_),
    .A2(_15550_),
    .B(_15138_),
    .Y(_15551_));
 NAND2x1_ASAP7_75t_R _23848_ (.A(net6179),
    .B(net5449),
    .Y(_15552_));
 AOI21x1_ASAP7_75t_R _23849_ (.A1(net5757),
    .A2(_15552_),
    .B(net5443),
    .Y(_15553_));
 NAND2x1_ASAP7_75t_R _23850_ (.A(net5765),
    .B(_15145_),
    .Y(_15554_));
 AOI21x1_ASAP7_75t_R _23851_ (.A1(_15553_),
    .A2(_15554_),
    .B(_15051_),
    .Y(_15555_));
 AOI21x1_ASAP7_75t_R _23852_ (.A1(net5770),
    .A2(_15186_),
    .B(_15358_),
    .Y(_15556_));
 NAND2x1_ASAP7_75t_R _23853_ (.A(_15547_),
    .B(_15556_),
    .Y(_15557_));
 NAND2x1_ASAP7_75t_R _23854_ (.A(_15555_),
    .B(_15557_),
    .Y(_15558_));
 NAND2x1_ASAP7_75t_R _23855_ (.A(net5765),
    .B(net4901),
    .Y(_15559_));
 AOI21x1_ASAP7_75t_R _23856_ (.A1(_15283_),
    .A2(_15559_),
    .B(_14995_),
    .Y(_15560_));
 NAND2x1_ASAP7_75t_R _23857_ (.A(net6172),
    .B(net5765),
    .Y(_15561_));
 AOI21x1_ASAP7_75t_R _23858_ (.A1(_15561_),
    .A2(_15398_),
    .B(net5749),
    .Y(_15562_));
 OAI21x1_ASAP7_75t_R _23859_ (.A1(net5443),
    .A2(_15560_),
    .B(_15562_),
    .Y(_15563_));
 AOI21x1_ASAP7_75t_R _23860_ (.A1(_15558_),
    .A2(_15563_),
    .B(_15080_),
    .Y(_15564_));
 AO21x1_ASAP7_75t_R _23861_ (.A1(_14995_),
    .A2(net5776),
    .B(net5443),
    .Y(_15565_));
 AND2x2_ASAP7_75t_R _23862_ (.A(net4518),
    .B(net4751),
    .Y(_15566_));
 AOI21x1_ASAP7_75t_R _23863_ (.A1(_01201_),
    .A2(net5753),
    .B(net5151),
    .Y(_15567_));
 OAI21x1_ASAP7_75t_R _23864_ (.A1(net5143),
    .A2(_15326_),
    .B(net5773),
    .Y(_15568_));
 AOI21x1_ASAP7_75t_R _23865_ (.A1(_15567_),
    .A2(_15568_),
    .B(net5748),
    .Y(_15569_));
 OAI21x1_ASAP7_75t_R _23866_ (.A1(_15565_),
    .A2(_15566_),
    .B(_15569_),
    .Y(_15570_));
 NOR2x1_ASAP7_75t_R _23867_ (.A(net5158),
    .B(_14976_),
    .Y(_15571_));
 AOI21x1_ASAP7_75t_R _23868_ (.A1(net5755),
    .A2(_15571_),
    .B(net5150),
    .Y(_15572_));
 INVx1_ASAP7_75t_R _23869_ (.A(_15069_),
    .Y(_15573_));
 AOI21x1_ASAP7_75t_R _23870_ (.A1(_15573_),
    .A2(_15449_),
    .B(net5443),
    .Y(_15574_));
 OAI21x1_ASAP7_75t_R _23871_ (.A1(_15572_),
    .A2(_15574_),
    .B(net5748),
    .Y(_15575_));
 AOI21x1_ASAP7_75t_R _23872_ (.A1(_15570_),
    .A2(_15575_),
    .B(net6174),
    .Y(_15576_));
 OAI21x1_ASAP7_75t_R _23873_ (.A1(_15564_),
    .A2(_15576_),
    .B(net6173),
    .Y(_15577_));
 OAI21x1_ASAP7_75t_R _23874_ (.A1(_15536_),
    .A2(_15551_),
    .B(_15577_),
    .Y(_00086_));
 NAND2x1_ASAP7_75t_R _23875_ (.A(net5763),
    .B(_15155_),
    .Y(_15578_));
 AND2x2_ASAP7_75t_R _23876_ (.A(net5443),
    .B(net5156),
    .Y(_15579_));
 AND3x1_ASAP7_75t_R _23877_ (.A(_15578_),
    .B(_15006_),
    .C(_15579_),
    .Y(_15580_));
 AO21x1_ASAP7_75t_R _23878_ (.A1(net5766),
    .A2(_15107_),
    .B(net5443),
    .Y(_15581_));
 OAI21x1_ASAP7_75t_R _23879_ (.A1(_15581_),
    .A2(_15533_),
    .B(net6174),
    .Y(_15582_));
 OAI21x1_ASAP7_75t_R _23880_ (.A1(_15580_),
    .A2(_15582_),
    .B(net5749),
    .Y(_15583_));
 AO21x1_ASAP7_75t_R _23881_ (.A1(_15192_),
    .A2(net4674),
    .B(net5753),
    .Y(_15584_));
 AO21x1_ASAP7_75t_R _23882_ (.A1(_14998_),
    .A2(net6175),
    .B(_01206_),
    .Y(_15585_));
 AO21x1_ASAP7_75t_R _23883_ (.A1(_15584_),
    .A2(_15585_),
    .B(net5148),
    .Y(_15586_));
 AO21x1_ASAP7_75t_R _23884_ (.A1(_15272_),
    .A2(_15270_),
    .B(net5757),
    .Y(_15587_));
 AO21x1_ASAP7_75t_R _23885_ (.A1(_15099_),
    .A2(net4753),
    .B(net5765),
    .Y(_15588_));
 AO21x1_ASAP7_75t_R _23886_ (.A1(_15587_),
    .A2(_15588_),
    .B(net5443),
    .Y(_15589_));
 AOI21x1_ASAP7_75t_R _23887_ (.A1(_15586_),
    .A2(_15589_),
    .B(net6174),
    .Y(_15590_));
 NOR2x1_ASAP7_75t_R _23888_ (.A(_15583_),
    .B(_15590_),
    .Y(_15591_));
 INVx1_ASAP7_75t_R _23889_ (.A(_15376_),
    .Y(_15592_));
 AOI21x1_ASAP7_75t_R _23890_ (.A1(net6172),
    .A2(net5776),
    .B(net5443),
    .Y(_15593_));
 OAI21x1_ASAP7_75t_R _23891_ (.A1(net5763),
    .A2(_15084_),
    .B(_15593_),
    .Y(_15594_));
 OAI21x1_ASAP7_75t_R _23892_ (.A1(_15592_),
    .A2(_15594_),
    .B(net6174),
    .Y(_15595_));
 OA21x2_ASAP7_75t_R _23893_ (.A1(net5141),
    .A2(net4904),
    .B(net5776),
    .Y(_15596_));
 OAI21x1_ASAP7_75t_R _23894_ (.A1(net5776),
    .A2(_15391_),
    .B(net5443),
    .Y(_15597_));
 NOR2x1_ASAP7_75t_R _23895_ (.A(_15596_),
    .B(_15597_),
    .Y(_15598_));
 NOR2x1_ASAP7_75t_R _23896_ (.A(_15595_),
    .B(_15598_),
    .Y(_15599_));
 INVx1_ASAP7_75t_R _23897_ (.A(_15221_),
    .Y(_15600_));
 NAND2x1_ASAP7_75t_R _23898_ (.A(_15593_),
    .B(_15478_),
    .Y(_15601_));
 NOR2x1_ASAP7_75t_R _23899_ (.A(_15600_),
    .B(_15601_),
    .Y(_01549_));
 OA21x2_ASAP7_75t_R _23900_ (.A1(net5766),
    .A2(_15445_),
    .B(net5443),
    .Y(_01550_));
 AO21x1_ASAP7_75t_R _23901_ (.A1(_01550_),
    .A2(_15006_),
    .B(net6174),
    .Y(_01551_));
 OAI21x1_ASAP7_75t_R _23902_ (.A1(_01549_),
    .A2(_01551_),
    .B(net5751),
    .Y(_01552_));
 OAI21x1_ASAP7_75t_R _23903_ (.A1(_15599_),
    .A2(_01552_),
    .B(_15138_),
    .Y(_01553_));
 AOI211x1_ASAP7_75t_R _23904_ (.A1(net5762),
    .A2(_15208_),
    .B(net4748),
    .C(net5154),
    .Y(_01554_));
 AOI21x1_ASAP7_75t_R _23905_ (.A1(net5450),
    .A2(net5761),
    .B(net5443),
    .Y(_01555_));
 NAND2x1_ASAP7_75t_R _23906_ (.A(_15177_),
    .B(_01555_),
    .Y(_01556_));
 AOI21x1_ASAP7_75t_R _23907_ (.A1(net5450),
    .A2(net5438),
    .B(net4570),
    .Y(_01557_));
 OAI21x1_ASAP7_75t_R _23908_ (.A1(_01556_),
    .A2(_01557_),
    .B(net5749),
    .Y(_01558_));
 OAI21x1_ASAP7_75t_R _23909_ (.A1(_01554_),
    .A2(_01558_),
    .B(net5750),
    .Y(_01559_));
 NAND2x1_ASAP7_75t_R _23910_ (.A(net5142),
    .B(net5133),
    .Y(_01560_));
 AO21x1_ASAP7_75t_R _23911_ (.A1(net5767),
    .A2(net5778),
    .B(net5443),
    .Y(_01561_));
 AO21x1_ASAP7_75t_R _23912_ (.A1(net5761),
    .A2(_01560_),
    .B(_01561_),
    .Y(_01562_));
 INVx1_ASAP7_75t_R _23913_ (.A(net5140),
    .Y(_01563_));
 AOI21x1_ASAP7_75t_R _23914_ (.A1(_15272_),
    .A2(_01563_),
    .B(net5757),
    .Y(_01564_));
 OAI21x1_ASAP7_75t_R _23915_ (.A1(_15284_),
    .A2(_01564_),
    .B(net5443),
    .Y(_01565_));
 AOI21x1_ASAP7_75t_R _23916_ (.A1(_01562_),
    .A2(_01565_),
    .B(net5749),
    .Y(_01566_));
 OAI21x1_ASAP7_75t_R _23917_ (.A1(_01559_),
    .A2(_01566_),
    .B(net6173),
    .Y(_01567_));
 AO21x1_ASAP7_75t_R _23918_ (.A1(net4901),
    .A2(net5776),
    .B(net5154),
    .Y(_01568_));
 OAI21x1_ASAP7_75t_R _23919_ (.A1(_15450_),
    .A2(_01568_),
    .B(net5751),
    .Y(_01569_));
 OA21x2_ASAP7_75t_R _23920_ (.A1(net5141),
    .A2(net4904),
    .B(net5759),
    .Y(_01570_));
 OAI21x1_ASAP7_75t_R _23921_ (.A1(net5146),
    .A2(_15510_),
    .B(net5153),
    .Y(_01571_));
 NOR2x1_ASAP7_75t_R _23922_ (.A(_01570_),
    .B(_01571_),
    .Y(_01572_));
 OAI21x1_ASAP7_75t_R _23923_ (.A1(_01569_),
    .A2(_01572_),
    .B(net6174),
    .Y(_01573_));
 AND2x2_ASAP7_75t_R _23924_ (.A(_15261_),
    .B(net5759),
    .Y(_01574_));
 NOR2x1_ASAP7_75t_R _23925_ (.A(net5001),
    .B(_15510_),
    .Y(_01575_));
 OAI21x1_ASAP7_75t_R _23926_ (.A1(_01574_),
    .A2(_01575_),
    .B(net5153),
    .Y(_01576_));
 NOR2x1_ASAP7_75t_R _23927_ (.A(net5137),
    .B(net4898),
    .Y(_01577_));
 OAI21x1_ASAP7_75t_R _23928_ (.A1(_15522_),
    .A2(_01577_),
    .B(net5443),
    .Y(_01578_));
 AOI21x1_ASAP7_75t_R _23929_ (.A1(_01578_),
    .A2(_01576_),
    .B(net5751),
    .Y(_01579_));
 NOR2x1_ASAP7_75t_R _23930_ (.A(_01573_),
    .B(_01579_),
    .Y(_01580_));
 OAI22x1_ASAP7_75t_R _23931_ (.A1(_15591_),
    .A2(_01553_),
    .B1(_01580_),
    .B2(_01567_),
    .Y(_00087_));
 NOR2x1_ASAP7_75t_R _23932_ (.A(net6661),
    .B(_00465_),
    .Y(_01581_));
 INVx1_ASAP7_75t_R _23933_ (.A(net6627),
    .Y(_01582_));
 XOR2x2_ASAP7_75t_R _23934_ (.A(_01582_),
    .B(_12812_),
    .Y(_01583_));
 XNOR2x2_ASAP7_75t_R _23935_ (.A(net6577),
    .B(_00670_),
    .Y(_01584_));
 XOR2x2_ASAP7_75t_R _23936_ (.A(net6547),
    .B(_00664_),
    .Y(_01585_));
 XOR2x2_ASAP7_75t_R _23937_ (.A(_01584_),
    .B(_01585_),
    .Y(_01586_));
 NAND2x1p5_ASAP7_75t_R _23938_ (.A(_01586_),
    .B(_01583_),
    .Y(_01587_));
 XOR2x2_ASAP7_75t_R _23939_ (.A(net6627),
    .B(_12812_),
    .Y(_01588_));
 XOR2x2_ASAP7_75t_R _23940_ (.A(_00670_),
    .B(net6577),
    .Y(_01589_));
 XOR2x2_ASAP7_75t_R _23941_ (.A(_01589_),
    .B(_01585_),
    .Y(_01590_));
 NAND2x1p5_ASAP7_75t_R _23942_ (.A(_01590_),
    .B(_01588_),
    .Y(_01591_));
 AOI21x1_ASAP7_75t_R _23943_ (.A1(_01591_),
    .A2(_01587_),
    .B(net6457),
    .Y(_01592_));
 OAI21x1_ASAP7_75t_R _23944_ (.A1(net6407),
    .A2(net6354),
    .B(net6474),
    .Y(_01593_));
 AND2x2_ASAP7_75t_R _23945_ (.A(net6460),
    .B(_00465_),
    .Y(_01594_));
 NAND2x1p5_ASAP7_75t_R _23946_ (.A(_01588_),
    .B(_01586_),
    .Y(_01595_));
 NAND2x1p5_ASAP7_75t_R _23947_ (.A(_01590_),
    .B(_01583_),
    .Y(_01596_));
 AOI21x1_ASAP7_75t_R _23948_ (.A1(_01596_),
    .A2(_01595_),
    .B(net6457),
    .Y(_01597_));
 OAI21x1_ASAP7_75t_R _23949_ (.A1(_01594_),
    .A2(net6353),
    .B(_08063_),
    .Y(_01598_));
 NAND2x1_ASAP7_75t_R _23950_ (.A(_01593_),
    .B(_01598_),
    .Y(_01599_));
 XOR2x2_ASAP7_75t_R _23952_ (.A(net6628),
    .B(net6601),
    .Y(_01600_));
 NAND2x1_ASAP7_75t_R _23953_ (.A(_12833_),
    .B(_01600_),
    .Y(_01601_));
 XNOR2x2_ASAP7_75t_R _23954_ (.A(net6628),
    .B(net6601),
    .Y(_01602_));
 NAND2x1_ASAP7_75t_R _23955_ (.A(net6548),
    .B(_01602_),
    .Y(_01603_));
 AOI21x1_ASAP7_75t_R _23956_ (.A1(_01601_),
    .A2(_01603_),
    .B(net6406),
    .Y(_01604_));
 XOR2x2_ASAP7_75t_R _23957_ (.A(net6601),
    .B(net6548),
    .Y(_01605_));
 NAND2x1_ASAP7_75t_R _23958_ (.A(net6628),
    .B(_01605_),
    .Y(_01606_));
 INVx1_ASAP7_75t_R _23959_ (.A(net6628),
    .Y(_01607_));
 XNOR2x2_ASAP7_75t_R _23960_ (.A(net6601),
    .B(net6548),
    .Y(_01608_));
 NAND2x1_ASAP7_75t_R _23961_ (.A(_01607_),
    .B(_01608_),
    .Y(_01609_));
 AOI21x1_ASAP7_75t_R _23962_ (.A1(_01606_),
    .A2(_01609_),
    .B(net6404),
    .Y(_01610_));
 NOR2x1_ASAP7_75t_R _23963_ (.A(_01604_),
    .B(_01610_),
    .Y(_01611_));
 AND2x2_ASAP7_75t_R _23964_ (.A(net6460),
    .B(_00466_),
    .Y(_01612_));
 AOI21x1_ASAP7_75t_R _23965_ (.A1(net6663),
    .A2(_01611_),
    .B(_01612_),
    .Y(_01613_));
 XOR2x2_ASAP7_75t_R _23966_ (.A(net6171),
    .B(_08046_),
    .Y(_01215_));
 NOR2x1_ASAP7_75t_R _23967_ (.A(net6662),
    .B(_00467_),
    .Y(_01614_));
 INVx1_ASAP7_75t_R _23968_ (.A(_01614_),
    .Y(_01615_));
 INVx1_ASAP7_75t_R _23969_ (.A(net6625),
    .Y(_01616_));
 NOR2x1_ASAP7_75t_R _23970_ (.A(_01616_),
    .B(_12859_),
    .Y(_01617_));
 NOR2x1_ASAP7_75t_R _23971_ (.A(net6625),
    .B(_12855_),
    .Y(_01618_));
 OAI21x1_ASAP7_75t_R _23972_ (.A1(_01617_),
    .A2(_01618_),
    .B(net6426),
    .Y(_01619_));
 INVx1_ASAP7_75t_R _23973_ (.A(_01619_),
    .Y(_01620_));
 NOR3x1_ASAP7_75t_R _23974_ (.A(_01618_),
    .B(_01617_),
    .C(net6426),
    .Y(_01621_));
 OAI21x1_ASAP7_75t_R _23975_ (.A1(_01620_),
    .A2(_01621_),
    .B(net6662),
    .Y(_01622_));
 INVx1_ASAP7_75t_R _23976_ (.A(_00943_),
    .Y(_01623_));
 AOI21x1_ASAP7_75t_R _23977_ (.A1(_01615_),
    .A2(_01622_),
    .B(_01623_),
    .Y(_01624_));
 NAND2x1_ASAP7_75t_R _23978_ (.A(_00467_),
    .B(net6460),
    .Y(_01625_));
 NAND2x1_ASAP7_75t_R _23979_ (.A(_01616_),
    .B(_12859_),
    .Y(_01626_));
 INVx1_ASAP7_75t_R _23980_ (.A(net6426),
    .Y(_01627_));
 NOR2x1_ASAP7_75t_R _23981_ (.A(net6574),
    .B(net6544),
    .Y(_01628_));
 AND2x2_ASAP7_75t_R _23982_ (.A(net6574),
    .B(net6544),
    .Y(_01629_));
 OAI21x1_ASAP7_75t_R _23983_ (.A1(_01628_),
    .A2(_01629_),
    .B(net6625),
    .Y(_01630_));
 NAND3x1_ASAP7_75t_R _23984_ (.A(_01626_),
    .B(_01627_),
    .C(_01630_),
    .Y(_01631_));
 NAND3x1_ASAP7_75t_R _23985_ (.A(_01631_),
    .B(net6662),
    .C(_01619_),
    .Y(_01632_));
 AOI21x1_ASAP7_75t_R _23986_ (.A1(_01625_),
    .A2(_01632_),
    .B(_00943_),
    .Y(_01633_));
 NOR2x1_ASAP7_75t_R _23987_ (.A(_01624_),
    .B(_01633_),
    .Y(_01634_));
 XOR2x2_ASAP7_75t_R _23990_ (.A(_01613_),
    .B(net6475),
    .Y(_01636_));
 AOI21x1_ASAP7_75t_R _23992_ (.A1(_01615_),
    .A2(_01622_),
    .B(_00943_),
    .Y(_01637_));
 AOI21x1_ASAP7_75t_R _23993_ (.A1(_01625_),
    .A2(_01632_),
    .B(_01623_),
    .Y(_01638_));
 NOR2x1_ASAP7_75t_R _23994_ (.A(_01637_),
    .B(_01638_),
    .Y(_01639_));
 NOR2x1_ASAP7_75t_R _23997_ (.A(net6662),
    .B(_00543_),
    .Y(_01641_));
 XNOR2x2_ASAP7_75t_R _23998_ (.A(_00603_),
    .B(_12908_),
    .Y(_01642_));
 XOR2x2_ASAP7_75t_R _23999_ (.A(net6573),
    .B(net6570),
    .Y(_01643_));
 XOR2x2_ASAP7_75t_R _24000_ (.A(_12907_),
    .B(_01643_),
    .Y(_01644_));
 NAND2x1_ASAP7_75t_R _24001_ (.A(_01642_),
    .B(_01644_),
    .Y(_01645_));
 OR2x2_ASAP7_75t_R _24002_ (.A(_01642_),
    .B(_01644_),
    .Y(_01646_));
 AOI21x1_ASAP7_75t_R _24003_ (.A1(_01645_),
    .A2(_01646_),
    .B(net6458),
    .Y(_01647_));
 OAI21x1_ASAP7_75t_R _24004_ (.A1(_01641_),
    .A2(_01647_),
    .B(_00946_),
    .Y(_01648_));
 AND2x2_ASAP7_75t_R _24005_ (.A(net6458),
    .B(_00543_),
    .Y(_01649_));
 XNOR2x2_ASAP7_75t_R _24006_ (.A(_01642_),
    .B(_01644_),
    .Y(_01650_));
 NOR2x1_ASAP7_75t_R _24007_ (.A(net6458),
    .B(_01650_),
    .Y(_01651_));
 OAI21x1_ASAP7_75t_R _24008_ (.A1(_01649_),
    .A2(_01651_),
    .B(_08069_),
    .Y(_01652_));
 NAND2x1_ASAP7_75t_R _24009_ (.A(_01648_),
    .B(_01652_),
    .Y(_01653_));
 INVx2_ASAP7_75t_R _24010_ (.A(_01653_),
    .Y(_01654_));
 XOR2x2_ASAP7_75t_R _24014_ (.A(_12885_),
    .B(_00602_),
    .Y(_01658_));
 XOR2x2_ASAP7_75t_R _24015_ (.A(net6574),
    .B(net6570),
    .Y(_01659_));
 XOR2x2_ASAP7_75t_R _24016_ (.A(_12889_),
    .B(_01659_),
    .Y(_01660_));
 NOR2x1_ASAP7_75t_R _24017_ (.A(_01658_),
    .B(_01660_),
    .Y(_01661_));
 XNOR2x2_ASAP7_75t_R _24018_ (.A(_00602_),
    .B(_12885_),
    .Y(_01662_));
 XOR2x2_ASAP7_75t_R _24019_ (.A(_12884_),
    .B(_01659_),
    .Y(_01663_));
 NOR2x1_ASAP7_75t_R _24020_ (.A(_01662_),
    .B(_01663_),
    .Y(_01664_));
 OAI21x1_ASAP7_75t_R _24021_ (.A1(_01661_),
    .A2(_01664_),
    .B(net6662),
    .Y(_01665_));
 NOR2x1_ASAP7_75t_R _24022_ (.A(net6661),
    .B(_00544_),
    .Y(_01666_));
 INVx1_ASAP7_75t_R _24023_ (.A(_01666_),
    .Y(_01667_));
 NAND3x1_ASAP7_75t_R _24024_ (.A(_01665_),
    .B(_00944_),
    .C(_01667_),
    .Y(_01668_));
 AO21x1_ASAP7_75t_R _24025_ (.A1(_01665_),
    .A2(_01667_),
    .B(_00944_),
    .Y(_01669_));
 NAND2x2_ASAP7_75t_R _24026_ (.A(_01668_),
    .B(_01669_),
    .Y(_01670_));
 OA21x2_ASAP7_75t_R _24027_ (.A1(net5280),
    .A2(net5431),
    .B(net5728),
    .Y(_01671_));
 OAI21x1_ASAP7_75t_R _24028_ (.A1(_01592_),
    .A2(_01581_),
    .B(_08063_),
    .Y(_01672_));
 OAI21x1_ASAP7_75t_R _24029_ (.A1(_01597_),
    .A2(_01594_),
    .B(net6474),
    .Y(_01673_));
 NAND2x1p5_ASAP7_75t_R _24030_ (.A(_01673_),
    .B(_01672_),
    .Y(_01674_));
 NOR2x1_ASAP7_75t_R _24031_ (.A(net5744),
    .B(net5724),
    .Y(_01675_));
 NAND2x1_ASAP7_75t_R _24032_ (.A(net5432),
    .B(_01675_),
    .Y(_01676_));
 INVx1_ASAP7_75t_R _24034_ (.A(_01212_),
    .Y(_01678_));
 NAND2x1_ASAP7_75t_R _24035_ (.A(_01678_),
    .B(net5433),
    .Y(_01679_));
 NOR2x1_ASAP7_75t_R _24036_ (.A(net5734),
    .B(_01679_),
    .Y(_01680_));
 AO21x1_ASAP7_75t_R _24037_ (.A1(_01671_),
    .A2(_01676_),
    .B(_01680_),
    .Y(_01681_));
 NAND3x1_ASAP7_75t_R _24038_ (.A(_01665_),
    .B(_08038_),
    .C(_01667_),
    .Y(_01682_));
 AO21x1_ASAP7_75t_R _24039_ (.A1(_01665_),
    .A2(_01667_),
    .B(_08038_),
    .Y(_01683_));
 NAND2x1_ASAP7_75t_R _24040_ (.A(_01682_),
    .B(_01683_),
    .Y(_01684_));
 OA21x2_ASAP7_75t_R _24042_ (.A1(_01679_),
    .A2(net5717),
    .B(net5429),
    .Y(_01686_));
 INVx1_ASAP7_75t_R _24043_ (.A(_01217_),
    .Y(_01687_));
 OAI21x1_ASAP7_75t_R _24044_ (.A1(net5130),
    .A2(net5430),
    .B(net5718),
    .Y(_01688_));
 INVx1_ASAP7_75t_R _24045_ (.A(_01688_),
    .Y(_01689_));
 NAND2x1_ASAP7_75t_R _24046_ (.A(_01689_),
    .B(_01676_),
    .Y(_01690_));
 XNOR2x2_ASAP7_75t_R _24047_ (.A(_00604_),
    .B(_00635_),
    .Y(_01691_));
 XOR2x2_ASAP7_75t_R _24048_ (.A(net6572),
    .B(_00668_),
    .Y(_01692_));
 XOR2x2_ASAP7_75t_R _24049_ (.A(_01692_),
    .B(_00700_),
    .Y(_01693_));
 INVx1_ASAP7_75t_R _24050_ (.A(_01693_),
    .Y(_01694_));
 NAND2x1_ASAP7_75t_R _24051_ (.A(_01691_),
    .B(_01694_),
    .Y(_01695_));
 INVx1_ASAP7_75t_R _24052_ (.A(_01691_),
    .Y(_01696_));
 NAND2x1_ASAP7_75t_R _24053_ (.A(_01696_),
    .B(_01693_),
    .Y(_01697_));
 AO21x1_ASAP7_75t_R _24054_ (.A1(_01695_),
    .A2(_01697_),
    .B(net6458),
    .Y(_01698_));
 OR2x2_ASAP7_75t_R _24055_ (.A(net6664),
    .B(_00542_),
    .Y(_01699_));
 AND2x2_ASAP7_75t_R _24056_ (.A(_01698_),
    .B(_01699_),
    .Y(_01700_));
 INVx1_ASAP7_75t_R _24057_ (.A(_00947_),
    .Y(_01701_));
 XOR2x2_ASAP7_75t_R _24058_ (.A(_01700_),
    .B(_01701_),
    .Y(_01702_));
 AOI21x1_ASAP7_75t_R _24059_ (.A1(_01686_),
    .A2(_01690_),
    .B(net5423),
    .Y(_01703_));
 OAI21x1_ASAP7_75t_R _24060_ (.A1(net5429),
    .A2(_01681_),
    .B(_01703_),
    .Y(_01704_));
 INVx1_ASAP7_75t_R _24061_ (.A(_01214_),
    .Y(_01705_));
 OAI21x1_ASAP7_75t_R _24062_ (.A1(net5741),
    .A2(net6169),
    .B(_01705_),
    .Y(_01706_));
 INVx1_ASAP7_75t_R _24063_ (.A(_01706_),
    .Y(_01707_));
 AOI21x1_ASAP7_75t_R _24064_ (.A1(net5742),
    .A2(net5746),
    .B(net5435),
    .Y(_01708_));
 OAI21x1_ASAP7_75t_R _24066_ (.A1(_01707_),
    .A2(_01708_),
    .B(net5730),
    .Y(_01710_));
 NAND2x1_ASAP7_75t_R _24067_ (.A(_01210_),
    .B(net5433),
    .Y(_01711_));
 NAND2x1_ASAP7_75t_R _24068_ (.A(net5744),
    .B(net5435),
    .Y(_01712_));
 AOI21x1_ASAP7_75t_R _24070_ (.A1(_01711_),
    .A2(_01712_),
    .B(net5728),
    .Y(_01714_));
 OAI21x1_ASAP7_75t_R _24071_ (.A1(net5741),
    .A2(net6169),
    .B(_01678_),
    .Y(_01715_));
 INVx1_ASAP7_75t_R _24072_ (.A(_01715_),
    .Y(_01716_));
 AO21x1_ASAP7_75t_R _24074_ (.A1(_01716_),
    .A2(net5733),
    .B(net5740),
    .Y(_01718_));
 NOR2x1_ASAP7_75t_R _24075_ (.A(_01714_),
    .B(_01718_),
    .Y(_01719_));
 NAND2x1_ASAP7_75t_R _24076_ (.A(_01710_),
    .B(_01719_),
    .Y(_01720_));
 INVx1_ASAP7_75t_R _24077_ (.A(_01211_),
    .Y(_01721_));
 OAI21x1_ASAP7_75t_R _24078_ (.A1(net5741),
    .A2(net6169),
    .B(_01721_),
    .Y(_01722_));
 INVx2_ASAP7_75t_R _24079_ (.A(_01722_),
    .Y(_01723_));
 AO21x1_ASAP7_75t_R _24080_ (.A1(_01723_),
    .A2(net5728),
    .B(net5427),
    .Y(_01724_));
 NOR2x1_ASAP7_75t_R _24081_ (.A(_01224_),
    .B(net5728),
    .Y(_01725_));
 OA21x2_ASAP7_75t_R _24082_ (.A1(_01724_),
    .A2(_01725_),
    .B(net5424),
    .Y(_01726_));
 XOR2x2_ASAP7_75t_R _24083_ (.A(_00669_),
    .B(_00701_),
    .Y(_01727_));
 XOR2x2_ASAP7_75t_R _24084_ (.A(_12959_),
    .B(_00605_),
    .Y(_01728_));
 XNOR2x2_ASAP7_75t_R _24085_ (.A(_01727_),
    .B(_01728_),
    .Y(_01729_));
 NOR2x1_ASAP7_75t_R _24086_ (.A(net6661),
    .B(_00541_),
    .Y(_01730_));
 AO21x1_ASAP7_75t_R _24087_ (.A1(_01729_),
    .A2(net6662),
    .B(_01730_),
    .Y(_01731_));
 XOR2x2_ASAP7_75t_R _24088_ (.A(_01731_),
    .B(_00948_),
    .Y(_01732_));
 INVx1_ASAP7_75t_R _24089_ (.A(_01732_),
    .Y(_01733_));
 AOI21x1_ASAP7_75t_R _24090_ (.A1(_01720_),
    .A2(_01726_),
    .B(net5715),
    .Y(_01734_));
 NAND2x1_ASAP7_75t_R _24091_ (.A(_01734_),
    .B(_01704_),
    .Y(_01735_));
 AOI21x1_ASAP7_75t_R _24092_ (.A1(net5281),
    .A2(net5432),
    .B(net5734),
    .Y(_01736_));
 INVx1_ASAP7_75t_R _24093_ (.A(_01736_),
    .Y(_01737_));
 NAND2x1_ASAP7_75t_R _24095_ (.A(_01210_),
    .B(net5436),
    .Y(_01739_));
 AO21x1_ASAP7_75t_R _24097_ (.A1(_01739_),
    .A2(_01679_),
    .B(net5717),
    .Y(_01741_));
 AOI21x1_ASAP7_75t_R _24099_ (.A1(_01737_),
    .A2(_01741_),
    .B(net5429),
    .Y(_01743_));
 OAI21x1_ASAP7_75t_R _24100_ (.A1(net5741),
    .A2(net6169),
    .B(net5254),
    .Y(_01744_));
 OAI21x1_ASAP7_75t_R _24101_ (.A1(net5746),
    .A2(net5435),
    .B(_01744_),
    .Y(_01745_));
 NAND2x1_ASAP7_75t_R _24102_ (.A(net5730),
    .B(_01745_),
    .Y(_01746_));
 NAND2x1_ASAP7_75t_R _24103_ (.A(net5744),
    .B(net5433),
    .Y(_01747_));
 NAND2x1_ASAP7_75t_R _24104_ (.A(net5280),
    .B(net5435),
    .Y(_01748_));
 AO21x1_ASAP7_75t_R _24106_ (.A1(net5126),
    .A2(_01748_),
    .B(net5734),
    .Y(_01750_));
 AOI21x1_ASAP7_75t_R _24108_ (.A1(net4567),
    .A2(_01750_),
    .B(net5739),
    .Y(_01752_));
 XOR2x2_ASAP7_75t_R _24109_ (.A(_01700_),
    .B(_00947_),
    .Y(_01753_));
 OAI21x1_ASAP7_75t_R _24111_ (.A1(_01743_),
    .A2(_01752_),
    .B(net5422),
    .Y(_01755_));
 NOR2x1_ASAP7_75t_R _24112_ (.A(net5744),
    .B(net5433),
    .Y(_01756_));
 NOR2x1_ASAP7_75t_R _24113_ (.A(net5734),
    .B(_01756_),
    .Y(_01757_));
 NOR2x1_ASAP7_75t_R _24114_ (.A(net5742),
    .B(net5724),
    .Y(_01758_));
 NAND2x1_ASAP7_75t_R _24115_ (.A(net5432),
    .B(_01758_),
    .Y(_01759_));
 OAI21x1_ASAP7_75t_R _24117_ (.A1(net5723),
    .A2(net4895),
    .B(net5428),
    .Y(_01761_));
 AO21x1_ASAP7_75t_R _24118_ (.A1(_01757_),
    .A2(net5124),
    .B(_01761_),
    .Y(_01762_));
 OA21x2_ASAP7_75t_R _24119_ (.A1(net5723),
    .A2(_01706_),
    .B(net5740),
    .Y(_01763_));
 OAI21x1_ASAP7_75t_R _24120_ (.A1(net5743),
    .A2(net6170),
    .B(_01687_),
    .Y(_01764_));
 NOR2x1_ASAP7_75t_R _24121_ (.A(_01764_),
    .B(net5723),
    .Y(_01765_));
 OA21x2_ASAP7_75t_R _24122_ (.A1(net6170),
    .A2(net5743),
    .B(net5254),
    .Y(_01766_));
 NOR2x1_ASAP7_75t_R _24123_ (.A(net5734),
    .B(_01766_),
    .Y(_01767_));
 NOR2x1_ASAP7_75t_R _24124_ (.A(_01765_),
    .B(_01767_),
    .Y(_01768_));
 AOI21x1_ASAP7_75t_R _24126_ (.A1(_01763_),
    .A2(_01768_),
    .B(net5422),
    .Y(_01770_));
 AOI21x1_ASAP7_75t_R _24127_ (.A1(_01762_),
    .A2(_01770_),
    .B(net6168),
    .Y(_01771_));
 XOR2x2_ASAP7_75t_R _24128_ (.A(net6542),
    .B(_00669_),
    .Y(_01772_));
 INVx1_ASAP7_75t_R _24129_ (.A(net6571),
    .Y(_01773_));
 XOR2x2_ASAP7_75t_R _24130_ (.A(_01772_),
    .B(net6403),
    .Y(_01774_));
 XOR2x2_ASAP7_75t_R _24131_ (.A(net6624),
    .B(_00637_),
    .Y(_01775_));
 XOR2x2_ASAP7_75t_R _24132_ (.A(_01774_),
    .B(_01775_),
    .Y(_01776_));
 NOR2x1_ASAP7_75t_R _24133_ (.A(net6661),
    .B(_00540_),
    .Y(_01777_));
 AO21x1_ASAP7_75t_R _24134_ (.A1(_01776_),
    .A2(net6661),
    .B(_01777_),
    .Y(_01778_));
 XOR2x2_ASAP7_75t_R _24135_ (.A(_01778_),
    .B(_00949_),
    .Y(_01779_));
 AOI21x1_ASAP7_75t_R _24137_ (.A1(_01755_),
    .A2(_01771_),
    .B(net6167),
    .Y(_01781_));
 NAND2x1_ASAP7_75t_R _24138_ (.A(_01781_),
    .B(_01735_),
    .Y(_01782_));
 NAND2x1_ASAP7_75t_R _24140_ (.A(net5742),
    .B(net5724),
    .Y(_01783_));
 AO21x1_ASAP7_75t_R _24141_ (.A1(_01783_),
    .A2(net5126),
    .B(net5725),
    .Y(_01784_));
 NAND2x1_ASAP7_75t_R _24142_ (.A(net5742),
    .B(net5747),
    .Y(_01785_));
 AO21x1_ASAP7_75t_R _24143_ (.A1(net5418),
    .A2(_01712_),
    .B(net5718),
    .Y(_01786_));
 AND3x1_ASAP7_75t_R _24144_ (.A(_01784_),
    .B(_01786_),
    .C(net5735),
    .Y(_01787_));
 NAND2x1_ASAP7_75t_R _24146_ (.A(net5280),
    .B(net5431),
    .Y(_01789_));
 NAND2x1_ASAP7_75t_R _24147_ (.A(_01789_),
    .B(_01739_),
    .Y(_01790_));
 AOI21x1_ASAP7_75t_R _24149_ (.A1(net5719),
    .A2(_01790_),
    .B(net5740),
    .Y(_01792_));
 OAI21x1_ASAP7_75t_R _24150_ (.A1(net5742),
    .A2(net5724),
    .B(net5434),
    .Y(_01793_));
 OAI21x1_ASAP7_75t_R _24151_ (.A1(net5743),
    .A2(net6170),
    .B(_01721_),
    .Y(_01794_));
 AO21x1_ASAP7_75t_R _24154_ (.A1(_01793_),
    .A2(net4744),
    .B(net5719),
    .Y(_01797_));
 AO21x1_ASAP7_75t_R _24155_ (.A1(_01792_),
    .A2(_01797_),
    .B(net5715),
    .Y(_01798_));
 NAND2x1_ASAP7_75t_R _24158_ (.A(net5277),
    .B(net5436),
    .Y(_01801_));
 NAND2x1_ASAP7_75t_R _24159_ (.A(net5721),
    .B(_01801_),
    .Y(_01802_));
 AO21x1_ASAP7_75t_R _24161_ (.A1(net5724),
    .A2(net5434),
    .B(net5744),
    .Y(_01804_));
 AOI21x1_ASAP7_75t_R _24163_ (.A1(net5725),
    .A2(_01804_),
    .B(net5429),
    .Y(_01806_));
 OAI21x1_ASAP7_75t_R _24164_ (.A1(net4998),
    .A2(_01802_),
    .B(_01806_),
    .Y(_01807_));
 NAND2x1_ASAP7_75t_R _24165_ (.A(net5436),
    .B(net5426),
    .Y(_01808_));
 NAND2x1_ASAP7_75t_R _24166_ (.A(_01736_),
    .B(_01808_),
    .Y(_01809_));
 NOR2x1_ASAP7_75t_R _24168_ (.A(net5719),
    .B(_01756_),
    .Y(_01811_));
 NOR2x1_ASAP7_75t_R _24169_ (.A(net5736),
    .B(_01811_),
    .Y(_01812_));
 AOI21x1_ASAP7_75t_R _24170_ (.A1(_01809_),
    .A2(_01812_),
    .B(net6168),
    .Y(_01813_));
 AOI21x1_ASAP7_75t_R _24172_ (.A1(_01807_),
    .A2(_01813_),
    .B(net5423),
    .Y(_01815_));
 OAI21x1_ASAP7_75t_R _24173_ (.A1(_01787_),
    .A2(_01798_),
    .B(_01815_),
    .Y(_01816_));
 INVx1_ASAP7_75t_R _24174_ (.A(_01794_),
    .Y(_01817_));
 INVx1_ASAP7_75t_R _24175_ (.A(_01210_),
    .Y(_01818_));
 NOR2x1_ASAP7_75t_R _24176_ (.A(_01818_),
    .B(net5433),
    .Y(_01819_));
 OAI21x1_ASAP7_75t_R _24177_ (.A1(_01817_),
    .A2(_01819_),
    .B(net5723),
    .Y(_01820_));
 OA21x2_ASAP7_75t_R _24178_ (.A1(net6170),
    .A2(net5743),
    .B(_01210_),
    .Y(_01821_));
 AOI21x1_ASAP7_75t_R _24179_ (.A1(net5728),
    .A2(_01821_),
    .B(net5740),
    .Y(_01822_));
 INVx1_ASAP7_75t_R _24180_ (.A(_01216_),
    .Y(_01823_));
 NOR2x1_ASAP7_75t_R _24181_ (.A(_01823_),
    .B(net5431),
    .Y(_01824_));
 NAND2x1_ASAP7_75t_R _24182_ (.A(net5728),
    .B(net4890),
    .Y(_01825_));
 NAND3x1_ASAP7_75t_R _24183_ (.A(_01820_),
    .B(_01822_),
    .C(_01825_),
    .Y(_01826_));
 NOR2x1_ASAP7_75t_R _24185_ (.A(_01744_),
    .B(net5733),
    .Y(_01828_));
 NOR2x1_ASAP7_75t_R _24186_ (.A(net5428),
    .B(_01828_),
    .Y(_01829_));
 NAND2x1_ASAP7_75t_R _24187_ (.A(net5435),
    .B(net5747),
    .Y(_01830_));
 AO21x1_ASAP7_75t_R _24188_ (.A1(_01830_),
    .A2(net4743),
    .B(net5719),
    .Y(_01831_));
 AOI21x1_ASAP7_75t_R _24189_ (.A1(_01829_),
    .A2(_01831_),
    .B(_01733_),
    .Y(_01832_));
 AOI21x1_ASAP7_75t_R _24190_ (.A1(_01826_),
    .A2(_01832_),
    .B(net5421),
    .Y(_01833_));
 NAND2x1_ASAP7_75t_R _24191_ (.A(net5437),
    .B(net5724),
    .Y(_01834_));
 AO21x1_ASAP7_75t_R _24192_ (.A1(net5123),
    .A2(_01679_),
    .B(net5717),
    .Y(_01835_));
 AOI21x1_ASAP7_75t_R _24193_ (.A1(net5124),
    .A2(_01757_),
    .B(net5739),
    .Y(_01836_));
 NAND2x1_ASAP7_75t_R _24194_ (.A(_01835_),
    .B(_01836_),
    .Y(_01837_));
 OAI21x1_ASAP7_75t_R _24195_ (.A1(net5744),
    .A2(net5724),
    .B(net5434),
    .Y(_01838_));
 NAND2x1_ASAP7_75t_R _24196_ (.A(net5433),
    .B(net5745),
    .Y(_01839_));
 AO21x1_ASAP7_75t_R _24197_ (.A1(_01838_),
    .A2(_01839_),
    .B(net5719),
    .Y(_01840_));
 NAND2x1_ASAP7_75t_R _24198_ (.A(net5277),
    .B(net5430),
    .Y(_01841_));
 AOI21x1_ASAP7_75t_R _24199_ (.A1(_01841_),
    .A2(_01757_),
    .B(net5429),
    .Y(_01842_));
 AOI21x1_ASAP7_75t_R _24200_ (.A1(_01840_),
    .A2(_01842_),
    .B(net6168),
    .Y(_01843_));
 NAND2x1_ASAP7_75t_R _24201_ (.A(_01837_),
    .B(_01843_),
    .Y(_01844_));
 INVx1_ASAP7_75t_R _24202_ (.A(_01779_),
    .Y(_01845_));
 AOI21x1_ASAP7_75t_R _24203_ (.A1(_01833_),
    .A2(_01844_),
    .B(_01845_),
    .Y(_01846_));
 NAND2x1_ASAP7_75t_R _24204_ (.A(_01816_),
    .B(_01846_),
    .Y(_01847_));
 NAND2x1_ASAP7_75t_R _24205_ (.A(_01847_),
    .B(_01782_),
    .Y(_00088_));
 AOI21x1_ASAP7_75t_R _24206_ (.A1(net5744),
    .A2(net5747),
    .B(net5431),
    .Y(_01848_));
 OAI21x1_ASAP7_75t_R _24207_ (.A1(net4996),
    .A2(_01848_),
    .B(net5722),
    .Y(_01849_));
 OAI21x1_ASAP7_75t_R _24208_ (.A1(net5277),
    .A2(net5435),
    .B(net4894),
    .Y(_01850_));
 AOI21x1_ASAP7_75t_R _24209_ (.A1(net5733),
    .A2(_01850_),
    .B(net5427),
    .Y(_01851_));
 NAND2x1_ASAP7_75t_R _24210_ (.A(_01849_),
    .B(_01851_),
    .Y(_01852_));
 NOR2x1_ASAP7_75t_R _24211_ (.A(net5742),
    .B(net5431),
    .Y(_01853_));
 AOI21x1_ASAP7_75t_R _24212_ (.A1(net5744),
    .A2(net5746),
    .B(net5435),
    .Y(_01854_));
 OAI21x1_ASAP7_75t_R _24214_ (.A1(net5121),
    .A2(_01854_),
    .B(net5732),
    .Y(_01856_));
 OA21x2_ASAP7_75t_R _24215_ (.A1(net4996),
    .A2(net5732),
    .B(net5427),
    .Y(_01857_));
 AOI21x1_ASAP7_75t_R _24216_ (.A1(_01856_),
    .A2(_01857_),
    .B(net5421),
    .Y(_01858_));
 NAND2x1_ASAP7_75t_R _24217_ (.A(_01852_),
    .B(_01858_),
    .Y(_01859_));
 OAI21x1_ASAP7_75t_R _24219_ (.A1(_01723_),
    .A2(_01821_),
    .B(net5719),
    .Y(_01861_));
 NOR2x1_ASAP7_75t_R _24220_ (.A(net5282),
    .B(net5435),
    .Y(_01862_));
 OAI21x1_ASAP7_75t_R _24222_ (.A1(_01862_),
    .A2(net5121),
    .B(net5728),
    .Y(_01864_));
 AOI21x1_ASAP7_75t_R _24223_ (.A1(_01861_),
    .A2(_01864_),
    .B(net5427),
    .Y(_01865_));
 NOR2x1_ASAP7_75t_R _24224_ (.A(net5744),
    .B(net5435),
    .Y(_01866_));
 OAI21x1_ASAP7_75t_R _24225_ (.A1(_01819_),
    .A2(_01866_),
    .B(net5726),
    .Y(_01867_));
 NOR2x1_ASAP7_75t_R _24226_ (.A(net5281),
    .B(net5435),
    .Y(_01868_));
 NOR2x1_ASAP7_75t_R _24227_ (.A(net5433),
    .B(net5724),
    .Y(_01869_));
 OAI21x1_ASAP7_75t_R _24228_ (.A1(_01868_),
    .A2(net5120),
    .B(net5723),
    .Y(_01870_));
 AOI21x1_ASAP7_75t_R _24229_ (.A1(_01867_),
    .A2(_01870_),
    .B(net5737),
    .Y(_01871_));
 OAI21x1_ASAP7_75t_R _24230_ (.A1(_01865_),
    .A2(_01871_),
    .B(net5421),
    .Y(_01872_));
 AOI21x1_ASAP7_75t_R _24232_ (.A1(_01872_),
    .A2(_01859_),
    .B(net6168),
    .Y(_01874_));
 AO21x1_ASAP7_75t_R _24235_ (.A1(net5718),
    .A2(_01226_),
    .B(net5738),
    .Y(_01877_));
 NAND2x1_ASAP7_75t_R _24236_ (.A(net5424),
    .B(_01877_),
    .Y(_01878_));
 AOI21x1_ASAP7_75t_R _24237_ (.A1(_01818_),
    .A2(net5437),
    .B(net5718),
    .Y(_01879_));
 NAND2x1_ASAP7_75t_R _24238_ (.A(net5742),
    .B(net5432),
    .Y(_01880_));
 AND2x2_ASAP7_75t_R _24239_ (.A(_01879_),
    .B(_01880_),
    .Y(_01881_));
 NOR2x1_ASAP7_75t_R _24240_ (.A(net5432),
    .B(net5727),
    .Y(_01882_));
 AOI21x1_ASAP7_75t_R _24241_ (.A1(net5419),
    .A2(_01882_),
    .B(net5428),
    .Y(_01883_));
 NAND2x1_ASAP7_75t_R _24242_ (.A(net5432),
    .B(net5718),
    .Y(_01884_));
 NOR2x1_ASAP7_75t_R _24243_ (.A(net5420),
    .B(_01884_),
    .Y(_01885_));
 INVx1_ASAP7_75t_R _24244_ (.A(_01885_),
    .Y(_01886_));
 NAND2x1_ASAP7_75t_R _24245_ (.A(_01883_),
    .B(_01886_),
    .Y(_01887_));
 AO21x1_ASAP7_75t_R _24246_ (.A1(_01671_),
    .A2(net5124),
    .B(net5740),
    .Y(_01888_));
 OAI21x1_ASAP7_75t_R _24247_ (.A1(_01881_),
    .A2(_01887_),
    .B(_01888_),
    .Y(_01889_));
 NOR2x1_ASAP7_75t_R _24248_ (.A(net5428),
    .B(net5422),
    .Y(_01890_));
 NOR2x1_ASAP7_75t_R _24249_ (.A(net5433),
    .B(net5746),
    .Y(_01891_));
 OAI21x1_ASAP7_75t_R _24250_ (.A1(_01866_),
    .A2(_01891_),
    .B(net5726),
    .Y(_01892_));
 AO31x2_ASAP7_75t_R _24251_ (.A1(_01890_),
    .A2(_01870_),
    .A3(_01892_),
    .B(net5715),
    .Y(_01893_));
 AOI21x1_ASAP7_75t_R _24252_ (.A1(_01878_),
    .A2(_01889_),
    .B(_01893_),
    .Y(_01894_));
 OAI21x1_ASAP7_75t_R _24253_ (.A1(_01874_),
    .A2(_01894_),
    .B(net6167),
    .Y(_01895_));
 NAND2x1_ASAP7_75t_R _24254_ (.A(net5433),
    .B(net5724),
    .Y(_01896_));
 NAND2x1_ASAP7_75t_R _24255_ (.A(net5719),
    .B(_01830_),
    .Y(_01897_));
 NAND3x1_ASAP7_75t_R _24256_ (.A(_01763_),
    .B(net5119),
    .C(_01897_),
    .Y(_01898_));
 OAI21x1_ASAP7_75t_R _24257_ (.A1(net5277),
    .A2(net5436),
    .B(_01722_),
    .Y(_01899_));
 AOI21x1_ASAP7_75t_R _24258_ (.A1(net5720),
    .A2(_01899_),
    .B(net5739),
    .Y(_01900_));
 AOI21x1_ASAP7_75t_R _24259_ (.A1(_01710_),
    .A2(_01900_),
    .B(net5422),
    .Y(_01901_));
 NAND2x1_ASAP7_75t_R _24260_ (.A(_01898_),
    .B(_01901_),
    .Y(_01902_));
 OAI21x1_ASAP7_75t_R _24261_ (.A1(_01817_),
    .A2(net5121),
    .B(net5720),
    .Y(_01903_));
 OAI21x1_ASAP7_75t_R _24262_ (.A1(_01868_),
    .A2(net5125),
    .B(net5726),
    .Y(_01904_));
 AOI21x1_ASAP7_75t_R _24263_ (.A1(_01903_),
    .A2(_01904_),
    .B(net5428),
    .Y(_01905_));
 NOR2x1_ASAP7_75t_R _24264_ (.A(net5742),
    .B(net5746),
    .Y(_01906_));
 OAI21x1_ASAP7_75t_R _24265_ (.A1(_01906_),
    .A2(_01869_),
    .B(net5726),
    .Y(_01907_));
 NAND2x1_ASAP7_75t_R _24266_ (.A(net5419),
    .B(_01882_),
    .Y(_01908_));
 AOI21x1_ASAP7_75t_R _24267_ (.A1(_01907_),
    .A2(_01908_),
    .B(net5738),
    .Y(_01909_));
 OAI21x1_ASAP7_75t_R _24269_ (.A1(_01905_),
    .A2(_01909_),
    .B(net5422),
    .Y(_01911_));
 AOI21x1_ASAP7_75t_R _24271_ (.A1(_01902_),
    .A2(_01911_),
    .B(net5715),
    .Y(_01913_));
 OAI21x1_ASAP7_75t_R _24272_ (.A1(_01707_),
    .A2(net4996),
    .B(net5722),
    .Y(_01914_));
 OAI21x1_ASAP7_75t_R _24273_ (.A1(_01821_),
    .A2(net5121),
    .B(net5733),
    .Y(_01915_));
 AOI21x1_ASAP7_75t_R _24274_ (.A1(_01914_),
    .A2(_01915_),
    .B(net5427),
    .Y(_01916_));
 INVx1_ASAP7_75t_R _24275_ (.A(_01744_),
    .Y(_01917_));
 NOR2x1_ASAP7_75t_R _24276_ (.A(net5742),
    .B(net5437),
    .Y(_01918_));
 OAI21x1_ASAP7_75t_R _24277_ (.A1(net4741),
    .A2(net5117),
    .B(net5732),
    .Y(_01919_));
 OAI21x1_ASAP7_75t_R _24278_ (.A1(_01866_),
    .A2(net5420),
    .B(net5723),
    .Y(_01920_));
 AOI21x1_ASAP7_75t_R _24279_ (.A1(_01919_),
    .A2(_01920_),
    .B(net5737),
    .Y(_01921_));
 OAI21x1_ASAP7_75t_R _24280_ (.A1(_01916_),
    .A2(_01921_),
    .B(net5424),
    .Y(_01922_));
 NAND2x1_ASAP7_75t_R _24281_ (.A(net5732),
    .B(_01854_),
    .Y(_01923_));
 INVx1_ASAP7_75t_R _24282_ (.A(_01219_),
    .Y(_01924_));
 OAI21x1_ASAP7_75t_R _24283_ (.A1(net5741),
    .A2(net6169),
    .B(_01924_),
    .Y(_01925_));
 INVx1_ASAP7_75t_R _24284_ (.A(_01925_),
    .Y(_01926_));
 NOR2x1_ASAP7_75t_R _24285_ (.A(net5435),
    .B(net5724),
    .Y(_01927_));
 OAI21x1_ASAP7_75t_R _24286_ (.A1(_01926_),
    .A2(_01927_),
    .B(net5723),
    .Y(_01928_));
 AOI21x1_ASAP7_75t_R _24287_ (.A1(_01923_),
    .A2(_01928_),
    .B(net5427),
    .Y(_01929_));
 NAND2x1_ASAP7_75t_R _24288_ (.A(net5732),
    .B(_01868_),
    .Y(_01930_));
 AOI21x1_ASAP7_75t_R _24290_ (.A1(_01930_),
    .A2(_01849_),
    .B(net5737),
    .Y(_01932_));
 OAI21x1_ASAP7_75t_R _24291_ (.A1(_01929_),
    .A2(_01932_),
    .B(net5421),
    .Y(_01933_));
 AOI21x1_ASAP7_75t_R _24292_ (.A1(_01922_),
    .A2(_01933_),
    .B(net6168),
    .Y(_01934_));
 OAI21x1_ASAP7_75t_R _24293_ (.A1(_01913_),
    .A2(_01934_),
    .B(_01845_),
    .Y(_01935_));
 NAND2x1_ASAP7_75t_R _24294_ (.A(_01935_),
    .B(_01895_),
    .Y(_00089_));
 OA21x2_ASAP7_75t_R _24295_ (.A1(net5723),
    .A2(_01228_),
    .B(net5737),
    .Y(_01936_));
 OAI21x1_ASAP7_75t_R _24296_ (.A1(net5742),
    .A2(net5431),
    .B(net5747),
    .Y(_01937_));
 NAND2x1_ASAP7_75t_R _24297_ (.A(net5723),
    .B(_01937_),
    .Y(_01938_));
 AOI21x1_ASAP7_75t_R _24298_ (.A1(_01936_),
    .A2(_01938_),
    .B(net5421),
    .Y(_01939_));
 OAI21x1_ASAP7_75t_R _24299_ (.A1(net5431),
    .A2(_01785_),
    .B(net5733),
    .Y(_01940_));
 NAND2x1_ASAP7_75t_R _24300_ (.A(_01223_),
    .B(net5723),
    .Y(_01941_));
 NAND3x1_ASAP7_75t_R _24301_ (.A(_01940_),
    .B(net5427),
    .C(_01941_),
    .Y(_01942_));
 AOI21x1_ASAP7_75t_R _24302_ (.A1(_01939_),
    .A2(_01942_),
    .B(_01733_),
    .Y(_01943_));
 AND2x2_ASAP7_75t_R _24303_ (.A(_01212_),
    .B(_01214_),
    .Y(_01944_));
 INVx1_ASAP7_75t_R _24304_ (.A(_01944_),
    .Y(_01945_));
 NAND2x1_ASAP7_75t_R _24305_ (.A(_01945_),
    .B(net5431),
    .Y(_01946_));
 AO21x1_ASAP7_75t_R _24306_ (.A1(_01793_),
    .A2(net4668),
    .B(net5728),
    .Y(_01947_));
 AOI21x1_ASAP7_75t_R _24307_ (.A1(net5124),
    .A2(_01671_),
    .B(net5428),
    .Y(_01948_));
 AO21x1_ASAP7_75t_R _24308_ (.A1(net4743),
    .A2(_01706_),
    .B(net5728),
    .Y(_01949_));
 AO21x1_ASAP7_75t_R _24309_ (.A1(_01949_),
    .A2(_01822_),
    .B(net5424),
    .Y(_01950_));
 AO21x1_ASAP7_75t_R _24310_ (.A1(_01947_),
    .A2(_01948_),
    .B(_01950_),
    .Y(_01951_));
 NAND2x1_ASAP7_75t_R _24311_ (.A(_01943_),
    .B(_01951_),
    .Y(_01952_));
 OA21x2_ASAP7_75t_R _24312_ (.A1(_01224_),
    .A2(net5723),
    .B(net5427),
    .Y(_01953_));
 OAI21x1_ASAP7_75t_R _24313_ (.A1(_01723_),
    .A2(net5127),
    .B(net5723),
    .Y(_01954_));
 AOI21x1_ASAP7_75t_R _24314_ (.A1(_01953_),
    .A2(_01954_),
    .B(net5424),
    .Y(_01955_));
 NAND2x1_ASAP7_75t_R _24315_ (.A(net5718),
    .B(_01834_),
    .Y(_01956_));
 AOI21x1_ASAP7_75t_R _24316_ (.A1(net5731),
    .A2(net4746),
    .B(net5428),
    .Y(_01957_));
 OAI21x1_ASAP7_75t_R _24317_ (.A1(_01866_),
    .A2(net4887),
    .B(_01957_),
    .Y(_01958_));
 AOI21x1_ASAP7_75t_R _24318_ (.A1(_01955_),
    .A2(_01958_),
    .B(net6168),
    .Y(_01959_));
 NAND2x1_ASAP7_75t_R _24319_ (.A(_01226_),
    .B(net5727),
    .Y(_01960_));
 OAI21x1_ASAP7_75t_R _24320_ (.A1(_01906_),
    .A2(_01869_),
    .B(net5721),
    .Y(_01961_));
 AOI21x1_ASAP7_75t_R _24321_ (.A1(_01960_),
    .A2(_01961_),
    .B(net5738),
    .Y(_01962_));
 AO21x1_ASAP7_75t_R _24322_ (.A1(_01789_),
    .A2(_01722_),
    .B(net5728),
    .Y(_01963_));
 AO21x1_ASAP7_75t_R _24323_ (.A1(_01839_),
    .A2(_01739_),
    .B(net5719),
    .Y(_01964_));
 AOI21x1_ASAP7_75t_R _24324_ (.A1(_01963_),
    .A2(_01964_),
    .B(net5429),
    .Y(_01965_));
 OAI21x1_ASAP7_75t_R _24325_ (.A1(_01962_),
    .A2(_01965_),
    .B(net5424),
    .Y(_01966_));
 AOI21x1_ASAP7_75t_R _24326_ (.A1(_01959_),
    .A2(_01966_),
    .B(net6167),
    .Y(_01967_));
 NAND2x1_ASAP7_75t_R _24327_ (.A(_01967_),
    .B(_01952_),
    .Y(_01968_));
 AO21x1_ASAP7_75t_R _24328_ (.A1(net4743),
    .A2(net5000),
    .B(net5732),
    .Y(_01969_));
 NOR2x1_ASAP7_75t_R _24329_ (.A(net5279),
    .B(net5433),
    .Y(_01970_));
 OAI21x1_ASAP7_75t_R _24330_ (.A1(_01970_),
    .A2(net5117),
    .B(net5732),
    .Y(_01971_));
 AOI21x1_ASAP7_75t_R _24331_ (.A1(_01969_),
    .A2(_01971_),
    .B(net5737),
    .Y(_01972_));
 NAND2x1_ASAP7_75t_R _24332_ (.A(_01764_),
    .B(net5723),
    .Y(_01973_));
 NOR2x1_ASAP7_75t_R _24333_ (.A(_01891_),
    .B(_01973_),
    .Y(_01974_));
 NAND2x1_ASAP7_75t_R _24334_ (.A(_01925_),
    .B(net5733),
    .Y(_01975_));
 OAI21x1_ASAP7_75t_R _24335_ (.A1(net5117),
    .A2(_01975_),
    .B(net5737),
    .Y(_01976_));
 NOR2x1_ASAP7_75t_R _24336_ (.A(_01974_),
    .B(_01976_),
    .Y(_01977_));
 OAI21x1_ASAP7_75t_R _24337_ (.A1(_01972_),
    .A2(_01977_),
    .B(net5421),
    .Y(_01978_));
 OA21x2_ASAP7_75t_R _24338_ (.A1(_01927_),
    .A2(net4670),
    .B(net5722),
    .Y(_01979_));
 OR2x2_ASAP7_75t_R _24339_ (.A(_01765_),
    .B(_01761_),
    .Y(_01980_));
 NOR2x1_ASAP7_75t_R _24340_ (.A(net5427),
    .B(_01765_),
    .Y(_01981_));
 NAND2x1_ASAP7_75t_R _24341_ (.A(_01706_),
    .B(net5723),
    .Y(_01982_));
 OAI21x1_ASAP7_75t_R _24342_ (.A1(net5117),
    .A2(_01982_),
    .B(_01975_),
    .Y(_01983_));
 AOI21x1_ASAP7_75t_R _24343_ (.A1(_01981_),
    .A2(_01983_),
    .B(net5421),
    .Y(_01984_));
 OAI21x1_ASAP7_75t_R _24344_ (.A1(_01979_),
    .A2(_01980_),
    .B(_01984_),
    .Y(_01985_));
 AOI21x1_ASAP7_75t_R _24345_ (.A1(_01978_),
    .A2(_01985_),
    .B(net6168),
    .Y(_01986_));
 OAI21x1_ASAP7_75t_R _24346_ (.A1(_01926_),
    .A2(_01868_),
    .B(net5732),
    .Y(_01987_));
 AOI21x1_ASAP7_75t_R _24347_ (.A1(_01987_),
    .A2(_01938_),
    .B(net5427),
    .Y(_01988_));
 OAI21x1_ASAP7_75t_R _24348_ (.A1(_01708_),
    .A2(_01982_),
    .B(net5427),
    .Y(_01989_));
 INVx1_ASAP7_75t_R _24349_ (.A(_01746_),
    .Y(_01990_));
 NOR2x1_ASAP7_75t_R _24350_ (.A(_01989_),
    .B(_01990_),
    .Y(_01991_));
 OAI21x1_ASAP7_75t_R _24351_ (.A1(_01988_),
    .A2(_01991_),
    .B(net5424),
    .Y(_01992_));
 OAI21x1_ASAP7_75t_R _24352_ (.A1(net4669),
    .A2(net5117),
    .B(net5723),
    .Y(_01993_));
 OAI21x1_ASAP7_75t_R _24353_ (.A1(net5747),
    .A2(net5431),
    .B(net4743),
    .Y(_01994_));
 NAND2x1_ASAP7_75t_R _24354_ (.A(net5733),
    .B(_01994_),
    .Y(_01995_));
 AOI21x1_ASAP7_75t_R _24355_ (.A1(_01993_),
    .A2(_01995_),
    .B(net5427),
    .Y(_01996_));
 NOR2x1_ASAP7_75t_R _24356_ (.A(net5277),
    .B(net5435),
    .Y(_01997_));
 OAI21x1_ASAP7_75t_R _24357_ (.A1(_01997_),
    .A2(_01848_),
    .B(net5723),
    .Y(_01998_));
 AOI21x1_ASAP7_75t_R _24358_ (.A1(_01940_),
    .A2(_01998_),
    .B(net5737),
    .Y(_01999_));
 OAI21x1_ASAP7_75t_R _24359_ (.A1(_01996_),
    .A2(_01999_),
    .B(net5421),
    .Y(_02000_));
 AOI21x1_ASAP7_75t_R _24360_ (.A1(_01992_),
    .A2(_02000_),
    .B(_01733_),
    .Y(_02001_));
 OAI21x1_ASAP7_75t_R _24361_ (.A1(_01986_),
    .A2(_02001_),
    .B(net6167),
    .Y(_02002_));
 NAND2x1_ASAP7_75t_R _24362_ (.A(_02002_),
    .B(_01968_),
    .Y(_00090_));
 INVx1_ASAP7_75t_R _24363_ (.A(net4893),
    .Y(_02003_));
 OAI21x1_ASAP7_75t_R _24364_ (.A1(_02003_),
    .A2(_01756_),
    .B(net5718),
    .Y(_02004_));
 AO21x1_ASAP7_75t_R _24365_ (.A1(net4744),
    .A2(net4889),
    .B(net5718),
    .Y(_02005_));
 AO21x1_ASAP7_75t_R _24366_ (.A1(_02004_),
    .A2(_02005_),
    .B(net5428),
    .Y(_02006_));
 INVx1_ASAP7_75t_R _24367_ (.A(_01714_),
    .Y(_02007_));
 AO21x1_ASAP7_75t_R _24368_ (.A1(_02007_),
    .A2(_01907_),
    .B(net5740),
    .Y(_02008_));
 AOI21x1_ASAP7_75t_R _24370_ (.A1(_02006_),
    .A2(_02008_),
    .B(net5424),
    .Y(_02010_));
 NOR2x1_ASAP7_75t_R _24371_ (.A(net5117),
    .B(_01975_),
    .Y(_02011_));
 AO21x1_ASAP7_75t_R _24372_ (.A1(_02011_),
    .A2(net5740),
    .B(net5422),
    .Y(_02012_));
 NAND2x1_ASAP7_75t_R _24373_ (.A(net5130),
    .B(net5434),
    .Y(_02013_));
 AOI21x1_ASAP7_75t_R _24375_ (.A1(_02013_),
    .A2(_01946_),
    .B(net5728),
    .Y(_02015_));
 AOI211x1_ASAP7_75t_R _24376_ (.A1(_01671_),
    .A2(net5124),
    .B(net4516),
    .C(net5740),
    .Y(_02016_));
 OAI21x1_ASAP7_75t_R _24377_ (.A1(_02012_),
    .A2(_02016_),
    .B(net5715),
    .Y(_02017_));
 NOR2x1_ASAP7_75t_R _24378_ (.A(_02010_),
    .B(_02017_),
    .Y(_02018_));
 INVx1_ASAP7_75t_R _24379_ (.A(_01766_),
    .Y(_02019_));
 NOR2x1_ASAP7_75t_R _24380_ (.A(net5721),
    .B(_02019_),
    .Y(_02020_));
 AOI21x1_ASAP7_75t_R _24381_ (.A1(net5422),
    .A2(_02020_),
    .B(_01680_),
    .Y(_02021_));
 AOI21x1_ASAP7_75t_R _24383_ (.A1(_01748_),
    .A2(net5119),
    .B(net5721),
    .Y(_02023_));
 OAI21x1_ASAP7_75t_R _24384_ (.A1(net4742),
    .A2(_02023_),
    .B(net5424),
    .Y(_02024_));
 AOI21x1_ASAP7_75t_R _24386_ (.A1(_02021_),
    .A2(_02024_),
    .B(net5428),
    .Y(_02026_));
 INVx1_ASAP7_75t_R _24387_ (.A(_01971_),
    .Y(_02027_));
 OAI21x1_ASAP7_75t_R _24389_ (.A1(net5731),
    .A2(net4891),
    .B(net5422),
    .Y(_02029_));
 OAI21x1_ASAP7_75t_R _24390_ (.A1(_02027_),
    .A2(_02029_),
    .B(net5428),
    .Y(_02030_));
 NAND2x1_ASAP7_75t_R _24391_ (.A(net4889),
    .B(net4668),
    .Y(_02031_));
 AOI21x1_ASAP7_75t_R _24392_ (.A1(net4743),
    .A2(_01712_),
    .B(net5719),
    .Y(_02032_));
 AOI211x1_ASAP7_75t_R _24393_ (.A1(_02031_),
    .A2(net5723),
    .B(_02032_),
    .C(net5422),
    .Y(_02033_));
 OAI21x1_ASAP7_75t_R _24394_ (.A1(_02030_),
    .A2(_02033_),
    .B(net6168),
    .Y(_02034_));
 OAI21x1_ASAP7_75t_R _24395_ (.A1(_02026_),
    .A2(_02034_),
    .B(net6167),
    .Y(_02035_));
 NAND2x1_ASAP7_75t_R _24396_ (.A(net5123),
    .B(net4745),
    .Y(_02036_));
 NAND2x1_ASAP7_75t_R _24397_ (.A(_01747_),
    .B(_01785_),
    .Y(_02037_));
 OA21x2_ASAP7_75t_R _24398_ (.A1(_02037_),
    .A2(net5718),
    .B(net5424),
    .Y(_02038_));
 OAI21x1_ASAP7_75t_R _24399_ (.A1(net5723),
    .A2(_01994_),
    .B(net5421),
    .Y(_02039_));
 OA21x2_ASAP7_75t_R _24400_ (.A1(_01997_),
    .A2(_01707_),
    .B(net5723),
    .Y(_02040_));
 OAI21x1_ASAP7_75t_R _24401_ (.A1(_02039_),
    .A2(_02040_),
    .B(net5427),
    .Y(_02041_));
 AOI21x1_ASAP7_75t_R _24402_ (.A1(_02036_),
    .A2(_02038_),
    .B(_02041_),
    .Y(_02042_));
 OAI21x1_ASAP7_75t_R _24403_ (.A1(net5732),
    .A2(net4741),
    .B(net5424),
    .Y(_02043_));
 OA21x2_ASAP7_75t_R _24404_ (.A1(net5120),
    .A2(net5117),
    .B(net5732),
    .Y(_02044_));
 OAI21x1_ASAP7_75t_R _24406_ (.A1(_02043_),
    .A2(_02044_),
    .B(net5737),
    .Y(_02046_));
 NAND2x1_ASAP7_75t_R _24407_ (.A(_01789_),
    .B(_01712_),
    .Y(_02047_));
 AOI21x1_ASAP7_75t_R _24408_ (.A1(net4999),
    .A2(_01711_),
    .B(net5729),
    .Y(_02048_));
 AOI211x1_ASAP7_75t_R _24409_ (.A1(_02047_),
    .A2(net5731),
    .B(_02048_),
    .C(net5424),
    .Y(_02049_));
 OAI21x1_ASAP7_75t_R _24410_ (.A1(_02046_),
    .A2(_02049_),
    .B(net6168),
    .Y(_02050_));
 OAI21x1_ASAP7_75t_R _24411_ (.A1(_02042_),
    .A2(_02050_),
    .B(_01845_),
    .Y(_02051_));
 NAND2x1_ASAP7_75t_R _24412_ (.A(_01884_),
    .B(_02037_),
    .Y(_02052_));
 OAI21x1_ASAP7_75t_R _24413_ (.A1(net5738),
    .A2(_02052_),
    .B(net5424),
    .Y(_02053_));
 OA21x2_ASAP7_75t_R _24414_ (.A1(_01970_),
    .A2(net4996),
    .B(net5732),
    .Y(_02054_));
 NAND2x1_ASAP7_75t_R _24415_ (.A(net5737),
    .B(_01928_),
    .Y(_02055_));
 NOR2x1_ASAP7_75t_R _24416_ (.A(_02054_),
    .B(_02055_),
    .Y(_02056_));
 OAI21x1_ASAP7_75t_R _24417_ (.A1(_02053_),
    .A2(_02056_),
    .B(net5715),
    .Y(_02057_));
 OA21x2_ASAP7_75t_R _24418_ (.A1(net4890),
    .A2(net4996),
    .B(net5732),
    .Y(_02058_));
 OA21x2_ASAP7_75t_R _24419_ (.A1(net5425),
    .A2(net5121),
    .B(net5722),
    .Y(_02059_));
 OAI21x1_ASAP7_75t_R _24420_ (.A1(_02058_),
    .A2(_02059_),
    .B(net5737),
    .Y(_02060_));
 NAND2x1_ASAP7_75t_R _24421_ (.A(net5728),
    .B(net4747),
    .Y(_02061_));
 OA21x2_ASAP7_75t_R _24422_ (.A1(_02061_),
    .A2(_01854_),
    .B(net5427),
    .Y(_02062_));
 OAI21x1_ASAP7_75t_R _24423_ (.A1(net4887),
    .A2(_02047_),
    .B(_02062_),
    .Y(_02063_));
 AOI21x1_ASAP7_75t_R _24424_ (.A1(_02063_),
    .A2(_02060_),
    .B(net5424),
    .Y(_02064_));
 NOR2x1_ASAP7_75t_R _24425_ (.A(_02057_),
    .B(_02064_),
    .Y(_02065_));
 OAI22x1_ASAP7_75t_R _24426_ (.A1(_02018_),
    .A2(_02035_),
    .B1(_02065_),
    .B2(_02051_),
    .Y(_00091_));
 NAND2x1_ASAP7_75t_R _24427_ (.A(net5726),
    .B(_01891_),
    .Y(_02066_));
 AOI21x1_ASAP7_75t_R _24428_ (.A1(net5733),
    .A2(_01821_),
    .B(net5428),
    .Y(_02067_));
 AND3x1_ASAP7_75t_R _24429_ (.A(_01870_),
    .B(_02066_),
    .C(_02067_),
    .Y(_02068_));
 AO21x1_ASAP7_75t_R _24430_ (.A1(_01880_),
    .A2(net4889),
    .B(net5718),
    .Y(_02069_));
 NOR2x1_ASAP7_75t_R _24431_ (.A(net5740),
    .B(_01882_),
    .Y(_02070_));
 AO21x1_ASAP7_75t_R _24432_ (.A1(_02069_),
    .A2(_02070_),
    .B(net5422),
    .Y(_02071_));
 OAI21x1_ASAP7_75t_R _24433_ (.A1(_02068_),
    .A2(_02071_),
    .B(net5715),
    .Y(_02072_));
 NOR2x1_ASAP7_75t_R _24434_ (.A(net5131),
    .B(net5433),
    .Y(_02073_));
 OA21x2_ASAP7_75t_R _24435_ (.A1(_02073_),
    .A2(net5719),
    .B(net5740),
    .Y(_02074_));
 AO21x1_ASAP7_75t_R _24436_ (.A1(net5420),
    .A2(net5437),
    .B(net5727),
    .Y(_02075_));
 AO21x1_ASAP7_75t_R _24437_ (.A1(_02074_),
    .A2(_02075_),
    .B(net5423),
    .Y(_02076_));
 AO21x1_ASAP7_75t_R _24438_ (.A1(net5281),
    .A2(net5432),
    .B(net5718),
    .Y(_02077_));
 OA21x2_ASAP7_75t_R _24439_ (.A1(net4568),
    .A2(_02077_),
    .B(_01836_),
    .Y(_02078_));
 NOR2x1_ASAP7_75t_R _24440_ (.A(_02076_),
    .B(_02078_),
    .Y(_02079_));
 OAI21x1_ASAP7_75t_R _24441_ (.A1(_02072_),
    .A2(_02079_),
    .B(net6167),
    .Y(_02080_));
 AND3x1_ASAP7_75t_R _24442_ (.A(net5123),
    .B(net5418),
    .C(net5725),
    .Y(_02081_));
 NOR2x1_ASAP7_75t_R _24443_ (.A(net5118),
    .B(net4896),
    .Y(_02082_));
 OR3x1_ASAP7_75t_R _24444_ (.A(_02081_),
    .B(net5429),
    .C(_02082_),
    .Y(_02083_));
 AND3x1_ASAP7_75t_R _24445_ (.A(_01784_),
    .B(_01741_),
    .C(net5429),
    .Y(_02084_));
 NOR2x1_ASAP7_75t_R _24446_ (.A(net5422),
    .B(_02084_),
    .Y(_02085_));
 INVx1_ASAP7_75t_R _24447_ (.A(net5127),
    .Y(_02086_));
 INVx1_ASAP7_75t_R _24448_ (.A(_01896_),
    .Y(_02087_));
 OAI22x1_ASAP7_75t_R _24449_ (.A1(_02086_),
    .A2(net5716),
    .B1(net4896),
    .B2(_02087_),
    .Y(_02088_));
 OAI21x1_ASAP7_75t_R _24450_ (.A1(net5278),
    .A2(net5719),
    .B(net5429),
    .Y(_02089_));
 AOI21x1_ASAP7_75t_R _24451_ (.A1(net5716),
    .A2(net4568),
    .B(_02089_),
    .Y(_02090_));
 AOI21x1_ASAP7_75t_R _24452_ (.A1(net5735),
    .A2(_02088_),
    .B(_02090_),
    .Y(_02091_));
 OAI21x1_ASAP7_75t_R _24453_ (.A1(net5423),
    .A2(_02091_),
    .B(net6168),
    .Y(_02092_));
 AOI21x1_ASAP7_75t_R _24454_ (.A1(_02083_),
    .A2(_02085_),
    .B(_02092_),
    .Y(_02093_));
 OA21x2_ASAP7_75t_R _24455_ (.A1(net4747),
    .A2(net5733),
    .B(net4892),
    .Y(_02094_));
 AOI21x1_ASAP7_75t_R _24456_ (.A1(_01763_),
    .A2(_02094_),
    .B(net5424),
    .Y(_02095_));
 AOI21x1_ASAP7_75t_R _24457_ (.A1(net5734),
    .A2(_01899_),
    .B(net5739),
    .Y(_02096_));
 NAND2x1_ASAP7_75t_R _24458_ (.A(_01690_),
    .B(_02096_),
    .Y(_02097_));
 AOI21x1_ASAP7_75t_R _24459_ (.A1(_02095_),
    .A2(_02097_),
    .B(net5715),
    .Y(_02098_));
 OAI21x1_ASAP7_75t_R _24460_ (.A1(net5120),
    .A2(_01708_),
    .B(net5720),
    .Y(_02099_));
 AOI21x1_ASAP7_75t_R _24461_ (.A1(_01987_),
    .A2(_02099_),
    .B(net5428),
    .Y(_02100_));
 AO21x1_ASAP7_75t_R _24462_ (.A1(_01830_),
    .A2(_01711_),
    .B(net5728),
    .Y(_02101_));
 AOI21x1_ASAP7_75t_R _24463_ (.A1(_01710_),
    .A2(_02101_),
    .B(net5740),
    .Y(_02102_));
 OAI21x1_ASAP7_75t_R _24464_ (.A1(_02100_),
    .A2(_02102_),
    .B(net5424),
    .Y(_02103_));
 NAND2x1_ASAP7_75t_R _24465_ (.A(_02103_),
    .B(_02098_),
    .Y(_02104_));
 OAI21x1_ASAP7_75t_R _24466_ (.A1(_01819_),
    .A2(_01927_),
    .B(net5720),
    .Y(_02105_));
 OAI21x1_ASAP7_75t_R _24467_ (.A1(net5425),
    .A2(_01891_),
    .B(net5726),
    .Y(_02106_));
 AOI21x1_ASAP7_75t_R _24468_ (.A1(_02105_),
    .A2(_02106_),
    .B(net5428),
    .Y(_02107_));
 AOI21x1_ASAP7_75t_R _24469_ (.A1(_01892_),
    .A2(_01961_),
    .B(net5738),
    .Y(_02108_));
 OAI21x1_ASAP7_75t_R _24470_ (.A1(_02107_),
    .A2(_02108_),
    .B(net5424),
    .Y(_02109_));
 NAND2x1_ASAP7_75t_R _24471_ (.A(net5739),
    .B(_01679_),
    .Y(_02110_));
 OA21x2_ASAP7_75t_R _24472_ (.A1(_01689_),
    .A2(_02110_),
    .B(net5422),
    .Y(_02111_));
 AO21x1_ASAP7_75t_R _24473_ (.A1(net5123),
    .A2(_01747_),
    .B(net5727),
    .Y(_02112_));
 AOI21x1_ASAP7_75t_R _24474_ (.A1(_01880_),
    .A2(_01879_),
    .B(net5740),
    .Y(_02113_));
 NAND2x1_ASAP7_75t_R _24475_ (.A(_02112_),
    .B(_02113_),
    .Y(_02114_));
 AOI21x1_ASAP7_75t_R _24476_ (.A1(_02111_),
    .A2(_02114_),
    .B(net6168),
    .Y(_02115_));
 AOI21x1_ASAP7_75t_R _24477_ (.A1(_02109_),
    .A2(_02115_),
    .B(net6167),
    .Y(_02116_));
 NAND2x1_ASAP7_75t_R _24478_ (.A(_02104_),
    .B(_02116_),
    .Y(_02117_));
 OAI21x1_ASAP7_75t_R _24479_ (.A1(_02080_),
    .A2(_02093_),
    .B(_02117_),
    .Y(_00092_));
 INVx1_ASAP7_75t_R _24480_ (.A(net5124),
    .Y(_02118_));
 OA21x2_ASAP7_75t_R _24481_ (.A1(_01823_),
    .A2(net5728),
    .B(net5427),
    .Y(_02119_));
 OA21x2_ASAP7_75t_R _24482_ (.A1(net5719),
    .A2(_02118_),
    .B(_02119_),
    .Y(_02120_));
 NAND2x1p5_ASAP7_75t_R _24483_ (.A(net4744),
    .B(net5728),
    .Y(_02121_));
 INVx1_ASAP7_75t_R _24484_ (.A(_01801_),
    .Y(_02122_));
 OA21x2_ASAP7_75t_R _24485_ (.A1(_02121_),
    .A2(_02122_),
    .B(net5740),
    .Y(_02123_));
 AO21x1_ASAP7_75t_R _24486_ (.A1(_01748_),
    .A2(net4743),
    .B(net5733),
    .Y(_02124_));
 AO21x1_ASAP7_75t_R _24487_ (.A1(_02123_),
    .A2(_02124_),
    .B(net5421),
    .Y(_02125_));
 AOI21x1_ASAP7_75t_R _24488_ (.A1(_01802_),
    .A2(_01763_),
    .B(net5423),
    .Y(_02126_));
 NOR2x1_ASAP7_75t_R _24489_ (.A(net4888),
    .B(net5435),
    .Y(_02127_));
 OA21x2_ASAP7_75t_R _24490_ (.A1(_02127_),
    .A2(net5728),
    .B(net5427),
    .Y(_02128_));
 OAI21x1_ASAP7_75t_R _24491_ (.A1(_02118_),
    .A2(_01940_),
    .B(_02128_),
    .Y(_02129_));
 AOI21x1_ASAP7_75t_R _24492_ (.A1(_02126_),
    .A2(_02129_),
    .B(_01733_),
    .Y(_02130_));
 OAI21x1_ASAP7_75t_R _24493_ (.A1(_02120_),
    .A2(_02125_),
    .B(_02130_),
    .Y(_02131_));
 NOR2x1_ASAP7_75t_R _24494_ (.A(net5718),
    .B(_01747_),
    .Y(_02132_));
 OAI21x1_ASAP7_75t_R _24495_ (.A1(_01926_),
    .A2(_01854_),
    .B(net5732),
    .Y(_02133_));
 OA21x2_ASAP7_75t_R _24496_ (.A1(_01748_),
    .A2(net5734),
    .B(net5739),
    .Y(_02134_));
 AOI21x1_ASAP7_75t_R _24497_ (.A1(_02133_),
    .A2(_02134_),
    .B(net5422),
    .Y(_02135_));
 OAI21x1_ASAP7_75t_R _24498_ (.A1(_02132_),
    .A2(_01762_),
    .B(_02135_),
    .Y(_02136_));
 NAND2x1_ASAP7_75t_R _24499_ (.A(_01767_),
    .B(_01808_),
    .Y(_02137_));
 AOI21x1_ASAP7_75t_R _24500_ (.A1(net5279),
    .A2(net5436),
    .B(net5721),
    .Y(_02138_));
 AOI21x1_ASAP7_75t_R _24501_ (.A1(net5119),
    .A2(_02138_),
    .B(net5429),
    .Y(_02139_));
 NAND2x1_ASAP7_75t_R _24502_ (.A(_02137_),
    .B(_02139_),
    .Y(_02140_));
 OA21x2_ASAP7_75t_R _24503_ (.A1(net5742),
    .A2(net5727),
    .B(net5429),
    .Y(_02141_));
 AOI21x1_ASAP7_75t_R _24504_ (.A1(_02141_),
    .A2(_01786_),
    .B(net5423),
    .Y(_02142_));
 AOI21x1_ASAP7_75t_R _24505_ (.A1(_02140_),
    .A2(_02142_),
    .B(net6168),
    .Y(_02143_));
 AOI21x1_ASAP7_75t_R _24506_ (.A1(_02136_),
    .A2(_02143_),
    .B(_01845_),
    .Y(_02144_));
 NAND2x1_ASAP7_75t_R _24507_ (.A(_02144_),
    .B(_02131_),
    .Y(_02145_));
 OA21x2_ASAP7_75t_R _24508_ (.A1(_01862_),
    .A2(net5128),
    .B(net5719),
    .Y(_02146_));
 AOI211x1_ASAP7_75t_R _24509_ (.A1(_01676_),
    .A2(_02138_),
    .B(_02146_),
    .C(net5429),
    .Y(_02147_));
 OAI21x1_ASAP7_75t_R _24510_ (.A1(net4886),
    .A2(_01737_),
    .B(_01835_),
    .Y(_02148_));
 OAI21x1_ASAP7_75t_R _24511_ (.A1(net5739),
    .A2(_02148_),
    .B(net5422),
    .Y(_02149_));
 NAND2x1_ASAP7_75t_R _24512_ (.A(_02077_),
    .B(_01883_),
    .Y(_02150_));
 OA21x2_ASAP7_75t_R _24513_ (.A1(net4996),
    .A2(net5718),
    .B(net5428),
    .Y(_02151_));
 AOI21x1_ASAP7_75t_R _24514_ (.A1(_02004_),
    .A2(_02151_),
    .B(net5422),
    .Y(_02152_));
 AOI21x1_ASAP7_75t_R _24515_ (.A1(_02150_),
    .A2(_02152_),
    .B(net6168),
    .Y(_02153_));
 OAI21x1_ASAP7_75t_R _24516_ (.A1(_02147_),
    .A2(_02149_),
    .B(_02153_),
    .Y(_02154_));
 INVx1_ASAP7_75t_R _24517_ (.A(_01767_),
    .Y(_02155_));
 OA21x2_ASAP7_75t_R _24518_ (.A1(_02155_),
    .A2(_01819_),
    .B(_01975_),
    .Y(_02156_));
 OA21x2_ASAP7_75t_R _24519_ (.A1(net4747),
    .A2(net5728),
    .B(net5737),
    .Y(_02157_));
 AO21x1_ASAP7_75t_R _24520_ (.A1(net5119),
    .A2(net4894),
    .B(net5721),
    .Y(_02158_));
 AOI21x1_ASAP7_75t_R _24521_ (.A1(_02157_),
    .A2(_02158_),
    .B(net5422),
    .Y(_02159_));
 OAI21x1_ASAP7_75t_R _24522_ (.A1(net5740),
    .A2(_02156_),
    .B(_02159_),
    .Y(_02160_));
 OA21x2_ASAP7_75t_R _24523_ (.A1(net5724),
    .A2(net5726),
    .B(net5428),
    .Y(_02161_));
 AOI21x1_ASAP7_75t_R _24524_ (.A1(_02106_),
    .A2(_02161_),
    .B(net5424),
    .Y(_02162_));
 OAI21x1_ASAP7_75t_R _24525_ (.A1(net4890),
    .A2(_01854_),
    .B(net5723),
    .Y(_02163_));
 OAI21x1_ASAP7_75t_R _24526_ (.A1(net5125),
    .A2(net5420),
    .B(net5726),
    .Y(_02164_));
 NAND3x1_ASAP7_75t_R _24527_ (.A(_02163_),
    .B(net5737),
    .C(_02164_),
    .Y(_02165_));
 AOI21x1_ASAP7_75t_R _24528_ (.A1(_02162_),
    .A2(_02165_),
    .B(net5715),
    .Y(_02166_));
 AOI21x1_ASAP7_75t_R _24529_ (.A1(_02160_),
    .A2(_02166_),
    .B(net6167),
    .Y(_02167_));
 NAND2x1_ASAP7_75t_R _24530_ (.A(_02154_),
    .B(_02167_),
    .Y(_02168_));
 NAND2x1_ASAP7_75t_R _24531_ (.A(_02145_),
    .B(_02168_),
    .Y(_00093_));
 AO21x1_ASAP7_75t_R _24532_ (.A1(net4892),
    .A2(net4894),
    .B(net5729),
    .Y(_02169_));
 NAND2x1_ASAP7_75t_R _24533_ (.A(_02169_),
    .B(_02067_),
    .Y(_02170_));
 NAND2x1_ASAP7_75t_R _24534_ (.A(_01221_),
    .B(_01227_),
    .Y(_02171_));
 AOI21x1_ASAP7_75t_R _24535_ (.A1(_02171_),
    .A2(net5725),
    .B(net5736),
    .Y(_02172_));
 OAI21x1_ASAP7_75t_R _24536_ (.A1(net5426),
    .A2(net4887),
    .B(_02172_),
    .Y(_02173_));
 NAND2x1_ASAP7_75t_R _24537_ (.A(_02170_),
    .B(_02173_),
    .Y(_02174_));
 AOI21x1_ASAP7_75t_R _24538_ (.A1(net5422),
    .A2(_02174_),
    .B(net6168),
    .Y(_02175_));
 NAND2x1_ASAP7_75t_R _24539_ (.A(net5116),
    .B(net5433),
    .Y(_02176_));
 AOI21x1_ASAP7_75t_R _24540_ (.A1(_02176_),
    .A2(_02013_),
    .B(net5719),
    .Y(_02177_));
 AOI21x1_ASAP7_75t_R _24541_ (.A1(net4897),
    .A2(_01793_),
    .B(net5728),
    .Y(_02178_));
 OAI21x1_ASAP7_75t_R _24542_ (.A1(net4667),
    .A2(_02178_),
    .B(net5429),
    .Y(_02179_));
 NAND2x1_ASAP7_75t_R _24543_ (.A(net4888),
    .B(net5435),
    .Y(_02180_));
 AOI21x1_ASAP7_75t_R _24544_ (.A1(net4892),
    .A2(_02180_),
    .B(net5728),
    .Y(_02181_));
 AOI21x1_ASAP7_75t_R _24545_ (.A1(net4999),
    .A2(_01880_),
    .B(net5719),
    .Y(_02182_));
 OAI21x1_ASAP7_75t_R _24546_ (.A1(_02181_),
    .A2(_02182_),
    .B(net5736),
    .Y(_02183_));
 NAND3x1_ASAP7_75t_R _24547_ (.A(_02179_),
    .B(net5423),
    .C(_02183_),
    .Y(_02184_));
 AOI21x1_ASAP7_75t_R _24548_ (.A1(_02175_),
    .A2(_02184_),
    .B(net6167),
    .Y(_02185_));
 AO21x1_ASAP7_75t_R _24549_ (.A1(net4890),
    .A2(net5729),
    .B(net5429),
    .Y(_02186_));
 NOR2x1_ASAP7_75t_R _24550_ (.A(net5425),
    .B(_01897_),
    .Y(_02187_));
 OAI21x1_ASAP7_75t_R _24551_ (.A1(_02186_),
    .A2(_02187_),
    .B(net5423),
    .Y(_02188_));
 AOI21x1_ASAP7_75t_R _24552_ (.A1(net5733),
    .A2(_01917_),
    .B(net5740),
    .Y(_02189_));
 OAI21x1_ASAP7_75t_R _24553_ (.A1(net5721),
    .A2(net4668),
    .B(_02189_),
    .Y(_02190_));
 OAI21x1_ASAP7_75t_R _24554_ (.A1(net5437),
    .A2(_01785_),
    .B(net5718),
    .Y(_02191_));
 NOR2x1_ASAP7_75t_R _24555_ (.A(net5121),
    .B(net5115),
    .Y(_02192_));
 NOR2x1_ASAP7_75t_R _24556_ (.A(_02190_),
    .B(_02192_),
    .Y(_02193_));
 NOR2x1_ASAP7_75t_R _24557_ (.A(_02188_),
    .B(_02193_),
    .Y(_02194_));
 NOR2x1_ASAP7_75t_R _24558_ (.A(_02073_),
    .B(_02121_),
    .Y(_02195_));
 AOI21x1_ASAP7_75t_R _24559_ (.A1(_01839_),
    .A2(_01838_),
    .B(net5727),
    .Y(_02196_));
 OAI21x1_ASAP7_75t_R _24560_ (.A1(_02195_),
    .A2(_02196_),
    .B(net5429),
    .Y(_02197_));
 NOR2x1_ASAP7_75t_R _24561_ (.A(net5429),
    .B(_02020_),
    .Y(_02198_));
 NAND2x1_ASAP7_75t_R _24562_ (.A(_01941_),
    .B(_01940_),
    .Y(_02199_));
 NAND2x1_ASAP7_75t_R _24563_ (.A(_02198_),
    .B(_02199_),
    .Y(_02200_));
 AOI21x1_ASAP7_75t_R _24564_ (.A1(_02197_),
    .A2(_02200_),
    .B(net5423),
    .Y(_02201_));
 OAI21x1_ASAP7_75t_R _24565_ (.A1(_02194_),
    .A2(_02201_),
    .B(net6168),
    .Y(_02202_));
 NOR2x1_ASAP7_75t_R _24566_ (.A(_02087_),
    .B(_01688_),
    .Y(_02203_));
 OAI21x1_ASAP7_75t_R _24567_ (.A1(net5132),
    .A2(_02203_),
    .B(net5735),
    .Y(_02204_));
 AND2x2_ASAP7_75t_R _24568_ (.A(_01989_),
    .B(net5424),
    .Y(_02205_));
 NAND2x1_ASAP7_75t_R _24569_ (.A(_02204_),
    .B(_02205_),
    .Y(_02206_));
 AO21x1_ASAP7_75t_R _24570_ (.A1(net5121),
    .A2(net5728),
    .B(net5429),
    .Y(_02207_));
 NOR2x1_ASAP7_75t_R _24571_ (.A(net4566),
    .B(_01802_),
    .Y(_02208_));
 OAI21x1_ASAP7_75t_R _24572_ (.A1(net5129),
    .A2(net5430),
    .B(net5727),
    .Y(_02209_));
 AOI21x1_ASAP7_75t_R _24573_ (.A1(_01222_),
    .A2(net5718),
    .B(net5736),
    .Y(_02210_));
 OAI21x1_ASAP7_75t_R _24574_ (.A1(_02087_),
    .A2(_02209_),
    .B(_02210_),
    .Y(_02211_));
 OAI21x1_ASAP7_75t_R _24575_ (.A1(_02207_),
    .A2(_02208_),
    .B(_02211_),
    .Y(_02212_));
 AOI21x1_ASAP7_75t_R _24576_ (.A1(net5422),
    .A2(_02212_),
    .B(net5715),
    .Y(_02213_));
 AOI21x1_ASAP7_75t_R _24577_ (.A1(_02206_),
    .A2(_02213_),
    .B(_01845_),
    .Y(_02214_));
 NAND2x1_ASAP7_75t_R _24578_ (.A(net5725),
    .B(net5122),
    .Y(_02215_));
 NAND2x1_ASAP7_75t_R _24579_ (.A(net5717),
    .B(_01783_),
    .Y(_02216_));
 NAND2x1_ASAP7_75t_R _24580_ (.A(_02215_),
    .B(_02216_),
    .Y(_02217_));
 AOI21x1_ASAP7_75t_R _24581_ (.A1(_01712_),
    .A2(_02217_),
    .B(net5429),
    .Y(_02218_));
 NAND2x1_ASAP7_75t_R _24582_ (.A(net5724),
    .B(net5727),
    .Y(_02219_));
 NAND2x1_ASAP7_75t_R _24583_ (.A(net5417),
    .B(_02037_),
    .Y(_02220_));
 OAI21x1_ASAP7_75t_R _24584_ (.A1(net5735),
    .A2(_02220_),
    .B(net5422),
    .Y(_02221_));
 NOR2x1_ASAP7_75t_R _24585_ (.A(_02218_),
    .B(_02221_),
    .Y(_02222_));
 AO21x1_ASAP7_75t_R _24586_ (.A1(_01830_),
    .A2(net5716),
    .B(net5429),
    .Y(_02223_));
 AND2x2_ASAP7_75t_R _24587_ (.A(_01804_),
    .B(net5725),
    .Y(_02224_));
 OAI21x1_ASAP7_75t_R _24588_ (.A1(_02223_),
    .A2(_02224_),
    .B(net5423),
    .Y(_02225_));
 NAND2x1_ASAP7_75t_R _24589_ (.A(net5734),
    .B(net4566),
    .Y(_02226_));
 AND3x1_ASAP7_75t_R _24590_ (.A(_02004_),
    .B(net5429),
    .C(_02226_),
    .Y(_02227_));
 NOR2x1_ASAP7_75t_R _24591_ (.A(_02225_),
    .B(_02227_),
    .Y(_02228_));
 OAI21x1_ASAP7_75t_R _24592_ (.A1(_02222_),
    .A2(_02228_),
    .B(net5715),
    .Y(_02229_));
 AOI22x1_ASAP7_75t_R _24593_ (.A1(_02185_),
    .A2(_02202_),
    .B1(_02214_),
    .B2(_02229_),
    .Y(_00094_));
 AND3x1_ASAP7_75t_R _24594_ (.A(net5719),
    .B(net4744),
    .C(net4999),
    .Y(_02230_));
 AOI21x1_ASAP7_75t_R _24595_ (.A1(_01811_),
    .A2(net5119),
    .B(_02230_),
    .Y(_02231_));
 INVx1_ASAP7_75t_R _24596_ (.A(_02189_),
    .Y(_02232_));
 AO21x1_ASAP7_75t_R _24597_ (.A1(_01683_),
    .A2(_01682_),
    .B(_01227_),
    .Y(_02233_));
 OAI21x1_ASAP7_75t_R _24598_ (.A1(net5717),
    .A2(net4892),
    .B(_02233_),
    .Y(_02234_));
 OAI21x1_ASAP7_75t_R _24599_ (.A1(_02232_),
    .A2(_02234_),
    .B(net5423),
    .Y(_02235_));
 AOI21x1_ASAP7_75t_R _24600_ (.A1(net5740),
    .A2(_02231_),
    .B(_02235_),
    .Y(_02236_));
 AND3x1_ASAP7_75t_R _24601_ (.A(_01669_),
    .B(_01668_),
    .C(_01218_),
    .Y(_02237_));
 OAI21x1_ASAP7_75t_R _24602_ (.A1(_02237_),
    .A2(_01718_),
    .B(net5422),
    .Y(_02238_));
 NAND2x1_ASAP7_75t_R _24603_ (.A(net5739),
    .B(_02219_),
    .Y(_02239_));
 AOI211x1_ASAP7_75t_R _24604_ (.A1(net5123),
    .A2(_01736_),
    .B(_02239_),
    .C(_02132_),
    .Y(_02240_));
 OAI21x1_ASAP7_75t_R _24605_ (.A1(_02238_),
    .A2(_02240_),
    .B(net6168),
    .Y(_02241_));
 OAI21x1_ASAP7_75t_R _24606_ (.A1(_02236_),
    .A2(_02241_),
    .B(_01845_),
    .Y(_02242_));
 AOI21x1_ASAP7_75t_R _24607_ (.A1(net5119),
    .A2(_01793_),
    .B(net5719),
    .Y(_02243_));
 OAI21x1_ASAP7_75t_R _24608_ (.A1(_02015_),
    .A2(_02243_),
    .B(net5736),
    .Y(_02244_));
 AOI21x1_ASAP7_75t_R _24609_ (.A1(_01711_),
    .A2(_01793_),
    .B(net5719),
    .Y(_02245_));
 OA21x2_ASAP7_75t_R _24610_ (.A1(_01824_),
    .A2(_01766_),
    .B(net5719),
    .Y(_02246_));
 OAI21x1_ASAP7_75t_R _24611_ (.A1(_02245_),
    .A2(_02246_),
    .B(net5429),
    .Y(_02247_));
 AOI21x1_ASAP7_75t_R _24612_ (.A1(_02244_),
    .A2(_02247_),
    .B(net5423),
    .Y(_02248_));
 AO21x1_ASAP7_75t_R _24613_ (.A1(net5128),
    .A2(net5728),
    .B(net5429),
    .Y(_02249_));
 NOR2x1_ASAP7_75t_R _24614_ (.A(net5425),
    .B(_01956_),
    .Y(_02250_));
 OAI21x1_ASAP7_75t_R _24615_ (.A1(_02249_),
    .A2(_02250_),
    .B(net5423),
    .Y(_02251_));
 AOI211x1_ASAP7_75t_R _24616_ (.A1(net5721),
    .A2(_01891_),
    .B(_01718_),
    .C(_01821_),
    .Y(_02252_));
 OAI21x1_ASAP7_75t_R _24617_ (.A1(_02251_),
    .A2(_02252_),
    .B(net5715),
    .Y(_02253_));
 NOR2x1_ASAP7_75t_R _24618_ (.A(_02248_),
    .B(_02253_),
    .Y(_02254_));
 NAND2x1_ASAP7_75t_R _24619_ (.A(net5742),
    .B(net5727),
    .Y(_02255_));
 AO21x1_ASAP7_75t_R _24620_ (.A1(_02112_),
    .A2(_02255_),
    .B(net5428),
    .Y(_02256_));
 NAND2x1_ASAP7_75t_R _24621_ (.A(net5428),
    .B(_01961_),
    .Y(_02257_));
 OA21x2_ASAP7_75t_R _24622_ (.A1(_01848_),
    .A2(_01927_),
    .B(net5726),
    .Y(_02258_));
 OA21x2_ASAP7_75t_R _24623_ (.A1(_02257_),
    .A2(_02258_),
    .B(net5422),
    .Y(_02259_));
 AO21x1_ASAP7_75t_R _24624_ (.A1(net4997),
    .A2(net5727),
    .B(net5740),
    .Y(_02260_));
 OAI21x1_ASAP7_75t_R _24625_ (.A1(_01885_),
    .A2(_02260_),
    .B(net5424),
    .Y(_02261_));
 OA21x2_ASAP7_75t_R _24626_ (.A1(_01848_),
    .A2(net4997),
    .B(net5727),
    .Y(_02262_));
 NAND2x1_ASAP7_75t_R _24627_ (.A(net5740),
    .B(_02191_),
    .Y(_02263_));
 NOR2x1_ASAP7_75t_R _24628_ (.A(_02262_),
    .B(_02263_),
    .Y(_02264_));
 OAI21x1_ASAP7_75t_R _24629_ (.A1(_02261_),
    .A2(_02264_),
    .B(net6168),
    .Y(_02265_));
 AOI21x1_ASAP7_75t_R _24630_ (.A1(_02256_),
    .A2(_02259_),
    .B(_02265_),
    .Y(_02266_));
 AOI21x1_ASAP7_75t_R _24631_ (.A1(_01722_),
    .A2(_02176_),
    .B(net5728),
    .Y(_02267_));
 OAI21x1_ASAP7_75t_R _24632_ (.A1(_02267_),
    .A2(_02032_),
    .B(net5736),
    .Y(_02268_));
 AOI21x1_ASAP7_75t_R _24633_ (.A1(net5126),
    .A2(_01830_),
    .B(net5728),
    .Y(_02269_));
 OAI21x1_ASAP7_75t_R _24634_ (.A1(_02177_),
    .A2(_02269_),
    .B(net5429),
    .Y(_02270_));
 AOI21x1_ASAP7_75t_R _24635_ (.A1(_02268_),
    .A2(_02270_),
    .B(net5421),
    .Y(_02271_));
 AO21x1_ASAP7_75t_R _24636_ (.A1(_01841_),
    .A2(net5725),
    .B(net5736),
    .Y(_02272_));
 OAI21x1_ASAP7_75t_R _24637_ (.A1(_02203_),
    .A2(_02272_),
    .B(net5421),
    .Y(_02273_));
 AOI21x1_ASAP7_75t_R _24638_ (.A1(_01711_),
    .A2(_01793_),
    .B(net5728),
    .Y(_02274_));
 OA21x2_ASAP7_75t_R _24639_ (.A1(net5745),
    .A2(net5434),
    .B(net5742),
    .Y(_02275_));
 OAI21x1_ASAP7_75t_R _24640_ (.A1(net5719),
    .A2(_02275_),
    .B(net5736),
    .Y(_02276_));
 NOR2x1_ASAP7_75t_R _24641_ (.A(_02274_),
    .B(_02276_),
    .Y(_02277_));
 OAI21x1_ASAP7_75t_R _24642_ (.A1(_02273_),
    .A2(_02277_),
    .B(net5715),
    .Y(_02278_));
 OAI21x1_ASAP7_75t_R _24643_ (.A1(_02271_),
    .A2(_02278_),
    .B(net6167),
    .Y(_02279_));
 OAI22x1_ASAP7_75t_R _24644_ (.A1(_02242_),
    .A2(_02254_),
    .B1(_02266_),
    .B2(_02279_),
    .Y(_00095_));
 NOR2x1_ASAP7_75t_R _24645_ (.A(net6671),
    .B(_00468_),
    .Y(_02280_));
 XOR2x2_ASAP7_75t_R _24646_ (.A(_00678_),
    .B(net6568),
    .Y(_02281_));
 INVx1_ASAP7_75t_R _24647_ (.A(net6565),
    .Y(_02282_));
 XOR2x2_ASAP7_75t_R _24648_ (.A(_02281_),
    .B(_02282_),
    .Y(_02283_));
 XOR2x2_ASAP7_75t_R _24649_ (.A(_10719_),
    .B(net6417),
    .Y(_02284_));
 NAND2x1_ASAP7_75t_R _24650_ (.A(_02283_),
    .B(_02284_),
    .Y(_02285_));
 XOR2x2_ASAP7_75t_R _24651_ (.A(_02281_),
    .B(net6565),
    .Y(_02286_));
 XOR2x2_ASAP7_75t_R _24652_ (.A(net6417),
    .B(_10717_),
    .Y(_02287_));
 NAND2x1p5_ASAP7_75t_R _24653_ (.A(_02287_),
    .B(_02286_),
    .Y(_02288_));
 AOI21x1_ASAP7_75t_R _24654_ (.A1(_02288_),
    .A2(_02285_),
    .B(net6462),
    .Y(_02289_));
 OAI21x1_ASAP7_75t_R _24655_ (.A1(_02280_),
    .A2(_02289_),
    .B(net6513),
    .Y(_02290_));
 AND2x2_ASAP7_75t_R _24656_ (.A(net6462),
    .B(_00468_),
    .Y(_02291_));
 NAND2x1_ASAP7_75t_R _24657_ (.A(_02286_),
    .B(_02284_),
    .Y(_02292_));
 NAND2x1p5_ASAP7_75t_R _24658_ (.A(_02287_),
    .B(_02283_),
    .Y(_02293_));
 AOI21x1_ASAP7_75t_R _24659_ (.A1(_02293_),
    .A2(_02292_),
    .B(net6462),
    .Y(_02294_));
 INVx1_ASAP7_75t_R _24660_ (.A(net6513),
    .Y(_02295_));
 OAI21x1_ASAP7_75t_R _24661_ (.A1(_02291_),
    .A2(net6352),
    .B(_02295_),
    .Y(_02296_));
 NAND2x1_ASAP7_75t_R _24662_ (.A(_02290_),
    .B(_02296_),
    .Y(_02297_));
 INVx1_ASAP7_75t_R _24664_ (.A(net6592),
    .Y(_02298_));
 XOR2x2_ASAP7_75t_R _24665_ (.A(net6650),
    .B(net6622),
    .Y(_02299_));
 NAND2x1_ASAP7_75t_R _24666_ (.A(_02298_),
    .B(_02299_),
    .Y(_02300_));
 INVx1_ASAP7_75t_R _24667_ (.A(_02299_),
    .Y(_02301_));
 NAND2x1_ASAP7_75t_R _24668_ (.A(net6592),
    .B(_02301_),
    .Y(_02302_));
 INVx2_ASAP7_75t_R _24669_ (.A(_02281_),
    .Y(_02303_));
 AOI21x1_ASAP7_75t_R _24670_ (.A1(_02300_),
    .A2(_02302_),
    .B(_02303_),
    .Y(_02304_));
 XOR2x2_ASAP7_75t_R _24671_ (.A(net6622),
    .B(net6592),
    .Y(_02305_));
 NOR2x1_ASAP7_75t_R _24672_ (.A(net6650),
    .B(_02305_),
    .Y(_02306_));
 XNOR2x2_ASAP7_75t_R _24673_ (.A(net6622),
    .B(net6592),
    .Y(_02307_));
 NOR2x1_ASAP7_75t_R _24674_ (.A(net6416),
    .B(_02307_),
    .Y(_02308_));
 OAI21x1_ASAP7_75t_R _24675_ (.A1(_02306_),
    .A2(_02308_),
    .B(_02303_),
    .Y(_02309_));
 INVx1_ASAP7_75t_R _24676_ (.A(_02309_),
    .Y(_02310_));
 OAI21x1_ASAP7_75t_R _24677_ (.A1(_02310_),
    .A2(_02304_),
    .B(net6671),
    .Y(_02311_));
 INVx1_ASAP7_75t_R _24678_ (.A(net6514),
    .Y(_02312_));
 NOR2x1_ASAP7_75t_R _24679_ (.A(net6671),
    .B(_00469_),
    .Y(_02313_));
 INVx1_ASAP7_75t_R _24680_ (.A(_02313_),
    .Y(_02314_));
 NAND3x1_ASAP7_75t_R _24681_ (.A(net6166),
    .B(_02312_),
    .C(_02314_),
    .Y(_02315_));
 AO21x1_ASAP7_75t_R _24682_ (.A1(net6166),
    .A2(_02314_),
    .B(_02312_),
    .Y(_02316_));
 NAND2x1_ASAP7_75t_R _24683_ (.A(_02315_),
    .B(_02316_),
    .Y(_01237_));
 NOR2x1_ASAP7_75t_R _24684_ (.A(net6671),
    .B(_00470_),
    .Y(_02317_));
 INVx1_ASAP7_75t_R _24685_ (.A(_02317_),
    .Y(_02318_));
 XOR2x2_ASAP7_75t_R _24686_ (.A(_00577_),
    .B(_00609_),
    .Y(_02319_));
 XOR2x2_ASAP7_75t_R _24687_ (.A(net6418),
    .B(net6564),
    .Y(_02320_));
 NOR2x1_ASAP7_75t_R _24688_ (.A(_02319_),
    .B(_02320_),
    .Y(_02321_));
 INVx1_ASAP7_75t_R _24689_ (.A(net6564),
    .Y(_02322_));
 NOR2x1_ASAP7_75t_R _24690_ (.A(_02322_),
    .B(net6418),
    .Y(_02323_));
 AND2x4_ASAP7_75t_R _24691_ (.A(net6418),
    .B(_02322_),
    .Y(_02324_));
 OAI21x1_ASAP7_75t_R _24692_ (.A1(_02323_),
    .A2(_02324_),
    .B(_02319_),
    .Y(_02325_));
 INVx2_ASAP7_75t_R _24693_ (.A(_02325_),
    .Y(_02326_));
 OAI21x1_ASAP7_75t_R _24694_ (.A1(_02321_),
    .A2(_02326_),
    .B(net6671),
    .Y(_02327_));
 INVx1_ASAP7_75t_R _24695_ (.A(net6538),
    .Y(_02328_));
 AOI21x1_ASAP7_75t_R _24696_ (.A1(_02318_),
    .A2(_02327_),
    .B(_02328_),
    .Y(_02329_));
 NAND2x1_ASAP7_75t_R _24697_ (.A(_00470_),
    .B(net6462),
    .Y(_02330_));
 INVx1_ASAP7_75t_R _24698_ (.A(_02319_),
    .Y(_02331_));
 XOR2x2_ASAP7_75t_R _24699_ (.A(net6418),
    .B(_02322_),
    .Y(_02332_));
 NAND2x1_ASAP7_75t_R _24700_ (.A(_02331_),
    .B(_02332_),
    .Y(_02333_));
 NAND3x1_ASAP7_75t_R _24701_ (.A(_02333_),
    .B(_02325_),
    .C(net6671),
    .Y(_02334_));
 AOI21x1_ASAP7_75t_R _24702_ (.A1(_02330_),
    .A2(_02334_),
    .B(net6538),
    .Y(_02335_));
 NOR2x2_ASAP7_75t_R _24703_ (.A(_02329_),
    .B(_02335_),
    .Y(_02336_));
 OAI21x1_ASAP7_75t_R _24705_ (.A1(_02289_),
    .A2(_02280_),
    .B(_02295_),
    .Y(_02337_));
 OAI21x1_ASAP7_75t_R _24706_ (.A1(_02294_),
    .A2(_02291_),
    .B(net6513),
    .Y(_02338_));
 NAND2x2_ASAP7_75t_R _24707_ (.A(_02338_),
    .B(_02337_),
    .Y(_01230_));
 AOI21x1_ASAP7_75t_R _24708_ (.A1(_02318_),
    .A2(_02327_),
    .B(net6538),
    .Y(_02339_));
 AOI21x1_ASAP7_75t_R _24709_ (.A1(_02330_),
    .A2(_02334_),
    .B(_02328_),
    .Y(_02340_));
 NOR2x2_ASAP7_75t_R _24711_ (.A(_02339_),
    .B(_02340_),
    .Y(_02342_));
 XOR2x2_ASAP7_75t_R _24713_ (.A(net6561),
    .B(_00677_),
    .Y(_02343_));
 XOR2x2_ASAP7_75t_R _24714_ (.A(_02343_),
    .B(net6594),
    .Y(_02344_));
 XOR2x2_ASAP7_75t_R _24715_ (.A(_02344_),
    .B(_10857_),
    .Y(_02345_));
 NOR2x1_ASAP7_75t_R _24716_ (.A(net6655),
    .B(_00561_),
    .Y(_02346_));
 AO21x1_ASAP7_75t_R _24717_ (.A1(_02345_),
    .A2(net6671),
    .B(_02346_),
    .Y(_02347_));
 XOR2x2_ASAP7_75t_R _24718_ (.A(_02347_),
    .B(net6534),
    .Y(_02348_));
 XOR2x2_ASAP7_75t_R _24720_ (.A(net6563),
    .B(net6560),
    .Y(_02350_));
 XOR2x2_ASAP7_75t_R _24721_ (.A(_10800_),
    .B(_02350_),
    .Y(_02351_));
 NAND2x1_ASAP7_75t_R _24722_ (.A(_13603_),
    .B(_02351_),
    .Y(_02352_));
 OA21x2_ASAP7_75t_R _24723_ (.A1(_02351_),
    .A2(_13603_),
    .B(net6671),
    .Y(_02353_));
 AND2x2_ASAP7_75t_R _24724_ (.A(net6462),
    .B(_00563_),
    .Y(_02354_));
 AOI21x1_ASAP7_75t_R _24725_ (.A1(_02352_),
    .A2(_02353_),
    .B(_02354_),
    .Y(_02355_));
 XOR2x2_ASAP7_75t_R _24726_ (.A(_02355_),
    .B(net6536),
    .Y(_02356_));
 INVx2_ASAP7_75t_R _24727_ (.A(_02356_),
    .Y(_02357_));
 INVx1_ASAP7_75t_R _24730_ (.A(net6563),
    .Y(_02360_));
 XOR2x2_ASAP7_75t_R _24731_ (.A(_13583_),
    .B(_02360_),
    .Y(_02361_));
 XNOR2x2_ASAP7_75t_R _24732_ (.A(_00673_),
    .B(net6560),
    .Y(_02362_));
 XOR2x2_ASAP7_75t_R _24733_ (.A(_00578_),
    .B(_00610_),
    .Y(_02363_));
 XOR2x2_ASAP7_75t_R _24734_ (.A(_02362_),
    .B(_02363_),
    .Y(_02364_));
 AOI21x1_ASAP7_75t_R _24735_ (.A1(_02361_),
    .A2(_02364_),
    .B(net6462),
    .Y(_02365_));
 NOR2x1_ASAP7_75t_R _24736_ (.A(_02361_),
    .B(_02364_),
    .Y(_02366_));
 INVx1_ASAP7_75t_R _24737_ (.A(_02366_),
    .Y(_02367_));
 AND2x2_ASAP7_75t_R _24738_ (.A(net6462),
    .B(_00564_),
    .Y(_02368_));
 AOI21x1_ASAP7_75t_R _24739_ (.A1(_02365_),
    .A2(_02367_),
    .B(_02368_),
    .Y(_02369_));
 XOR2x2_ASAP7_75t_R _24740_ (.A(_02369_),
    .B(net6537),
    .Y(_02370_));
 INVx1_ASAP7_75t_R _24742_ (.A(_01235_),
    .Y(_02372_));
 OAI21x1_ASAP7_75t_R _24743_ (.A1(net5710),
    .A2(net6164),
    .B(_02372_),
    .Y(_02373_));
 NAND2x1_ASAP7_75t_R _24744_ (.A(net5702),
    .B(_02373_),
    .Y(_02374_));
 NOR2x1_ASAP7_75t_R _24745_ (.A(net5416),
    .B(net5413),
    .Y(_02375_));
 INVx2_ASAP7_75t_R _24746_ (.A(_02370_),
    .Y(_02376_));
 OAI21x1_ASAP7_75t_R _24749_ (.A1(net5710),
    .A2(net6164),
    .B(net5058),
    .Y(_02379_));
 NAND2x1_ASAP7_75t_R _24750_ (.A(net5411),
    .B(_02379_),
    .Y(_02380_));
 OAI21x1_ASAP7_75t_R _24751_ (.A1(net5712),
    .A2(net6165),
    .B(net4722),
    .Y(_02381_));
 INVx2_ASAP7_75t_R _24752_ (.A(net4565),
    .Y(_02382_));
 OAI22x1_ASAP7_75t_R _24753_ (.A1(net4446),
    .A2(_02375_),
    .B1(_02380_),
    .B2(net4468),
    .Y(_02383_));
 INVx1_ASAP7_75t_R _24754_ (.A(_02311_),
    .Y(_02384_));
 OAI21x1_ASAP7_75t_R _24755_ (.A1(_02313_),
    .A2(_02384_),
    .B(_02312_),
    .Y(_02385_));
 NAND3x1_ASAP7_75t_R _24756_ (.A(_02311_),
    .B(net6514),
    .C(_02314_),
    .Y(_02386_));
 NAND2x1p5_ASAP7_75t_R _24757_ (.A(_02386_),
    .B(_02385_),
    .Y(_02387_));
 AOI21x1_ASAP7_75t_R _24758_ (.A1(net5113),
    .A2(net5414),
    .B(net5409),
    .Y(_02388_));
 INVx1_ASAP7_75t_R _24759_ (.A(_02388_),
    .Y(_02389_));
 INVx1_ASAP7_75t_R _24760_ (.A(_02339_),
    .Y(_02390_));
 NAND3x1_ASAP7_75t_R _24761_ (.A(_02327_),
    .B(net6538),
    .C(_02318_),
    .Y(_02391_));
 AOI21x1_ASAP7_75t_R _24762_ (.A1(_02390_),
    .A2(_02391_),
    .B(_02372_),
    .Y(_02392_));
 INVx2_ASAP7_75t_R _24763_ (.A(net5712),
    .Y(_02393_));
 NAND3x1_ASAP7_75t_R _24764_ (.A(_02327_),
    .B(_02328_),
    .C(_02318_),
    .Y(_02394_));
 AOI21x1_ASAP7_75t_R _24765_ (.A1(_02393_),
    .A2(_02394_),
    .B(net4804),
    .Y(_02395_));
 OAI21x1_ASAP7_75t_R _24768_ (.A1(_02392_),
    .A2(net4666),
    .B(net5411),
    .Y(_02398_));
 AOI21x1_ASAP7_75t_R _24770_ (.A1(_02389_),
    .A2(_02398_),
    .B(net5708),
    .Y(_02400_));
 AOI21x1_ASAP7_75t_R _24771_ (.A1(net5708),
    .A2(_02383_),
    .B(_02400_),
    .Y(_02401_));
 INVx1_ASAP7_75t_R _24772_ (.A(_10776_),
    .Y(_02402_));
 XOR2x2_ASAP7_75t_R _24773_ (.A(_10743_),
    .B(_10803_),
    .Y(_02403_));
 NOR2x1_ASAP7_75t_R _24774_ (.A(_02402_),
    .B(_02403_),
    .Y(_02404_));
 XOR2x2_ASAP7_75t_R _24775_ (.A(_10743_),
    .B(net6561),
    .Y(_02405_));
 NOR2x1_ASAP7_75t_R _24776_ (.A(_10776_),
    .B(_02405_),
    .Y(_02406_));
 OAI21x1_ASAP7_75t_R _24777_ (.A1(_02404_),
    .A2(_02406_),
    .B(net6671),
    .Y(_02407_));
 NOR2x1_ASAP7_75t_R _24778_ (.A(net6655),
    .B(_00562_),
    .Y(_02408_));
 INVx1_ASAP7_75t_R _24779_ (.A(_02408_),
    .Y(_02409_));
 NAND3x1_ASAP7_75t_R _24780_ (.A(_02407_),
    .B(net6535),
    .C(_02409_),
    .Y(_02410_));
 AO21x1_ASAP7_75t_R _24781_ (.A1(_02407_),
    .A2(_02409_),
    .B(net6535),
    .Y(_02411_));
 NAND2x1_ASAP7_75t_R _24782_ (.A(_02410_),
    .B(_02411_),
    .Y(_02412_));
 INVx1_ASAP7_75t_R _24783_ (.A(_02412_),
    .Y(_02413_));
 OAI21x1_ASAP7_75t_R _24786_ (.A1(net6163),
    .A2(_02401_),
    .B(net5405),
    .Y(_02416_));
 INVx1_ASAP7_75t_R _24787_ (.A(_01238_),
    .Y(_02417_));
 NOR2x1_ASAP7_75t_R _24789_ (.A(_02417_),
    .B(net5414),
    .Y(_02419_));
 INVx1_ASAP7_75t_R _24790_ (.A(_02419_),
    .Y(_02420_));
 INVx1_ASAP7_75t_R _24791_ (.A(_01231_),
    .Y(_02421_));
 AO21x1_ASAP7_75t_R _24792_ (.A1(_02391_),
    .A2(_02390_),
    .B(_02421_),
    .Y(_02422_));
 AO21x1_ASAP7_75t_R _24795_ (.A1(_02420_),
    .A2(_02422_),
    .B(net5703),
    .Y(_02425_));
 AO21x1_ASAP7_75t_R _24796_ (.A1(_02391_),
    .A2(_02390_),
    .B(net5059),
    .Y(_02426_));
 NOR2x1_ASAP7_75t_R _24797_ (.A(net5410),
    .B(_02382_),
    .Y(_02427_));
 AOI21x1_ASAP7_75t_R _24798_ (.A1(_02426_),
    .A2(_02427_),
    .B(net5709),
    .Y(_02428_));
 NOR2x1_ASAP7_75t_R _24799_ (.A(net5714),
    .B(net5416),
    .Y(_02429_));
 OAI21x1_ASAP7_75t_R _24800_ (.A1(net5113),
    .A2(net5414),
    .B(net5706),
    .Y(_02430_));
 NOR2x1_ASAP7_75t_R _24801_ (.A(net5112),
    .B(net4885),
    .Y(_02431_));
 NAND2x1_ASAP7_75t_R _24803_ (.A(net5714),
    .B(net5113),
    .Y(_02432_));
 NAND2x1_ASAP7_75t_R _24804_ (.A(net5416),
    .B(net5413),
    .Y(_02433_));
 NAND2x1_ASAP7_75t_R _24805_ (.A(_02432_),
    .B(_02433_),
    .Y(_02434_));
 OAI21x1_ASAP7_75t_R _24807_ (.A1(net5703),
    .A2(_02434_),
    .B(net5707),
    .Y(_02436_));
 OAI21x1_ASAP7_75t_R _24808_ (.A1(_02431_),
    .A2(_02436_),
    .B(net6163),
    .Y(_02437_));
 AOI21x1_ASAP7_75t_R _24809_ (.A1(_02425_),
    .A2(_02428_),
    .B(_02437_),
    .Y(_02438_));
 XOR2x2_ASAP7_75t_R _24810_ (.A(_13623_),
    .B(net6445),
    .Y(_02439_));
 XOR2x2_ASAP7_75t_R _24811_ (.A(_02439_),
    .B(_10697_),
    .Y(_02440_));
 NOR2x1_ASAP7_75t_R _24812_ (.A(net6655),
    .B(_00560_),
    .Y(_02441_));
 AO21x1_ASAP7_75t_R _24813_ (.A1(_02440_),
    .A2(net6671),
    .B(_02441_),
    .Y(_02442_));
 XOR2x2_ASAP7_75t_R _24814_ (.A(_02442_),
    .B(_00844_),
    .Y(_02443_));
 OAI21x1_ASAP7_75t_R _24815_ (.A1(_02416_),
    .A2(_02438_),
    .B(_02443_),
    .Y(_02444_));
 INVx1_ASAP7_75t_R _24816_ (.A(_01241_),
    .Y(_02445_));
 AO21x1_ASAP7_75t_R _24817_ (.A1(_02394_),
    .A2(_02393_),
    .B(_02445_),
    .Y(_02446_));
 AOI21x1_ASAP7_75t_R _24818_ (.A1(net5113),
    .A2(net5414),
    .B(net5706),
    .Y(_02447_));
 NAND2x1_ASAP7_75t_R _24819_ (.A(net5711),
    .B(net5412),
    .Y(_02448_));
 INVx1_ASAP7_75t_R _24820_ (.A(_02374_),
    .Y(_02449_));
 AOI221x1_ASAP7_75t_R _24823_ (.A1(net4665),
    .A2(_02447_),
    .B1(_02448_),
    .B2(_02449_),
    .C(net6162),
    .Y(_02452_));
 AO21x1_ASAP7_75t_R _24824_ (.A1(_02394_),
    .A2(_02393_),
    .B(net5059),
    .Y(_02453_));
 AND2x2_ASAP7_75t_R _24825_ (.A(_02447_),
    .B(_02453_),
    .Y(_02454_));
 NOR2x1_ASAP7_75t_R _24826_ (.A(net5714),
    .B(net5412),
    .Y(_02455_));
 NAND2x1_ASAP7_75t_R _24827_ (.A(net5704),
    .B(_02455_),
    .Y(_02456_));
 INVx1_ASAP7_75t_R _24829_ (.A(_01233_),
    .Y(_02458_));
 OA21x2_ASAP7_75t_R _24830_ (.A1(net6165),
    .A2(net5712),
    .B(_02458_),
    .Y(_02459_));
 NAND2x1_ASAP7_75t_R _24831_ (.A(net5702),
    .B(_02459_),
    .Y(_02460_));
 NAND3x1_ASAP7_75t_R _24833_ (.A(_02456_),
    .B(_02460_),
    .C(net6162),
    .Y(_02462_));
 INVx1_ASAP7_75t_R _24834_ (.A(_02348_),
    .Y(_02463_));
 OAI21x1_ASAP7_75t_R _24836_ (.A1(_02454_),
    .A2(_02462_),
    .B(net5698),
    .Y(_02465_));
 NOR2x1_ASAP7_75t_R _24837_ (.A(_02452_),
    .B(_02465_),
    .Y(_02466_));
 INVx1_ASAP7_75t_R _24838_ (.A(net4723),
    .Y(_02467_));
 OAI21x1_ASAP7_75t_R _24839_ (.A1(net5712),
    .A2(net6165),
    .B(net4562),
    .Y(_02468_));
 AO21x1_ASAP7_75t_R _24841_ (.A1(_02422_),
    .A2(_02468_),
    .B(net5703),
    .Y(_02470_));
 OA21x2_ASAP7_75t_R _24842_ (.A1(net6164),
    .A2(net5710),
    .B(_01238_),
    .Y(_02471_));
 NAND2x1_ASAP7_75t_R _24843_ (.A(net5703),
    .B(_02471_),
    .Y(_02472_));
 AOI21x1_ASAP7_75t_R _24845_ (.A1(_02393_),
    .A2(_02394_),
    .B(_02421_),
    .Y(_02474_));
 AOI21x1_ASAP7_75t_R _24846_ (.A1(net5705),
    .A2(net4512),
    .B(net5709),
    .Y(_02475_));
 AND3x1_ASAP7_75t_R _24847_ (.A(_02470_),
    .B(_02472_),
    .C(_02475_),
    .Y(_02476_));
 OAI21x1_ASAP7_75t_R _24849_ (.A1(net5710),
    .A2(net6164),
    .B(net4722),
    .Y(_02478_));
 NAND2x1p5_ASAP7_75t_R _24850_ (.A(_02478_),
    .B(net5406),
    .Y(_02479_));
 INVx2_ASAP7_75t_R _24851_ (.A(_02479_),
    .Y(_02480_));
 NOR2x1_ASAP7_75t_R _24852_ (.A(net5409),
    .B(net4565),
    .Y(_02481_));
 AOI211x1_ASAP7_75t_R _24853_ (.A1(net5703),
    .A2(_02455_),
    .B(_02480_),
    .C(_02481_),
    .Y(_02482_));
 OAI21x1_ASAP7_75t_R _24854_ (.A1(net6162),
    .A2(_02482_),
    .B(net6163),
    .Y(_02483_));
 OAI21x1_ASAP7_75t_R _24857_ (.A1(_02476_),
    .A2(_02483_),
    .B(net5700),
    .Y(_02486_));
 NOR2x1_ASAP7_75t_R _24858_ (.A(_02466_),
    .B(_02486_),
    .Y(_02487_));
 INVx1_ASAP7_75t_R _24859_ (.A(_01236_),
    .Y(_02488_));
 OAI21x1_ASAP7_75t_R _24860_ (.A1(net5710),
    .A2(net6164),
    .B(_02488_),
    .Y(_02489_));
 NOR2x1_ASAP7_75t_R _24861_ (.A(net5409),
    .B(_02489_),
    .Y(_02490_));
 AO21x1_ASAP7_75t_R _24862_ (.A1(_02447_),
    .A2(_02453_),
    .B(net5708),
    .Y(_02491_));
 NOR2x1_ASAP7_75t_R _24863_ (.A(_02490_),
    .B(_02491_),
    .Y(_02492_));
 INVx1_ASAP7_75t_R _24865_ (.A(_01239_),
    .Y(_02494_));
 OAI21x1_ASAP7_75t_R _24866_ (.A1(net5712),
    .A2(net6165),
    .B(_02494_),
    .Y(_02495_));
 NAND2x2_ASAP7_75t_R _24868_ (.A(net4565),
    .B(net5409),
    .Y(_02497_));
 OA21x2_ASAP7_75t_R _24869_ (.A1(net5409),
    .A2(net4663),
    .B(_02497_),
    .Y(_02498_));
 NOR2x1_ASAP7_75t_R _24870_ (.A(net6162),
    .B(_02490_),
    .Y(_02499_));
 AO21x1_ASAP7_75t_R _24871_ (.A1(_02498_),
    .A2(_02499_),
    .B(net6163),
    .Y(_02500_));
 OAI21x1_ASAP7_75t_R _24873_ (.A1(net5712),
    .A2(net6165),
    .B(net4806),
    .Y(_02502_));
 OAI21x1_ASAP7_75t_R _24874_ (.A1(net5408),
    .A2(_02502_),
    .B(net6162),
    .Y(_02503_));
 NOR2x1_ASAP7_75t_R _24875_ (.A(_02490_),
    .B(_02503_),
    .Y(_02504_));
 NOR2x1_ASAP7_75t_R _24876_ (.A(net4809),
    .B(_02336_),
    .Y(_02505_));
 INVx1_ASAP7_75t_R _24877_ (.A(_02505_),
    .Y(_02506_));
 OAI21x1_ASAP7_75t_R _24878_ (.A1(net5710),
    .A2(net6164),
    .B(_02458_),
    .Y(_02507_));
 NOR2x1_ASAP7_75t_R _24879_ (.A(net5409),
    .B(_02507_),
    .Y(_02508_));
 AOI21x1_ASAP7_75t_R _24880_ (.A1(_02447_),
    .A2(_02506_),
    .B(_02508_),
    .Y(_02509_));
 NAND2x1_ASAP7_75t_R _24881_ (.A(_02504_),
    .B(_02509_),
    .Y(_02510_));
 INVx1_ASAP7_75t_R _24882_ (.A(_01246_),
    .Y(_02511_));
 OAI21x1_ASAP7_75t_R _24884_ (.A1(net5710),
    .A2(net6164),
    .B(_02467_),
    .Y(_02513_));
 NAND2x1p5_ASAP7_75t_R _24885_ (.A(_02513_),
    .B(net5704),
    .Y(_02514_));
 OAI21x1_ASAP7_75t_R _24886_ (.A1(_02511_),
    .A2(net5704),
    .B(net4433),
    .Y(_02515_));
 AOI21x1_ASAP7_75t_R _24887_ (.A1(net5708),
    .A2(_02515_),
    .B(_02463_),
    .Y(_02516_));
 AOI21x1_ASAP7_75t_R _24889_ (.A1(_02510_),
    .A2(_02516_),
    .B(net5405),
    .Y(_02518_));
 OAI21x1_ASAP7_75t_R _24890_ (.A1(_02492_),
    .A2(_02500_),
    .B(_02518_),
    .Y(_02519_));
 AO21x1_ASAP7_75t_R _24891_ (.A1(net5412),
    .A2(net4804),
    .B(net5702),
    .Y(_02520_));
 NOR2x1_ASAP7_75t_R _24892_ (.A(_02421_),
    .B(net5412),
    .Y(_02521_));
 OAI21x1_ASAP7_75t_R _24893_ (.A1(net4514),
    .A2(_02521_),
    .B(net5702),
    .Y(_02522_));
 AOI21x1_ASAP7_75t_R _24895_ (.A1(_02520_),
    .A2(_02522_),
    .B(net6162),
    .Y(_02524_));
 NOR2x1_ASAP7_75t_R _24896_ (.A(net5113),
    .B(net5414),
    .Y(_02525_));
 OAI21x1_ASAP7_75t_R _24897_ (.A1(net4881),
    .A2(_02525_),
    .B(net5407),
    .Y(_02526_));
 AOI21x1_ASAP7_75t_R _24898_ (.A1(net5412),
    .A2(net5714),
    .B(_02376_),
    .Y(_02527_));
 NAND2x1_ASAP7_75t_R _24899_ (.A(_02513_),
    .B(_02527_),
    .Y(_02528_));
 AOI21x1_ASAP7_75t_R _24900_ (.A1(_02526_),
    .A2(_02528_),
    .B(net5708),
    .Y(_02529_));
 OAI21x1_ASAP7_75t_R _24901_ (.A1(_02524_),
    .A2(_02529_),
    .B(_02463_),
    .Y(_02530_));
 AOI21x1_ASAP7_75t_R _24902_ (.A1(net5407),
    .A2(net4513),
    .B(net6162),
    .Y(_02531_));
 AOI21x1_ASAP7_75t_R _24903_ (.A1(_02393_),
    .A2(_02394_),
    .B(_02372_),
    .Y(_02532_));
 OAI21x1_ASAP7_75t_R _24905_ (.A1(_02532_),
    .A2(net4881),
    .B(net5705),
    .Y(_02534_));
 AOI21x1_ASAP7_75t_R _24906_ (.A1(_02531_),
    .A2(_02534_),
    .B(_02463_),
    .Y(_02535_));
 AOI21x1_ASAP7_75t_R _24907_ (.A1(_02390_),
    .A2(_02391_),
    .B(net5060),
    .Y(_02536_));
 OAI21x1_ASAP7_75t_R _24909_ (.A1(_02532_),
    .A2(net4880),
    .B(net5407),
    .Y(_02538_));
 NAND3x1_ASAP7_75t_R _24911_ (.A(_02538_),
    .B(_02460_),
    .C(net6162),
    .Y(_02540_));
 AOI21x1_ASAP7_75t_R _24912_ (.A1(_02535_),
    .A2(_02540_),
    .B(net5700),
    .Y(_02541_));
 AOI21x1_ASAP7_75t_R _24913_ (.A1(_02530_),
    .A2(_02541_),
    .B(_02443_),
    .Y(_02542_));
 NAND2x1_ASAP7_75t_R _24914_ (.A(_02542_),
    .B(_02519_),
    .Y(_02543_));
 OAI21x1_ASAP7_75t_R _24915_ (.A1(_02444_),
    .A2(_02487_),
    .B(_02543_),
    .Y(_00096_));
 INVx1_ASAP7_75t_R _24916_ (.A(_02443_),
    .Y(_02544_));
 OA21x2_ASAP7_75t_R _24918_ (.A1(net6165),
    .A2(net5712),
    .B(_02445_),
    .Y(_02546_));
 INVx1_ASAP7_75t_R _24919_ (.A(_02507_),
    .Y(_02547_));
 OA21x2_ASAP7_75t_R _24920_ (.A1(_02546_),
    .A2(_02547_),
    .B(net5705),
    .Y(_02548_));
 OA21x2_ASAP7_75t_R _24922_ (.A1(net6164),
    .A2(net5710),
    .B(net5059),
    .Y(_02550_));
 OAI21x1_ASAP7_75t_R _24923_ (.A1(_02382_),
    .A2(_02550_),
    .B(net5411),
    .Y(_02551_));
 NAND2x1_ASAP7_75t_R _24924_ (.A(net5707),
    .B(_02551_),
    .Y(_02552_));
 NOR2x1_ASAP7_75t_R _24925_ (.A(_02548_),
    .B(_02552_),
    .Y(_02553_));
 AO21x1_ASAP7_75t_R _24926_ (.A1(net4564),
    .A2(net5408),
    .B(net5708),
    .Y(_02554_));
 INVx1_ASAP7_75t_R _24927_ (.A(_02453_),
    .Y(_02555_));
 NOR2x1_ASAP7_75t_R _24928_ (.A(_02555_),
    .B(_02389_),
    .Y(_02556_));
 OAI21x1_ASAP7_75t_R _24929_ (.A1(_02554_),
    .A2(_02556_),
    .B(net5700),
    .Y(_02557_));
 OAI21x1_ASAP7_75t_R _24931_ (.A1(net5411),
    .A2(_02433_),
    .B(net5707),
    .Y(_02559_));
 OAI21x1_ASAP7_75t_R _24932_ (.A1(_02505_),
    .A2(net4466),
    .B(net4445),
    .Y(_02560_));
 NOR2x1_ASAP7_75t_R _24933_ (.A(_02559_),
    .B(_02560_),
    .Y(_02561_));
 INVx1_ASAP7_75t_R _24934_ (.A(_02395_),
    .Y(_02562_));
 NAND2x1_ASAP7_75t_R _24935_ (.A(net5714),
    .B(_02336_),
    .Y(_02563_));
 AOI21x1_ASAP7_75t_R _24936_ (.A1(_02562_),
    .A2(_02563_),
    .B(net5703),
    .Y(_02564_));
 NOR2x1_ASAP7_75t_R _24937_ (.A(net4809),
    .B(net5412),
    .Y(_02565_));
 OAI21x1_ASAP7_75t_R _24938_ (.A1(_02565_),
    .A2(net4885),
    .B(net6162),
    .Y(_02566_));
 OAI21x1_ASAP7_75t_R _24939_ (.A1(net4443),
    .A2(_02566_),
    .B(net5405),
    .Y(_02567_));
 OAI22x1_ASAP7_75t_R _24940_ (.A1(_02553_),
    .A2(_02557_),
    .B1(_02561_),
    .B2(_02567_),
    .Y(_02568_));
 NOR2x1_ASAP7_75t_R _24941_ (.A(net6162),
    .B(_02564_),
    .Y(_02569_));
 NOR2x1_ASAP7_75t_R _24942_ (.A(net5711),
    .B(net5412),
    .Y(_02570_));
 NOR2x1_ASAP7_75t_R _24943_ (.A(_02570_),
    .B(net4885),
    .Y(_02571_));
 NOR2x1_ASAP7_75t_R _24944_ (.A(net5404),
    .B(_02571_),
    .Y(_02572_));
 INVx1_ASAP7_75t_R _24945_ (.A(_01248_),
    .Y(_02573_));
 NAND2x1_ASAP7_75t_R _24946_ (.A(net5411),
    .B(net5700),
    .Y(_02574_));
 OAI21x1_ASAP7_75t_R _24947_ (.A1(_02573_),
    .A2(_02574_),
    .B(net6162),
    .Y(_02575_));
 INVx1_ASAP7_75t_R _24948_ (.A(net5059),
    .Y(_02576_));
 AO21x1_ASAP7_75t_R _24949_ (.A1(_02394_),
    .A2(_02393_),
    .B(_02576_),
    .Y(_02577_));
 INVx1_ASAP7_75t_R _24950_ (.A(_02471_),
    .Y(_02578_));
 AOI21x1_ASAP7_75t_R _24951_ (.A1(_02577_),
    .A2(_02578_),
    .B(net5411),
    .Y(_02579_));
 OAI21x1_ASAP7_75t_R _24952_ (.A1(_02575_),
    .A2(_02579_),
    .B(net6163),
    .Y(_02580_));
 AND2x2_ASAP7_75t_R _24953_ (.A(_02373_),
    .B(net5410),
    .Y(_02581_));
 OAI21x1_ASAP7_75t_R _24954_ (.A1(net4809),
    .A2(net5412),
    .B(net5706),
    .Y(_02582_));
 NOR2x1_ASAP7_75t_R _24955_ (.A(net6162),
    .B(net5701),
    .Y(_02583_));
 OAI21x1_ASAP7_75t_R _24956_ (.A1(_02375_),
    .A2(_02582_),
    .B(_02583_),
    .Y(_02584_));
 AOI21x1_ASAP7_75t_R _24957_ (.A1(net4882),
    .A2(net4442),
    .B(_02584_),
    .Y(_02585_));
 AOI211x1_ASAP7_75t_R _24958_ (.A1(net4426),
    .A2(_02572_),
    .B(_02580_),
    .C(_02585_),
    .Y(_02586_));
 AOI21x1_ASAP7_75t_R _24959_ (.A1(net5696),
    .A2(_02568_),
    .B(_02586_),
    .Y(_02587_));
 AOI21x1_ASAP7_75t_R _24960_ (.A1(net5411),
    .A2(_02392_),
    .B(net5708),
    .Y(_02588_));
 NAND2x1_ASAP7_75t_R _24961_ (.A(net5711),
    .B(net5113),
    .Y(_02589_));
 NAND2x1_ASAP7_75t_R _24962_ (.A(_02589_),
    .B(_02527_),
    .Y(_02590_));
 AOI21x1_ASAP7_75t_R _24963_ (.A1(_02588_),
    .A2(_02590_),
    .B(net5700),
    .Y(_02591_));
 AOI21x1_ASAP7_75t_R _24964_ (.A1(net4564),
    .A2(_02447_),
    .B(net6162),
    .Y(_02592_));
 NAND2x1_ASAP7_75t_R _24965_ (.A(net5113),
    .B(net5413),
    .Y(_02593_));
 AO21x1_ASAP7_75t_R _24966_ (.A1(_02593_),
    .A2(_02562_),
    .B(net5411),
    .Y(_02594_));
 NAND2x1_ASAP7_75t_R _24967_ (.A(_02592_),
    .B(_02594_),
    .Y(_02595_));
 AOI21x1_ASAP7_75t_R _24968_ (.A1(_02591_),
    .A2(_02595_),
    .B(net5698),
    .Y(_02596_));
 AO21x1_ASAP7_75t_R _24969_ (.A1(net4511),
    .A2(net4661),
    .B(net5408),
    .Y(_02597_));
 NAND2x1p5_ASAP7_75t_R _24970_ (.A(_02446_),
    .B(_02480_),
    .Y(_02598_));
 AOI21x1_ASAP7_75t_R _24971_ (.A1(_02597_),
    .A2(_02598_),
    .B(net5708),
    .Y(_02599_));
 NAND2x1_ASAP7_75t_R _24972_ (.A(_01250_),
    .B(net5408),
    .Y(_02600_));
 AO21x1_ASAP7_75t_R _24973_ (.A1(_02448_),
    .A2(net4511),
    .B(net5408),
    .Y(_02601_));
 AOI21x1_ASAP7_75t_R _24974_ (.A1(net4879),
    .A2(_02601_),
    .B(net6162),
    .Y(_02602_));
 OAI21x1_ASAP7_75t_R _24976_ (.A1(_02599_),
    .A2(_02602_),
    .B(net5700),
    .Y(_02604_));
 NAND2x1_ASAP7_75t_R _24977_ (.A(_02596_),
    .B(_02604_),
    .Y(_02605_));
 NAND2x1_ASAP7_75t_R _24978_ (.A(net5113),
    .B(net5412),
    .Y(_02606_));
 INVx2_ASAP7_75t_R _24979_ (.A(_02514_),
    .Y(_02607_));
 NAND2x1p5_ASAP7_75t_R _24980_ (.A(_02606_),
    .B(_02607_),
    .Y(_02608_));
 NAND2x1_ASAP7_75t_R _24981_ (.A(net5711),
    .B(net5415),
    .Y(_02609_));
 AOI21x1_ASAP7_75t_R _24982_ (.A1(_02609_),
    .A2(_02447_),
    .B(net5709),
    .Y(_02610_));
 AOI21x1_ASAP7_75t_R _24983_ (.A1(_02610_),
    .A2(_02608_),
    .B(net5404),
    .Y(_02611_));
 INVx1_ASAP7_75t_R _24984_ (.A(_02489_),
    .Y(_02612_));
 NOR2x1_ASAP7_75t_R _24985_ (.A(_02612_),
    .B(_02497_),
    .Y(_02613_));
 AOI21x1_ASAP7_75t_R _24986_ (.A1(net5415),
    .A2(net5413),
    .B(net5407),
    .Y(_02614_));
 INVx1_ASAP7_75t_R _24987_ (.A(_02474_),
    .Y(_02615_));
 AND2x2_ASAP7_75t_R _24988_ (.A(_02614_),
    .B(_02615_),
    .Y(_02616_));
 OAI21x1_ASAP7_75t_R _24989_ (.A1(_02613_),
    .A2(_02616_),
    .B(net5708),
    .Y(_02617_));
 NAND2x1_ASAP7_75t_R _24990_ (.A(_02617_),
    .B(_02611_),
    .Y(_02618_));
 AOI21x1_ASAP7_75t_R _24991_ (.A1(net5703),
    .A2(net4666),
    .B(net5708),
    .Y(_02619_));
 AOI21x1_ASAP7_75t_R _24992_ (.A1(_02619_),
    .A2(_02551_),
    .B(net5700),
    .Y(_02620_));
 AOI21x1_ASAP7_75t_R _24993_ (.A1(net5058),
    .A2(_02336_),
    .B(net5703),
    .Y(_02621_));
 AOI21x1_ASAP7_75t_R _24994_ (.A1(_02448_),
    .A2(_02621_),
    .B(net6162),
    .Y(_02622_));
 OAI21x1_ASAP7_75t_R _24995_ (.A1(net5411),
    .A2(_02577_),
    .B(_02622_),
    .Y(_02623_));
 AOI21x1_ASAP7_75t_R _24996_ (.A1(_02620_),
    .A2(_02623_),
    .B(net6163),
    .Y(_02624_));
 AOI21x1_ASAP7_75t_R _24997_ (.A1(_02624_),
    .A2(_02618_),
    .B(_02443_),
    .Y(_02625_));
 NAND2x1_ASAP7_75t_R _24998_ (.A(_02625_),
    .B(_02605_),
    .Y(_02626_));
 OAI21x1_ASAP7_75t_R _24999_ (.A1(_02544_),
    .A2(_02587_),
    .B(_02626_),
    .Y(_00097_));
 INVx1_ASAP7_75t_R _25000_ (.A(_02379_),
    .Y(_02627_));
 AO21x1_ASAP7_75t_R _25001_ (.A1(net5412),
    .A2(net4804),
    .B(net5407),
    .Y(_02628_));
 NOR2x1_ASAP7_75t_R _25002_ (.A(_02627_),
    .B(_02628_),
    .Y(_02629_));
 NAND2x1_ASAP7_75t_R _25003_ (.A(net5714),
    .B(net5412),
    .Y(_02630_));
 AND2x2_ASAP7_75t_R _25004_ (.A(_02581_),
    .B(_02630_),
    .Y(_02631_));
 OAI21x1_ASAP7_75t_R _25005_ (.A1(_02629_),
    .A2(_02631_),
    .B(net5709),
    .Y(_02632_));
 NAND2x1_ASAP7_75t_R _25006_ (.A(net5409),
    .B(_02489_),
    .Y(_02633_));
 OA21x2_ASAP7_75t_R _25007_ (.A1(_02633_),
    .A2(net4508),
    .B(net6162),
    .Y(_02634_));
 AOI21x1_ASAP7_75t_R _25008_ (.A1(_02528_),
    .A2(_02634_),
    .B(net5404),
    .Y(_02635_));
 NAND2x1_ASAP7_75t_R _25009_ (.A(_02632_),
    .B(_02635_),
    .Y(_02636_));
 NAND2x1_ASAP7_75t_R _25010_ (.A(net5416),
    .B(net5412),
    .Y(_02637_));
 NAND3x1_ASAP7_75t_R _25011_ (.A(_02637_),
    .B(net5411),
    .C(net4509),
    .Y(_02638_));
 AO21x1_ASAP7_75t_R _25012_ (.A1(_02563_),
    .A2(net4563),
    .B(net5411),
    .Y(_02639_));
 AOI21x1_ASAP7_75t_R _25013_ (.A1(_02638_),
    .A2(_02639_),
    .B(net6162),
    .Y(_02640_));
 AO21x1_ASAP7_75t_R _25014_ (.A1(net5413),
    .A2(_02576_),
    .B(net5706),
    .Y(_02641_));
 NOR2x1_ASAP7_75t_R _25015_ (.A(net4884),
    .B(_02336_),
    .Y(_02642_));
 OA211x2_ASAP7_75t_R _25016_ (.A1(_02641_),
    .A2(_02642_),
    .B(net6162),
    .C(net4446),
    .Y(_02643_));
 OAI21x1_ASAP7_75t_R _25017_ (.A1(_02640_),
    .A2(_02643_),
    .B(net5405),
    .Y(_02644_));
 AOI21x1_ASAP7_75t_R _25018_ (.A1(_02636_),
    .A2(_02644_),
    .B(net5698),
    .Y(_02645_));
 NAND2x1_ASAP7_75t_R _25019_ (.A(_02489_),
    .B(_02495_),
    .Y(_02646_));
 AOI21x1_ASAP7_75t_R _25020_ (.A1(net5704),
    .A2(_02646_),
    .B(net5708),
    .Y(_02647_));
 AO21x1_ASAP7_75t_R _25021_ (.A1(_02630_),
    .A2(net4510),
    .B(net5705),
    .Y(_02648_));
 NAND2x1_ASAP7_75t_R _25022_ (.A(_02647_),
    .B(_02648_),
    .Y(_02649_));
 OA21x2_ASAP7_75t_R _25023_ (.A1(_02495_),
    .A2(net5409),
    .B(net5708),
    .Y(_02650_));
 OAI21x1_ASAP7_75t_R _25024_ (.A1(net5710),
    .A2(net6164),
    .B(_02445_),
    .Y(_02651_));
 NAND2x1_ASAP7_75t_R _25025_ (.A(net5705),
    .B(_02651_),
    .Y(_02652_));
 OAI21x1_ASAP7_75t_R _25026_ (.A1(_02525_),
    .A2(_02633_),
    .B(_02652_),
    .Y(_02653_));
 AOI21x1_ASAP7_75t_R _25027_ (.A1(_02650_),
    .A2(_02653_),
    .B(net5405),
    .Y(_02654_));
 NAND2x1_ASAP7_75t_R _25028_ (.A(_02649_),
    .B(_02654_),
    .Y(_02655_));
 INVx1_ASAP7_75t_R _25029_ (.A(_02651_),
    .Y(_02656_));
 OAI21x1_ASAP7_75t_R _25030_ (.A1(_02656_),
    .A2(_02430_),
    .B(net5708),
    .Y(_02657_));
 INVx1_ASAP7_75t_R _25031_ (.A(_02495_),
    .Y(_02658_));
 AOI211x1_ASAP7_75t_R _25032_ (.A1(net5414),
    .A2(net5711),
    .B(_02658_),
    .C(net5705),
    .Y(_02659_));
 NOR2x1_ASAP7_75t_R _25033_ (.A(_02657_),
    .B(_02659_),
    .Y(_02660_));
 AOI21x1_ASAP7_75t_R _25034_ (.A1(net4561),
    .A2(_02468_),
    .B(net5705),
    .Y(_02661_));
 INVx1_ASAP7_75t_R _25035_ (.A(_02661_),
    .Y(_02662_));
 AOI21x1_ASAP7_75t_R _25036_ (.A1(net5060),
    .A2(net5413),
    .B(net5406),
    .Y(_02663_));
 NAND2x1_ASAP7_75t_R _25037_ (.A(_02606_),
    .B(_02663_),
    .Y(_02664_));
 AOI21x1_ASAP7_75t_R _25038_ (.A1(_02662_),
    .A2(_02664_),
    .B(net5708),
    .Y(_02665_));
 OAI21x1_ASAP7_75t_R _25039_ (.A1(_02660_),
    .A2(_02665_),
    .B(net5405),
    .Y(_02666_));
 NAND2x1_ASAP7_75t_R _25040_ (.A(_02655_),
    .B(_02666_),
    .Y(_02667_));
 OAI21x1_ASAP7_75t_R _25041_ (.A1(net6163),
    .A2(_02667_),
    .B(_02443_),
    .Y(_02668_));
 AND2x2_ASAP7_75t_R _25042_ (.A(_02527_),
    .B(_02422_),
    .Y(_02669_));
 NAND2x1p5_ASAP7_75t_R _25043_ (.A(net5409),
    .B(net4465),
    .Y(_02670_));
 NOR2x1_ASAP7_75t_R _25044_ (.A(_02419_),
    .B(_02670_),
    .Y(_02671_));
 OA21x2_ASAP7_75t_R _25045_ (.A1(_02669_),
    .A2(_02671_),
    .B(net5708),
    .Y(_02672_));
 OAI21x1_ASAP7_75t_R _25046_ (.A1(net5711),
    .A2(net5413),
    .B(net5410),
    .Y(_02673_));
 OAI21x1_ASAP7_75t_R _25047_ (.A1(_02429_),
    .A2(_02673_),
    .B(net6162),
    .Y(_02674_));
 INVx1_ASAP7_75t_R _25048_ (.A(_02674_),
    .Y(_02675_));
 NAND2x1_ASAP7_75t_R _25049_ (.A(_01248_),
    .B(net5703),
    .Y(_02676_));
 AO21x1_ASAP7_75t_R _25050_ (.A1(_02675_),
    .A2(_02676_),
    .B(net5404),
    .Y(_02677_));
 OA21x2_ASAP7_75t_R _25051_ (.A1(net5409),
    .A2(_01246_),
    .B(net6162),
    .Y(_02678_));
 AO21x1_ASAP7_75t_R _25052_ (.A1(net4661),
    .A2(net4465),
    .B(net5704),
    .Y(_02679_));
 AOI21x1_ASAP7_75t_R _25053_ (.A1(_02678_),
    .A2(_02679_),
    .B(net5700),
    .Y(_02680_));
 AOI21x1_ASAP7_75t_R _25054_ (.A1(net4464),
    .A2(_02527_),
    .B(net6162),
    .Y(_02681_));
 AO21x1_ASAP7_75t_R _25055_ (.A1(_02637_),
    .A2(_02563_),
    .B(net5703),
    .Y(_02682_));
 NAND2x1_ASAP7_75t_R _25056_ (.A(_02681_),
    .B(_02682_),
    .Y(_02683_));
 AOI21x1_ASAP7_75t_R _25057_ (.A1(_02680_),
    .A2(_02683_),
    .B(net6163),
    .Y(_02684_));
 OAI21x1_ASAP7_75t_R _25058_ (.A1(_02672_),
    .A2(_02677_),
    .B(_02684_),
    .Y(_02685_));
 OAI21x1_ASAP7_75t_R _25059_ (.A1(_01251_),
    .A2(net5410),
    .B(net5709),
    .Y(_02686_));
 NAND2x1_ASAP7_75t_R _25060_ (.A(net6537),
    .B(_02369_),
    .Y(_02687_));
 INVx1_ASAP7_75t_R _25061_ (.A(net6537),
    .Y(_02688_));
 INVx1_ASAP7_75t_R _25062_ (.A(_02369_),
    .Y(_02689_));
 NAND2x1_ASAP7_75t_R _25063_ (.A(_02688_),
    .B(_02689_),
    .Y(_02690_));
 INVx1_ASAP7_75t_R _25064_ (.A(_01245_),
    .Y(_02691_));
 AOI21x1_ASAP7_75t_R _25065_ (.A1(_02687_),
    .A2(_02690_),
    .B(_02691_),
    .Y(_02692_));
 AOI21x1_ASAP7_75t_R _25066_ (.A1(net5706),
    .A2(net4515),
    .B(_02692_),
    .Y(_02693_));
 AOI21x1_ASAP7_75t_R _25067_ (.A1(net6162),
    .A2(_02693_),
    .B(net5404),
    .Y(_02694_));
 OAI21x1_ASAP7_75t_R _25068_ (.A1(_02686_),
    .A2(_02631_),
    .B(_02694_),
    .Y(_02695_));
 AO21x1_ASAP7_75t_R _25069_ (.A1(net4510),
    .A2(_02468_),
    .B(net5705),
    .Y(_02696_));
 AOI21x1_ASAP7_75t_R _25070_ (.A1(_02475_),
    .A2(_02696_),
    .B(net5700),
    .Y(_02697_));
 AND2x2_ASAP7_75t_R _25071_ (.A(_01233_),
    .B(net4805),
    .Y(_02698_));
 INVx1_ASAP7_75t_R _25072_ (.A(_02698_),
    .Y(_02699_));
 AO21x1_ASAP7_75t_R _25073_ (.A1(_02394_),
    .A2(_02393_),
    .B(_02699_),
    .Y(_02700_));
 INVx1_ASAP7_75t_R _25074_ (.A(_02700_),
    .Y(_02701_));
 AO21x1_ASAP7_75t_R _25075_ (.A1(_02391_),
    .A2(_02390_),
    .B(_01238_),
    .Y(_02702_));
 AOI21x1_ASAP7_75t_R _25076_ (.A1(_02576_),
    .A2(net5412),
    .B(net5407),
    .Y(_02703_));
 AOI21x1_ASAP7_75t_R _25077_ (.A1(_02702_),
    .A2(_02703_),
    .B(net6162),
    .Y(_02704_));
 OAI21x1_ASAP7_75t_R _25078_ (.A1(_02641_),
    .A2(_02701_),
    .B(_02704_),
    .Y(_02705_));
 AOI21x1_ASAP7_75t_R _25079_ (.A1(_02697_),
    .A2(_02705_),
    .B(net5699),
    .Y(_02706_));
 AOI21x1_ASAP7_75t_R _25080_ (.A1(_02695_),
    .A2(_02706_),
    .B(_02443_),
    .Y(_02707_));
 NAND2x1_ASAP7_75t_R _25081_ (.A(_02685_),
    .B(_02707_),
    .Y(_02708_));
 OAI21x1_ASAP7_75t_R _25082_ (.A1(_02645_),
    .A2(_02668_),
    .B(_02708_),
    .Y(_00098_));
 AOI21x1_ASAP7_75t_R _25083_ (.A1(net4560),
    .A2(_02615_),
    .B(net5703),
    .Y(_02709_));
 NOR2x1_ASAP7_75t_R _25084_ (.A(net5113),
    .B(net5412),
    .Y(_02710_));
 OA21x2_ASAP7_75t_R _25085_ (.A1(_02710_),
    .A2(_02419_),
    .B(net5703),
    .Y(_02711_));
 OAI21x1_ASAP7_75t_R _25086_ (.A1(_02709_),
    .A2(_02711_),
    .B(net5708),
    .Y(_02712_));
 OAI21x1_ASAP7_75t_R _25087_ (.A1(_02612_),
    .A2(_02546_),
    .B(net5409),
    .Y(_02713_));
 AO21x1_ASAP7_75t_R _25088_ (.A1(_02639_),
    .A2(_02713_),
    .B(net5708),
    .Y(_02714_));
 AOI21x1_ASAP7_75t_R _25089_ (.A1(_02712_),
    .A2(_02714_),
    .B(net5700),
    .Y(_02715_));
 AO21x1_ASAP7_75t_R _25090_ (.A1(_02637_),
    .A2(_02563_),
    .B(net5411),
    .Y(_02716_));
 NOR2x1_ASAP7_75t_R _25091_ (.A(net6162),
    .B(_02480_),
    .Y(_02717_));
 AO21x1_ASAP7_75t_R _25092_ (.A1(_02716_),
    .A2(_02717_),
    .B(net5405),
    .Y(_02718_));
 OA21x2_ASAP7_75t_R _25093_ (.A1(_02710_),
    .A2(net5112),
    .B(net5703),
    .Y(_02719_));
 AOI21x1_ASAP7_75t_R _25094_ (.A1(net4467),
    .A2(_02563_),
    .B(net5703),
    .Y(_02720_));
 NOR3x1_ASAP7_75t_R _25095_ (.A(_02719_),
    .B(_02720_),
    .C(net5708),
    .Y(_02721_));
 OAI21x1_ASAP7_75t_R _25096_ (.A1(_02718_),
    .A2(_02721_),
    .B(net6163),
    .Y(_02722_));
 OAI21x1_ASAP7_75t_R _25097_ (.A1(_02715_),
    .A2(_02722_),
    .B(_02544_),
    .Y(_02723_));
 OAI21x1_ASAP7_75t_R _25098_ (.A1(net4442),
    .A2(_02719_),
    .B(net6162),
    .Y(_02724_));
 NAND2x1_ASAP7_75t_R _25099_ (.A(net4467),
    .B(_02663_),
    .Y(_02725_));
 NAND2x1_ASAP7_75t_R _25100_ (.A(_02448_),
    .B(_02621_),
    .Y(_02726_));
 AO21x1_ASAP7_75t_R _25101_ (.A1(_02725_),
    .A2(_02726_),
    .B(net6162),
    .Y(_02727_));
 AOI21x1_ASAP7_75t_R _25102_ (.A1(_02724_),
    .A2(_02727_),
    .B(net5405),
    .Y(_02728_));
 AOI21x1_ASAP7_75t_R _25103_ (.A1(_02432_),
    .A2(_02433_),
    .B(net5703),
    .Y(_02729_));
 AOI21x1_ASAP7_75t_R _25104_ (.A1(net4563),
    .A2(_02578_),
    .B(net5411),
    .Y(_02730_));
 OAI21x1_ASAP7_75t_R _25105_ (.A1(_02729_),
    .A2(_02730_),
    .B(net5708),
    .Y(_02731_));
 AOI21x1_ASAP7_75t_R _25106_ (.A1(net4464),
    .A2(_02577_),
    .B(net5411),
    .Y(_02732_));
 INVx1_ASAP7_75t_R _25107_ (.A(_02392_),
    .Y(_02733_));
 AOI21x1_ASAP7_75t_R _25108_ (.A1(_02733_),
    .A2(_02420_),
    .B(net5703),
    .Y(_02734_));
 OAI21x1_ASAP7_75t_R _25109_ (.A1(_02732_),
    .A2(_02734_),
    .B(net6162),
    .Y(_02735_));
 AOI21x1_ASAP7_75t_R _25110_ (.A1(_02731_),
    .A2(_02735_),
    .B(net5700),
    .Y(_02736_));
 NOR3x1_ASAP7_75t_R _25111_ (.A(_02728_),
    .B(net6163),
    .C(_02736_),
    .Y(_02737_));
 OAI21x1_ASAP7_75t_R _25112_ (.A1(net4559),
    .A2(_02574_),
    .B(_02531_),
    .Y(_02738_));
 AO21x1_ASAP7_75t_R _25113_ (.A1(net5414),
    .A2(_02417_),
    .B(net5407),
    .Y(_02739_));
 NAND2x1_ASAP7_75t_R _25114_ (.A(net5700),
    .B(_02630_),
    .Y(_02740_));
 NAND2x1_ASAP7_75t_R _25115_ (.A(net5404),
    .B(_02481_),
    .Y(_02741_));
 OAI21x1_ASAP7_75t_R _25116_ (.A1(_02739_),
    .A2(_02740_),
    .B(_02741_),
    .Y(_02742_));
 OAI21x1_ASAP7_75t_R _25117_ (.A1(_02738_),
    .A2(_02742_),
    .B(net6163),
    .Y(_02743_));
 OA21x2_ASAP7_75t_R _25118_ (.A1(net4663),
    .A2(net5704),
    .B(net5405),
    .Y(_02744_));
 NAND2x1_ASAP7_75t_R _25119_ (.A(_02744_),
    .B(_02664_),
    .Y(_02745_));
 NAND2x1_ASAP7_75t_R _25120_ (.A(_02700_),
    .B(_02621_),
    .Y(_02746_));
 AOI21x1_ASAP7_75t_R _25121_ (.A1(net4565),
    .A2(_02388_),
    .B(net5405),
    .Y(_02747_));
 NAND2x1_ASAP7_75t_R _25122_ (.A(_02746_),
    .B(_02747_),
    .Y(_02748_));
 AOI21x1_ASAP7_75t_R _25123_ (.A1(_02745_),
    .A2(_02748_),
    .B(net5708),
    .Y(_02749_));
 NOR2x1_ASAP7_75t_R _25124_ (.A(_02743_),
    .B(_02749_),
    .Y(_02750_));
 NAND2x1_ASAP7_75t_R _25125_ (.A(net5700),
    .B(_02657_),
    .Y(_02751_));
 OA21x2_ASAP7_75t_R _25126_ (.A1(net6165),
    .A2(net5712),
    .B(_02699_),
    .Y(_02752_));
 OAI21x1_ASAP7_75t_R _25127_ (.A1(net4880),
    .A2(_02752_),
    .B(net5407),
    .Y(_02753_));
 NAND2x1_ASAP7_75t_R _25128_ (.A(_02702_),
    .B(_02703_),
    .Y(_02754_));
 AOI21x1_ASAP7_75t_R _25129_ (.A1(_02753_),
    .A2(_02754_),
    .B(net5708),
    .Y(_02755_));
 OAI21x1_ASAP7_75t_R _25130_ (.A1(_02751_),
    .A2(_02755_),
    .B(_02463_),
    .Y(_02756_));
 AOI21x1_ASAP7_75t_R _25131_ (.A1(_02447_),
    .A2(_02506_),
    .B(net5709),
    .Y(_02757_));
 NAND2x1_ASAP7_75t_R _25132_ (.A(_02590_),
    .B(_02757_),
    .Y(_02758_));
 AO21x1_ASAP7_75t_R _25133_ (.A1(_02651_),
    .A2(_02468_),
    .B(net5407),
    .Y(_02759_));
 AOI21x1_ASAP7_75t_R _25134_ (.A1(net5407),
    .A2(_02658_),
    .B(net6162),
    .Y(_02760_));
 NAND3x1_ASAP7_75t_R _25135_ (.A(net5407),
    .B(net5414),
    .C(net5113),
    .Y(_02761_));
 NAND3x1_ASAP7_75t_R _25136_ (.A(_02759_),
    .B(_02760_),
    .C(_02761_),
    .Y(_02762_));
 AOI21x1_ASAP7_75t_R _25137_ (.A1(_02758_),
    .A2(_02762_),
    .B(net5700),
    .Y(_02763_));
 NOR2x1_ASAP7_75t_R _25138_ (.A(_02756_),
    .B(_02763_),
    .Y(_02764_));
 OAI21x1_ASAP7_75t_R _25139_ (.A1(_02750_),
    .A2(_02764_),
    .B(_02443_),
    .Y(_02765_));
 OAI21x1_ASAP7_75t_R _25140_ (.A1(_02723_),
    .A2(_02737_),
    .B(_02765_),
    .Y(_00099_));
 AO21x1_ASAP7_75t_R _25141_ (.A1(net4809),
    .A2(net5413),
    .B(_02673_),
    .Y(_02766_));
 NAND2x1_ASAP7_75t_R _25142_ (.A(net5714),
    .B(net5416),
    .Y(_02767_));
 AO21x1_ASAP7_75t_R _25143_ (.A1(_02448_),
    .A2(_02767_),
    .B(net5410),
    .Y(_02768_));
 AO21x1_ASAP7_75t_R _25144_ (.A1(_02766_),
    .A2(_02768_),
    .B(net6162),
    .Y(_02769_));
 OA21x2_ASAP7_75t_R _25145_ (.A1(_02674_),
    .A2(_02571_),
    .B(net5701),
    .Y(_02770_));
 AO21x1_ASAP7_75t_R _25146_ (.A1(net5413),
    .A2(net5060),
    .B(net5702),
    .Y(_02771_));
 INVx1_ASAP7_75t_R _25147_ (.A(net4514),
    .Y(_02772_));
 AO21x1_ASAP7_75t_R _25148_ (.A1(_02771_),
    .A2(_02772_),
    .B(net6162),
    .Y(_02773_));
 NOR2x1_ASAP7_75t_R _25149_ (.A(_02375_),
    .B(_02582_),
    .Y(_02774_));
 NAND2x1_ASAP7_75t_R _25150_ (.A(net5711),
    .B(net5413),
    .Y(_02775_));
 AOI21x1_ASAP7_75t_R _25151_ (.A1(_02775_),
    .A2(_02637_),
    .B(net5703),
    .Y(_02776_));
 OAI21x1_ASAP7_75t_R _25152_ (.A1(_02774_),
    .A2(_02776_),
    .B(net6162),
    .Y(_02777_));
 AOI21x1_ASAP7_75t_R _25153_ (.A1(_02773_),
    .A2(_02777_),
    .B(net5701),
    .Y(_02778_));
 AOI211x1_ASAP7_75t_R _25154_ (.A1(_02769_),
    .A2(_02770_),
    .B(_02778_),
    .C(net6163),
    .Y(_02779_));
 AO21x1_ASAP7_75t_R _25155_ (.A1(_02563_),
    .A2(_02615_),
    .B(net5703),
    .Y(_02780_));
 AND2x2_ASAP7_75t_R _25156_ (.A(_02780_),
    .B(_02504_),
    .Y(_02781_));
 OAI21x1_ASAP7_75t_R _25157_ (.A1(_02627_),
    .A2(_02628_),
    .B(net5709),
    .Y(_02782_));
 AO21x1_ASAP7_75t_R _25158_ (.A1(_02394_),
    .A2(_02393_),
    .B(net4806),
    .Y(_02783_));
 AND3x1_ASAP7_75t_R _25159_ (.A(_02775_),
    .B(_02783_),
    .C(net5411),
    .Y(_02784_));
 OAI21x1_ASAP7_75t_R _25160_ (.A1(_02782_),
    .A2(_02784_),
    .B(net5701),
    .Y(_02785_));
 INVx2_ASAP7_75t_R _25161_ (.A(_02513_),
    .Y(_02786_));
 OAI21x1_ASAP7_75t_R _25162_ (.A1(_02786_),
    .A2(_02546_),
    .B(net5704),
    .Y(_02787_));
 AOI21x1_ASAP7_75t_R _25163_ (.A1(_02538_),
    .A2(_02787_),
    .B(net5708),
    .Y(_02788_));
 AO21x1_ASAP7_75t_R _25164_ (.A1(net4511),
    .A2(net4663),
    .B(net5409),
    .Y(_02789_));
 AO21x1_ASAP7_75t_R _25165_ (.A1(net4663),
    .A2(net4465),
    .B(net5704),
    .Y(_02790_));
 AOI21x1_ASAP7_75t_R _25166_ (.A1(_02789_),
    .A2(_02790_),
    .B(net6162),
    .Y(_02791_));
 OAI21x1_ASAP7_75t_R _25167_ (.A1(_02788_),
    .A2(_02791_),
    .B(net5404),
    .Y(_02792_));
 OAI21x1_ASAP7_75t_R _25168_ (.A1(_02781_),
    .A2(_02785_),
    .B(_02792_),
    .Y(_02793_));
 OAI21x1_ASAP7_75t_R _25169_ (.A1(net5696),
    .A2(_02793_),
    .B(_02544_),
    .Y(_02794_));
 AO21x1_ASAP7_75t_R _25170_ (.A1(_02637_),
    .A2(_02589_),
    .B(net5703),
    .Y(_02795_));
 AO21x1_ASAP7_75t_R _25171_ (.A1(_02795_),
    .A2(net4444),
    .B(net5709),
    .Y(_02796_));
 INVx1_ASAP7_75t_R _25172_ (.A(_02536_),
    .Y(_02797_));
 AO21x1_ASAP7_75t_R _25173_ (.A1(_02606_),
    .A2(_02797_),
    .B(net5702),
    .Y(_02798_));
 AO21x1_ASAP7_75t_R _25174_ (.A1(_02798_),
    .A2(_02768_),
    .B(net6162),
    .Y(_02799_));
 AOI21x1_ASAP7_75t_R _25175_ (.A1(_02796_),
    .A2(_02799_),
    .B(net5697),
    .Y(_02800_));
 AO21x1_ASAP7_75t_R _25176_ (.A1(_02606_),
    .A2(net4660),
    .B(net5407),
    .Y(_02801_));
 NAND2x1_ASAP7_75t_R _25177_ (.A(net5413),
    .B(net5406),
    .Y(_02802_));
 AND2x2_ASAP7_75t_R _25178_ (.A(_02802_),
    .B(net6162),
    .Y(_02803_));
 AO21x1_ASAP7_75t_R _25179_ (.A1(_02801_),
    .A2(_02803_),
    .B(net6163),
    .Y(_02804_));
 AO21x1_ASAP7_75t_R _25180_ (.A1(_02775_),
    .A2(_02615_),
    .B(_02376_),
    .Y(_02805_));
 AND2x2_ASAP7_75t_R _25181_ (.A(_02569_),
    .B(_02805_),
    .Y(_02806_));
 OAI21x1_ASAP7_75t_R _25182_ (.A1(_02804_),
    .A2(_02806_),
    .B(net5701),
    .Y(_02807_));
 OA21x2_ASAP7_75t_R _25183_ (.A1(net5407),
    .A2(_02576_),
    .B(net6162),
    .Y(_02808_));
 AOI21x1_ASAP7_75t_R _25184_ (.A1(_02670_),
    .A2(_02808_),
    .B(_02463_),
    .Y(_02809_));
 NOR2x1_ASAP7_75t_R _25185_ (.A(net5713),
    .B(net5414),
    .Y(_02810_));
 OA21x2_ASAP7_75t_R _25186_ (.A1(_02502_),
    .A2(net5407),
    .B(net5709),
    .Y(_02811_));
 OAI21x1_ASAP7_75t_R _25187_ (.A1(_02810_),
    .A2(_02771_),
    .B(_02811_),
    .Y(_02812_));
 AOI21x1_ASAP7_75t_R _25188_ (.A1(_02809_),
    .A2(_02812_),
    .B(net5700),
    .Y(_02813_));
 NOR2x1_ASAP7_75t_R _25189_ (.A(_02786_),
    .B(_02628_),
    .Y(_02814_));
 AO21x1_ASAP7_75t_R _25190_ (.A1(net5413),
    .A2(net4807),
    .B(net5406),
    .Y(_02815_));
 AOI21x1_ASAP7_75t_R _25191_ (.A1(net5406),
    .A2(_02426_),
    .B(net6162),
    .Y(_02816_));
 AOI21x1_ASAP7_75t_R _25192_ (.A1(_02815_),
    .A2(_02816_),
    .B(net6163),
    .Y(_02817_));
 OAI21x1_ASAP7_75t_R _25193_ (.A1(_02491_),
    .A2(_02814_),
    .B(_02817_),
    .Y(_02818_));
 AOI21x1_ASAP7_75t_R _25194_ (.A1(_02813_),
    .A2(_02818_),
    .B(_02544_),
    .Y(_02819_));
 OAI21x1_ASAP7_75t_R _25195_ (.A1(_02800_),
    .A2(_02807_),
    .B(_02819_),
    .Y(_02820_));
 OAI21x1_ASAP7_75t_R _25196_ (.A1(_02779_),
    .A2(_02794_),
    .B(_02820_),
    .Y(_00100_));
 INVx1_ASAP7_75t_R _25197_ (.A(_02630_),
    .Y(_02821_));
 OAI22x1_ASAP7_75t_R _25198_ (.A1(_02815_),
    .A2(_02821_),
    .B1(net4722),
    .B2(_02802_),
    .Y(_02822_));
 AO21x1_ASAP7_75t_R _25199_ (.A1(net4660),
    .A2(net5702),
    .B(net5709),
    .Y(_02823_));
 NOR2x1p5_ASAP7_75t_R _25200_ (.A(_02521_),
    .B(_02497_),
    .Y(_02824_));
 OAI21x1_ASAP7_75t_R _25201_ (.A1(_02823_),
    .A2(_02824_),
    .B(net5700),
    .Y(_02825_));
 AO21x1_ASAP7_75t_R _25202_ (.A1(_02822_),
    .A2(net5709),
    .B(_02825_),
    .Y(_02826_));
 OA21x2_ASAP7_75t_R _25203_ (.A1(net5706),
    .A2(net5714),
    .B(net6162),
    .Y(_02827_));
 AOI21x1_ASAP7_75t_R _25204_ (.A1(_02827_),
    .A2(_02768_),
    .B(net5701),
    .Y(_02828_));
 AO21x1_ASAP7_75t_R _25205_ (.A1(_02578_),
    .A2(_02577_),
    .B(net5703),
    .Y(_02829_));
 AO21x1_ASAP7_75t_R _25206_ (.A1(_02593_),
    .A2(_02767_),
    .B(net5410),
    .Y(_02830_));
 AO21x1_ASAP7_75t_R _25207_ (.A1(_02829_),
    .A2(_02830_),
    .B(net6162),
    .Y(_02831_));
 NAND2x1_ASAP7_75t_R _25208_ (.A(_02828_),
    .B(_02831_),
    .Y(_02832_));
 AOI21x1_ASAP7_75t_R _25209_ (.A1(_02832_),
    .A2(_02826_),
    .B(net5697),
    .Y(_02833_));
 NOR2x1_ASAP7_75t_R _25210_ (.A(net6162),
    .B(_02392_),
    .Y(_02834_));
 AO21x1_ASAP7_75t_R _25211_ (.A1(_02628_),
    .A2(_02834_),
    .B(net5404),
    .Y(_02835_));
 AOI21x1_ASAP7_75t_R _25212_ (.A1(net4662),
    .A2(_02593_),
    .B(net5702),
    .Y(_02836_));
 NOR3x1_ASAP7_75t_R _25213_ (.A(_02836_),
    .B(net5709),
    .C(_02427_),
    .Y(_02837_));
 OAI21x1_ASAP7_75t_R _25214_ (.A1(_02835_),
    .A2(_02837_),
    .B(net5697),
    .Y(_02838_));
 AO21x1_ASAP7_75t_R _25215_ (.A1(net5412),
    .A2(_02458_),
    .B(net4664),
    .Y(_02839_));
 AOI221x1_ASAP7_75t_R _25216_ (.A1(net4659),
    .A2(_02663_),
    .B1(net5407),
    .B2(_02839_),
    .C(net6162),
    .Y(_02840_));
 OA21x2_ASAP7_75t_R _25217_ (.A1(_02656_),
    .A2(net4666),
    .B(net5409),
    .Y(_02841_));
 OAI21x1_ASAP7_75t_R _25218_ (.A1(_02841_),
    .A2(_02462_),
    .B(net5404),
    .Y(_02842_));
 NOR2x1_ASAP7_75t_R _25219_ (.A(_02840_),
    .B(_02842_),
    .Y(_02843_));
 OAI21x1_ASAP7_75t_R _25220_ (.A1(_02838_),
    .A2(_02843_),
    .B(_02544_),
    .Y(_02844_));
 AND2x2_ASAP7_75t_R _25221_ (.A(_02663_),
    .B(_02448_),
    .Y(_02845_));
 AOI21x1_ASAP7_75t_R _25222_ (.A1(net4563),
    .A2(net4442),
    .B(_02845_),
    .Y(_02846_));
 OAI22x1_ASAP7_75t_R _25223_ (.A1(net4885),
    .A2(net5112),
    .B1(net5113),
    .B2(net5703),
    .Y(_02847_));
 OAI21x1_ASAP7_75t_R _25224_ (.A1(net5707),
    .A2(_02847_),
    .B(net5404),
    .Y(_02848_));
 AOI21x1_ASAP7_75t_R _25225_ (.A1(net5707),
    .A2(_02846_),
    .B(_02848_),
    .Y(_02849_));
 OA21x2_ASAP7_75t_R _25226_ (.A1(_02525_),
    .A2(_02612_),
    .B(net5704),
    .Y(_02850_));
 NOR2x1_ASAP7_75t_R _25227_ (.A(_02850_),
    .B(_02491_),
    .Y(_02851_));
 OA21x2_ASAP7_75t_R _25228_ (.A1(_02578_),
    .A2(net5703),
    .B(net5709),
    .Y(_02852_));
 NAND2x1_ASAP7_75t_R _25229_ (.A(_02379_),
    .B(_02703_),
    .Y(_02853_));
 AO21x1_ASAP7_75t_R _25230_ (.A1(_02852_),
    .A2(_02853_),
    .B(net5404),
    .Y(_02854_));
 OAI21x1_ASAP7_75t_R _25231_ (.A1(_02851_),
    .A2(_02854_),
    .B(net5699),
    .Y(_02855_));
 INVx1_ASAP7_75t_R _25232_ (.A(_02702_),
    .Y(_02856_));
 AO21x1_ASAP7_75t_R _25233_ (.A1(net4565),
    .A2(net4660),
    .B(net5407),
    .Y(_02857_));
 OAI21x1_ASAP7_75t_R _25234_ (.A1(_02497_),
    .A2(_02856_),
    .B(_02857_),
    .Y(_02858_));
 NOR2x1_ASAP7_75t_R _25235_ (.A(_02417_),
    .B(net5705),
    .Y(_02859_));
 AOI21x1_ASAP7_75t_R _25236_ (.A1(net5705),
    .A2(net4883),
    .B(_02859_),
    .Y(_02860_));
 AOI21x1_ASAP7_75t_R _25237_ (.A1(net6162),
    .A2(_02860_),
    .B(net5404),
    .Y(_02861_));
 OAI21x1_ASAP7_75t_R _25238_ (.A1(net6162),
    .A2(_02858_),
    .B(_02861_),
    .Y(_02862_));
 AOI21x1_ASAP7_75t_R _25239_ (.A1(net5408),
    .A2(_02700_),
    .B(net5709),
    .Y(_02863_));
 OAI21x1_ASAP7_75t_R _25240_ (.A1(_02555_),
    .A2(net4446),
    .B(_02863_),
    .Y(_02864_));
 AOI21x1_ASAP7_75t_R _25241_ (.A1(_02380_),
    .A2(_02499_),
    .B(net5700),
    .Y(_02865_));
 AOI21x1_ASAP7_75t_R _25242_ (.A1(_02864_),
    .A2(_02865_),
    .B(_02463_),
    .Y(_02866_));
 AOI21x1_ASAP7_75t_R _25243_ (.A1(_02862_),
    .A2(_02866_),
    .B(_02544_),
    .Y(_02867_));
 OAI21x1_ASAP7_75t_R _25244_ (.A1(_02849_),
    .A2(_02855_),
    .B(_02867_),
    .Y(_02868_));
 OAI21x1_ASAP7_75t_R _25245_ (.A1(_02844_),
    .A2(_02833_),
    .B(_02868_),
    .Y(_00101_));
 NOR2x1_ASAP7_75t_R _25246_ (.A(net5711),
    .B(net5114),
    .Y(_02869_));
 OAI21x1_ASAP7_75t_R _25247_ (.A1(_02869_),
    .A2(_02810_),
    .B(net5406),
    .Y(_02870_));
 NAND2x1_ASAP7_75t_R _25248_ (.A(_01243_),
    .B(_01249_),
    .Y(_02871_));
 AOI21x1_ASAP7_75t_R _25249_ (.A1(net5702),
    .A2(_02871_),
    .B(net5709),
    .Y(_02872_));
 AND2x2_ASAP7_75t_R _25250_ (.A(_02870_),
    .B(_02872_),
    .Y(_02873_));
 INVx1_ASAP7_75t_R _25251_ (.A(_02760_),
    .Y(_02874_));
 NAND2x1_ASAP7_75t_R _25252_ (.A(net5702),
    .B(net4512),
    .Y(_02875_));
 OAI21x1_ASAP7_75t_R _25253_ (.A1(net4808),
    .A2(_02802_),
    .B(_02875_),
    .Y(_02876_));
 OAI21x1_ASAP7_75t_R _25254_ (.A1(_02874_),
    .A2(_02876_),
    .B(net5404),
    .Y(_02877_));
 OAI21x1_ASAP7_75t_R _25255_ (.A1(_02873_),
    .A2(_02877_),
    .B(net5699),
    .Y(_02878_));
 AO21x1_ASAP7_75t_R _25256_ (.A1(_02391_),
    .A2(_02390_),
    .B(_02698_),
    .Y(_02879_));
 AOI21x1_ASAP7_75t_R _25257_ (.A1(net4662),
    .A2(_02879_),
    .B(net5702),
    .Y(_02880_));
 NOR2x1_ASAP7_75t_R _25258_ (.A(_02525_),
    .B(net4433),
    .Y(_02881_));
 OAI21x1_ASAP7_75t_R _25259_ (.A1(_02880_),
    .A2(_02881_),
    .B(net5709),
    .Y(_02882_));
 OA21x2_ASAP7_75t_R _25260_ (.A1(net4513),
    .A2(_02550_),
    .B(net5407),
    .Y(_02883_));
 AND2x2_ASAP7_75t_R _25261_ (.A(_02663_),
    .B(_02446_),
    .Y(_02884_));
 OAI21x1_ASAP7_75t_R _25262_ (.A1(_02883_),
    .A2(_02884_),
    .B(net6162),
    .Y(_02885_));
 AOI21x1_ASAP7_75t_R _25263_ (.A1(_02882_),
    .A2(_02885_),
    .B(net5404),
    .Y(_02886_));
 OAI21x1_ASAP7_75t_R _25264_ (.A1(_02878_),
    .A2(_02886_),
    .B(_02544_),
    .Y(_02887_));
 AND3x1_ASAP7_75t_R _25265_ (.A(_02433_),
    .B(_02783_),
    .C(net5410),
    .Y(_02888_));
 AO21x1_ASAP7_75t_R _25266_ (.A1(_02607_),
    .A2(_02700_),
    .B(net5404),
    .Y(_02889_));
 NOR2x1_ASAP7_75t_R _25267_ (.A(_02888_),
    .B(_02889_),
    .Y(_02890_));
 AND2x2_ASAP7_75t_R _25268_ (.A(_02581_),
    .B(_02448_),
    .Y(_02891_));
 INVx1_ASAP7_75t_R _25269_ (.A(_02468_),
    .Y(_02892_));
 OAI21x1_ASAP7_75t_R _25270_ (.A1(_02892_),
    .A2(_02815_),
    .B(net5404),
    .Y(_02893_));
 OAI21x1_ASAP7_75t_R _25271_ (.A1(_02891_),
    .A2(_02893_),
    .B(net6162),
    .Y(_02894_));
 NOR2x1_ASAP7_75t_R _25272_ (.A(_02894_),
    .B(_02890_),
    .Y(_02895_));
 INVx1_ASAP7_75t_R _25273_ (.A(_02783_),
    .Y(_02896_));
 AO21x1_ASAP7_75t_R _25274_ (.A1(net5413),
    .A2(net5714),
    .B(net5706),
    .Y(_02897_));
 OAI21x1_ASAP7_75t_R _25275_ (.A1(_02896_),
    .A2(_02897_),
    .B(_02472_),
    .Y(_02898_));
 OAI21x1_ASAP7_75t_R _25276_ (.A1(net5410),
    .A2(net4563),
    .B(net5404),
    .Y(_02899_));
 NOR2x1_ASAP7_75t_R _25277_ (.A(_02899_),
    .B(_02693_),
    .Y(_02900_));
 AOI21x1_ASAP7_75t_R _25278_ (.A1(net5701),
    .A2(_02898_),
    .B(_02900_),
    .Y(_02901_));
 OAI21x1_ASAP7_75t_R _25279_ (.A1(net6162),
    .A2(_02901_),
    .B(net6163),
    .Y(_02902_));
 NOR2x1_ASAP7_75t_R _25280_ (.A(_02902_),
    .B(_02895_),
    .Y(_02903_));
 AO21x1_ASAP7_75t_R _25281_ (.A1(_02433_),
    .A2(_02589_),
    .B(net5703),
    .Y(_02904_));
 OA21x2_ASAP7_75t_R _25282_ (.A1(_02821_),
    .A2(net4446),
    .B(net5404),
    .Y(_02905_));
 AO21x1_ASAP7_75t_R _25283_ (.A1(_02892_),
    .A2(net5702),
    .B(net5404),
    .Y(_02906_));
 OAI21x1_ASAP7_75t_R _25284_ (.A1(_02836_),
    .A2(_02906_),
    .B(net6162),
    .Y(_02907_));
 AOI21x1_ASAP7_75t_R _25285_ (.A1(_02904_),
    .A2(_02905_),
    .B(_02907_),
    .Y(_02908_));
 OA21x2_ASAP7_75t_R _25286_ (.A1(net5413),
    .A2(net4884),
    .B(net5703),
    .Y(_02909_));
 AOI21x1_ASAP7_75t_R _25287_ (.A1(_02432_),
    .A2(_02637_),
    .B(net5703),
    .Y(_02910_));
 AOI211x1_ASAP7_75t_R _25288_ (.A1(net4658),
    .A2(_02433_),
    .B(_02910_),
    .C(net5701),
    .Y(_02911_));
 NAND2x1_ASAP7_75t_R _25289_ (.A(_02606_),
    .B(_02449_),
    .Y(_02912_));
 AND2x2_ASAP7_75t_R _25290_ (.A(_02600_),
    .B(net5700),
    .Y(_02913_));
 AO21x1_ASAP7_75t_R _25291_ (.A1(_02912_),
    .A2(_02913_),
    .B(net6162),
    .Y(_02914_));
 OAI21x1_ASAP7_75t_R _25292_ (.A1(_02911_),
    .A2(_02914_),
    .B(net5697),
    .Y(_02915_));
 NOR2x1_ASAP7_75t_R _25293_ (.A(_02908_),
    .B(_02915_),
    .Y(_02916_));
 AND3x1_ASAP7_75t_R _25294_ (.A(net4467),
    .B(_02379_),
    .C(net5411),
    .Y(_02917_));
 OAI21x1_ASAP7_75t_R _25295_ (.A1(_02559_),
    .A2(_02917_),
    .B(net5404),
    .Y(_02918_));
 AO21x1_ASAP7_75t_R _25296_ (.A1(net5410),
    .A2(_01244_),
    .B(net5709),
    .Y(_02919_));
 NOR2x1_ASAP7_75t_R _25297_ (.A(_02919_),
    .B(_02845_),
    .Y(_02920_));
 OAI21x1_ASAP7_75t_R _25298_ (.A1(_02918_),
    .A2(_02920_),
    .B(net6163),
    .Y(_02921_));
 INVx1_ASAP7_75t_R _25299_ (.A(_02634_),
    .Y(_02922_));
 OAI21x1_ASAP7_75t_R _25300_ (.A1(_02810_),
    .A2(_02771_),
    .B(_02739_),
    .Y(_02923_));
 NAND2x1_ASAP7_75t_R _25301_ (.A(net5709),
    .B(_02923_),
    .Y(_02924_));
 AOI21x1_ASAP7_75t_R _25302_ (.A1(_02922_),
    .A2(_02924_),
    .B(net5404),
    .Y(_02925_));
 OAI21x1_ASAP7_75t_R _25303_ (.A1(_02921_),
    .A2(_02925_),
    .B(_02443_),
    .Y(_02926_));
 OAI22x1_ASAP7_75t_R _25304_ (.A1(_02903_),
    .A2(_02887_),
    .B1(_02916_),
    .B2(_02926_),
    .Y(_00102_));
 OAI21x1_ASAP7_75t_R _25305_ (.A1(net4468),
    .A2(_02389_),
    .B(_02598_),
    .Y(_02927_));
 AOI21x1_ASAP7_75t_R _25306_ (.A1(_02446_),
    .A2(_02663_),
    .B(net5709),
    .Y(_02928_));
 AOI21x1_ASAP7_75t_R _25307_ (.A1(_02928_),
    .A2(_02682_),
    .B(net5405),
    .Y(_02929_));
 OAI21x1_ASAP7_75t_R _25308_ (.A1(_02927_),
    .A2(net6162),
    .B(_02929_),
    .Y(_02930_));
 AOI21x1_ASAP7_75t_R _25309_ (.A1(_02783_),
    .A2(_02388_),
    .B(net6162),
    .Y(_02931_));
 OAI21x1_ASAP7_75t_R _25310_ (.A1(_02505_),
    .A2(_02641_),
    .B(_02931_),
    .Y(_02932_));
 AO21x1_ASAP7_75t_R _25311_ (.A1(_02630_),
    .A2(_02797_),
    .B(net5702),
    .Y(_02933_));
 NOR2x1_ASAP7_75t_R _25312_ (.A(net5709),
    .B(_02909_),
    .Y(_02934_));
 AOI21x1_ASAP7_75t_R _25313_ (.A1(_02933_),
    .A2(_02934_),
    .B(net5701),
    .Y(_02935_));
 AOI21x1_ASAP7_75t_R _25314_ (.A1(_02932_),
    .A2(_02935_),
    .B(net6163),
    .Y(_02936_));
 NAND2x1_ASAP7_75t_R _25315_ (.A(_02936_),
    .B(_02930_),
    .Y(_02937_));
 NOR2x1_ASAP7_75t_R _25316_ (.A(_02576_),
    .B(net5703),
    .Y(_02938_));
 NAND2x1_ASAP7_75t_R _25317_ (.A(net5412),
    .B(_02938_),
    .Y(_02939_));
 NOR2x1_ASAP7_75t_R _25318_ (.A(net5709),
    .B(_02481_),
    .Y(_02940_));
 AOI21x1_ASAP7_75t_R _25319_ (.A1(_02939_),
    .A2(_02940_),
    .B(net5404),
    .Y(_02941_));
 AOI21x1_ASAP7_75t_R _25320_ (.A1(net5411),
    .A2(_02783_),
    .B(net6162),
    .Y(_02942_));
 INVx1_ASAP7_75t_R _25321_ (.A(_02550_),
    .Y(_02943_));
 AO21x1_ASAP7_75t_R _25322_ (.A1(_02943_),
    .A2(net4563),
    .B(net5411),
    .Y(_02944_));
 NAND2x1_ASAP7_75t_R _25323_ (.A(_02942_),
    .B(_02944_),
    .Y(_02945_));
 AOI21x1_ASAP7_75t_R _25324_ (.A1(_02941_),
    .A2(_02945_),
    .B(net5697),
    .Y(_02946_));
 AO21x1_ASAP7_75t_R _25325_ (.A1(_02943_),
    .A2(_02630_),
    .B(net5411),
    .Y(_02947_));
 NAND2x1_ASAP7_75t_R _25326_ (.A(_02675_),
    .B(_02947_),
    .Y(_02948_));
 NAND2x1_ASAP7_75t_R _25327_ (.A(net5706),
    .B(net5113),
    .Y(_02949_));
 OAI21x1_ASAP7_75t_R _25328_ (.A1(_02375_),
    .A2(_02897_),
    .B(_02949_),
    .Y(_02950_));
 AOI21x1_ASAP7_75t_R _25329_ (.A1(net5709),
    .A2(_02950_),
    .B(net5701),
    .Y(_02951_));
 NAND2x1_ASAP7_75t_R _25330_ (.A(_02948_),
    .B(_02951_),
    .Y(_02952_));
 AOI21x1_ASAP7_75t_R _25331_ (.A1(_02946_),
    .A2(_02952_),
    .B(_02544_),
    .Y(_02953_));
 NAND2x1_ASAP7_75t_R _25332_ (.A(_02953_),
    .B(_02937_),
    .Y(_02954_));
 OAI21x1_ASAP7_75t_R _25333_ (.A1(net4512),
    .A2(_02550_),
    .B(net5702),
    .Y(_02955_));
 OAI21x1_ASAP7_75t_R _25334_ (.A1(_02382_),
    .A2(net4881),
    .B(net5407),
    .Y(_02956_));
 AOI21x1_ASAP7_75t_R _25335_ (.A1(_02955_),
    .A2(_02956_),
    .B(net5709),
    .Y(_02957_));
 OAI21x1_ASAP7_75t_R _25336_ (.A1(_02550_),
    .A2(_02810_),
    .B(net5702),
    .Y(_02958_));
 AOI21x1_ASAP7_75t_R _25337_ (.A1(_02753_),
    .A2(_02958_),
    .B(net6162),
    .Y(_02959_));
 OAI21x1_ASAP7_75t_R _25338_ (.A1(_02957_),
    .A2(_02959_),
    .B(net5404),
    .Y(_02960_));
 NAND2x1_ASAP7_75t_R _25339_ (.A(net4664),
    .B(net5702),
    .Y(_02961_));
 AOI21x1_ASAP7_75t_R _25340_ (.A1(_02961_),
    .A2(_02870_),
    .B(net6162),
    .Y(_02962_));
 OAI21x1_ASAP7_75t_R _25341_ (.A1(net4512),
    .A2(_02547_),
    .B(net5705),
    .Y(_02963_));
 OAI21x1_ASAP7_75t_R _25342_ (.A1(net4512),
    .A2(_02455_),
    .B(net5407),
    .Y(_02964_));
 AOI21x1_ASAP7_75t_R _25343_ (.A1(_02963_),
    .A2(_02964_),
    .B(net5708),
    .Y(_02965_));
 OAI21x1_ASAP7_75t_R _25344_ (.A1(_02962_),
    .A2(_02965_),
    .B(net5700),
    .Y(_02966_));
 AOI21x1_ASAP7_75t_R _25345_ (.A1(_02960_),
    .A2(_02966_),
    .B(net6163),
    .Y(_02967_));
 OA21x2_ASAP7_75t_R _25346_ (.A1(_02508_),
    .A2(_02938_),
    .B(net6162),
    .Y(_02968_));
 OAI21x1_ASAP7_75t_R _25347_ (.A1(_02532_),
    .A2(_02455_),
    .B(net5705),
    .Y(_02969_));
 OAI21x1_ASAP7_75t_R _25348_ (.A1(net4666),
    .A2(_02570_),
    .B(net5409),
    .Y(_02970_));
 AOI21x1_ASAP7_75t_R _25349_ (.A1(_02969_),
    .A2(_02970_),
    .B(net6162),
    .Y(_02971_));
 OAI21x1_ASAP7_75t_R _25350_ (.A1(_02968_),
    .A2(_02971_),
    .B(net5404),
    .Y(_02972_));
 AO21x1_ASAP7_75t_R _25351_ (.A1(_02690_),
    .A2(_02687_),
    .B(_01249_),
    .Y(_02973_));
 AO21x1_ASAP7_75t_R _25352_ (.A1(_02495_),
    .A2(net4561),
    .B(net5406),
    .Y(_02974_));
 AOI21x1_ASAP7_75t_R _25353_ (.A1(_02973_),
    .A2(_02974_),
    .B(net5709),
    .Y(_02975_));
 AOI211x1_ASAP7_75t_R _25354_ (.A1(_02614_),
    .A2(_02630_),
    .B(_02661_),
    .C(net6162),
    .Y(_02976_));
 OAI21x1_ASAP7_75t_R _25355_ (.A1(_02975_),
    .A2(_02976_),
    .B(net5700),
    .Y(_02977_));
 AOI21x1_ASAP7_75t_R _25356_ (.A1(_02972_),
    .A2(_02977_),
    .B(net5699),
    .Y(_02978_));
 OAI21x1_ASAP7_75t_R _25357_ (.A1(_02967_),
    .A2(_02978_),
    .B(_02544_),
    .Y(_02979_));
 NAND2x1_ASAP7_75t_R _25358_ (.A(_02979_),
    .B(_02954_),
    .Y(_00103_));
 NOR2x1_ASAP7_75t_R _25359_ (.A(net6668),
    .B(_00471_),
    .Y(_02980_));
 XOR2x2_ASAP7_75t_R _25360_ (.A(_00686_),
    .B(_00679_),
    .Y(_02981_));
 INVx1_ASAP7_75t_R _25361_ (.A(net6558),
    .Y(_02982_));
 XOR2x2_ASAP7_75t_R _25362_ (.A(_02982_),
    .B(_02981_),
    .Y(_02983_));
 XOR2x2_ASAP7_75t_R _25363_ (.A(_14217_),
    .B(_11430_),
    .Y(_02984_));
 NAND2x1p5_ASAP7_75t_R _25364_ (.A(_02984_),
    .B(_02983_),
    .Y(_02985_));
 XOR2x2_ASAP7_75t_R _25365_ (.A(net6558),
    .B(_02981_),
    .Y(_02986_));
 XOR2x2_ASAP7_75t_R _25366_ (.A(_11428_),
    .B(_14217_),
    .Y(_02987_));
 NAND2x1p5_ASAP7_75t_R _25367_ (.A(_02987_),
    .B(_02986_),
    .Y(_02988_));
 AOI21x1_ASAP7_75t_R _25368_ (.A1(_02988_),
    .A2(_02985_),
    .B(net6463),
    .Y(_02989_));
 OAI21x1_ASAP7_75t_R _25369_ (.A1(_02989_),
    .A2(_02980_),
    .B(net6493),
    .Y(_02990_));
 AND2x2_ASAP7_75t_R _25370_ (.A(net6464),
    .B(_00471_),
    .Y(_02991_));
 NAND2x1p5_ASAP7_75t_R _25371_ (.A(_02984_),
    .B(_02986_),
    .Y(_02992_));
 NAND2x1p5_ASAP7_75t_R _25372_ (.A(_02987_),
    .B(_02983_),
    .Y(_02993_));
 AOI21x1_ASAP7_75t_R _25373_ (.A1(_02993_),
    .A2(_02992_),
    .B(net6463),
    .Y(_02994_));
 OAI21x1_ASAP7_75t_R _25374_ (.A1(_02994_),
    .A2(_02991_),
    .B(_08746_),
    .Y(_02995_));
 NAND2x2_ASAP7_75t_R _25375_ (.A(net6161),
    .B(net6160),
    .Y(_01260_));
 NOR2x1_ASAP7_75t_R _25376_ (.A(net6673),
    .B(_00472_),
    .Y(_02996_));
 INVx1_ASAP7_75t_R _25377_ (.A(net6587),
    .Y(_02997_));
 XOR2x2_ASAP7_75t_R _25378_ (.A(_00583_),
    .B(_00615_),
    .Y(_02998_));
 NAND2x1_ASAP7_75t_R _25379_ (.A(_02997_),
    .B(_02998_),
    .Y(_02999_));
 OR2x2_ASAP7_75t_R _25380_ (.A(_02997_),
    .B(_02998_),
    .Y(_03000_));
 INVx1_ASAP7_75t_R _25381_ (.A(net6401),
    .Y(_03001_));
 AOI21x1_ASAP7_75t_R _25382_ (.A1(_02999_),
    .A2(_03000_),
    .B(_03001_),
    .Y(_03002_));
 XOR2x2_ASAP7_75t_R _25383_ (.A(_02998_),
    .B(net6587),
    .Y(_03003_));
 NOR2x1_ASAP7_75t_R _25384_ (.A(net6401),
    .B(_03003_),
    .Y(_03004_));
 OAI21x1_ASAP7_75t_R _25385_ (.A1(_03002_),
    .A2(_03004_),
    .B(net6669),
    .Y(_03005_));
 INVx1_ASAP7_75t_R _25386_ (.A(_03005_),
    .Y(_03006_));
 OAI21x1_ASAP7_75t_R _25387_ (.A1(net6399),
    .A2(_03006_),
    .B(net6494),
    .Y(_03007_));
 INVx1_ASAP7_75t_R _25388_ (.A(net6494),
    .Y(_03008_));
 INVx1_ASAP7_75t_R _25389_ (.A(_02996_),
    .Y(_03009_));
 NAND3x1_ASAP7_75t_R _25390_ (.A(net6351),
    .B(_03008_),
    .C(_03009_),
    .Y(_03010_));
 NAND2x1_ASAP7_75t_R _25391_ (.A(_03007_),
    .B(_03010_),
    .Y(_03011_));
 NOR2x1_ASAP7_75t_R _25393_ (.A(net6670),
    .B(_00473_),
    .Y(_03012_));
 INVx1_ASAP7_75t_R _25394_ (.A(_03012_),
    .Y(_03013_));
 XOR2x2_ASAP7_75t_R _25395_ (.A(_00585_),
    .B(_00617_),
    .Y(_03014_));
 XOR2x2_ASAP7_75t_R _25396_ (.A(net6414),
    .B(net6557),
    .Y(_03015_));
 NOR2x1_ASAP7_75t_R _25397_ (.A(_03014_),
    .B(_03015_),
    .Y(_03016_));
 INVx1_ASAP7_75t_R _25398_ (.A(net6557),
    .Y(_03017_));
 NOR2x1_ASAP7_75t_R _25399_ (.A(_03017_),
    .B(net6414),
    .Y(_03018_));
 AND2x2_ASAP7_75t_R _25400_ (.A(net6414),
    .B(_03017_),
    .Y(_03019_));
 OAI21x1_ASAP7_75t_R _25401_ (.A1(_03018_),
    .A2(_03019_),
    .B(_03014_),
    .Y(_03020_));
 INVx1_ASAP7_75t_R _25402_ (.A(_03020_),
    .Y(_03021_));
 OAI21x1_ASAP7_75t_R _25403_ (.A1(_03016_),
    .A2(_03021_),
    .B(net6670),
    .Y(_03022_));
 INVx1_ASAP7_75t_R _25404_ (.A(net6511),
    .Y(_03023_));
 AOI21x1_ASAP7_75t_R _25405_ (.A1(_03013_),
    .A2(_03022_),
    .B(_03023_),
    .Y(_03024_));
 NAND2x1_ASAP7_75t_R _25406_ (.A(_00473_),
    .B(net6463),
    .Y(_03025_));
 INVx1_ASAP7_75t_R _25407_ (.A(_03014_),
    .Y(_03026_));
 XOR2x2_ASAP7_75t_R _25408_ (.A(net6414),
    .B(_03017_),
    .Y(_03027_));
 NAND2x1_ASAP7_75t_R _25409_ (.A(_03026_),
    .B(_03027_),
    .Y(_03028_));
 NAND3x1_ASAP7_75t_R _25410_ (.A(_03028_),
    .B(_03020_),
    .C(net6670),
    .Y(_03029_));
 AOI21x1_ASAP7_75t_R _25411_ (.A1(_03025_),
    .A2(_03029_),
    .B(net6511),
    .Y(_03030_));
 NOR2x2_ASAP7_75t_R _25412_ (.A(_03024_),
    .B(_03030_),
    .Y(_03031_));
 AND2x2_ASAP7_75t_R _25414_ (.A(_02995_),
    .B(_02990_),
    .Y(_03032_));
 AOI21x1_ASAP7_75t_R _25416_ (.A1(_03013_),
    .A2(_03022_),
    .B(net6511),
    .Y(_03033_));
 AOI21x1_ASAP7_75t_R _25417_ (.A1(_03025_),
    .A2(_03029_),
    .B(_03023_),
    .Y(_03034_));
 NOR2x2_ASAP7_75t_R _25418_ (.A(_03033_),
    .B(_03034_),
    .Y(_03035_));
 NOR2x1_ASAP7_75t_R _25420_ (.A(net5694),
    .B(net5402),
    .Y(_03036_));
 OAI21x1_ASAP7_75t_R _25422_ (.A1(net6399),
    .A2(_03006_),
    .B(_03008_),
    .Y(_03038_));
 NAND3x1_ASAP7_75t_R _25423_ (.A(_03005_),
    .B(net6494),
    .C(_03009_),
    .Y(_03039_));
 NAND2x2_ASAP7_75t_R _25424_ (.A(_03038_),
    .B(_03039_),
    .Y(_01253_));
 XNOR2x2_ASAP7_75t_R _25425_ (.A(_00682_),
    .B(_14276_),
    .Y(_03040_));
 XNOR2x2_ASAP7_75t_R _25426_ (.A(_00681_),
    .B(net6554),
    .Y(_03041_));
 XOR2x2_ASAP7_75t_R _25427_ (.A(_00586_),
    .B(_00618_),
    .Y(_03042_));
 XOR2x2_ASAP7_75t_R _25428_ (.A(_03041_),
    .B(_03042_),
    .Y(_03043_));
 NOR2x1_ASAP7_75t_R _25429_ (.A(_03040_),
    .B(_03043_),
    .Y(_03044_));
 XOR2x2_ASAP7_75t_R _25430_ (.A(_14276_),
    .B(_00682_),
    .Y(_03045_));
 XNOR2x2_ASAP7_75t_R _25431_ (.A(_03042_),
    .B(_03041_),
    .Y(_03046_));
 OAI21x1_ASAP7_75t_R _25432_ (.A1(_03045_),
    .A2(_03046_),
    .B(net6666),
    .Y(_03047_));
 NAND2x1_ASAP7_75t_R _25433_ (.A(_00505_),
    .B(net6461),
    .Y(_03048_));
 OAI21x1_ASAP7_75t_R _25434_ (.A1(_03044_),
    .A2(_03047_),
    .B(_03048_),
    .Y(_03049_));
 XNOR2x2_ASAP7_75t_R _25435_ (.A(net6510),
    .B(_03049_),
    .Y(_03050_));
 OAI21x1_ASAP7_75t_R _25437_ (.A1(net5399),
    .A2(net5395),
    .B(net6155),
    .Y(_03052_));
 NOR2x1_ASAP7_75t_R _25438_ (.A(net5110),
    .B(_03052_),
    .Y(_03053_));
 NOR2x1_ASAP7_75t_R _25439_ (.A(net5400),
    .B(net5395),
    .Y(_03054_));
 XOR2x2_ASAP7_75t_R _25440_ (.A(_03049_),
    .B(net6510),
    .Y(_03055_));
 OA21x2_ASAP7_75t_R _25443_ (.A1(_03054_),
    .A2(net5111),
    .B(net6151),
    .Y(_03058_));
 XOR2x2_ASAP7_75t_R _25444_ (.A(_00682_),
    .B(net6554),
    .Y(_03059_));
 XOR2x2_ASAP7_75t_R _25445_ (.A(_11503_),
    .B(_03059_),
    .Y(_03060_));
 NAND2x1_ASAP7_75t_R _25446_ (.A(_14299_),
    .B(_03060_),
    .Y(_03061_));
 OA21x2_ASAP7_75t_R _25447_ (.A1(_03060_),
    .A2(_14299_),
    .B(net6666),
    .Y(_03062_));
 AND2x2_ASAP7_75t_R _25448_ (.A(net6461),
    .B(_00504_),
    .Y(_03063_));
 AOI21x1_ASAP7_75t_R _25449_ (.A1(_03061_),
    .A2(_03062_),
    .B(_03063_),
    .Y(_03064_));
 XOR2x2_ASAP7_75t_R _25450_ (.A(_03064_),
    .B(net6509),
    .Y(_03065_));
 INVx2_ASAP7_75t_R _25451_ (.A(_03065_),
    .Y(_03066_));
 OAI21x1_ASAP7_75t_R _25454_ (.A1(_03053_),
    .A2(_03058_),
    .B(net5687),
    .Y(_03069_));
 OA21x2_ASAP7_75t_R _25455_ (.A1(net6158),
    .A2(net5692),
    .B(net5055),
    .Y(_03070_));
 AOI21x1_ASAP7_75t_R _25456_ (.A1(_03020_),
    .A2(_03028_),
    .B(net6463),
    .Y(_03071_));
 OAI21x1_ASAP7_75t_R _25457_ (.A1(_03012_),
    .A2(_03071_),
    .B(_03023_),
    .Y(_03072_));
 NAND3x1_ASAP7_75t_R _25458_ (.A(_03022_),
    .B(net6511),
    .C(_03013_),
    .Y(_03073_));
 INVx1_ASAP7_75t_R _25459_ (.A(_01254_),
    .Y(_03074_));
 AOI21x1_ASAP7_75t_R _25460_ (.A1(_03072_),
    .A2(_03073_),
    .B(_03074_),
    .Y(_03075_));
 OA21x2_ASAP7_75t_R _25461_ (.A1(_03070_),
    .A2(_03075_),
    .B(net6151),
    .Y(_03076_));
 AO21x1_ASAP7_75t_R _25462_ (.A1(_03073_),
    .A2(_03072_),
    .B(_01263_),
    .Y(_03077_));
 OAI21x1_ASAP7_75t_R _25465_ (.A1(net5692),
    .A2(net6158),
    .B(_01255_),
    .Y(_03080_));
 AND3x1_ASAP7_75t_R _25467_ (.A(_03077_),
    .B(net6154),
    .C(net4740),
    .Y(_03082_));
 OAI21x1_ASAP7_75t_R _25470_ (.A1(_03076_),
    .A2(_03082_),
    .B(net6144),
    .Y(_03085_));
 INVx1_ASAP7_75t_R _25471_ (.A(_11483_),
    .Y(_03086_));
 XOR2x2_ASAP7_75t_R _25472_ (.A(_11454_),
    .B(_11508_),
    .Y(_03087_));
 NOR2x1_ASAP7_75t_R _25473_ (.A(_03086_),
    .B(_03087_),
    .Y(_03088_));
 AND2x2_ASAP7_75t_R _25474_ (.A(_03087_),
    .B(_03086_),
    .Y(_03089_));
 OAI21x1_ASAP7_75t_R _25475_ (.A1(_03088_),
    .A2(_03089_),
    .B(net6666),
    .Y(_03090_));
 NOR2x1_ASAP7_75t_R _25476_ (.A(net6665),
    .B(_00503_),
    .Y(_03091_));
 INVx1_ASAP7_75t_R _25477_ (.A(_03091_),
    .Y(_03092_));
 NAND3x1_ASAP7_75t_R _25478_ (.A(_03090_),
    .B(_00874_),
    .C(_03092_),
    .Y(_03093_));
 AO21x1_ASAP7_75t_R _25479_ (.A1(_03090_),
    .A2(_03092_),
    .B(_00874_),
    .Y(_03094_));
 NAND2x1_ASAP7_75t_R _25480_ (.A(_03093_),
    .B(_03094_),
    .Y(_03095_));
 AOI21x1_ASAP7_75t_R _25483_ (.A1(_03069_),
    .A2(_03085_),
    .B(net5681),
    .Y(_03098_));
 XOR2x2_ASAP7_75t_R _25484_ (.A(_14363_),
    .B(net6440),
    .Y(_03099_));
 XOR2x2_ASAP7_75t_R _25485_ (.A(_03099_),
    .B(_11411_),
    .Y(_03100_));
 NOR2x1_ASAP7_75t_R _25486_ (.A(net6665),
    .B(_00501_),
    .Y(_03101_));
 AO21x1_ASAP7_75t_R _25487_ (.A1(_03100_),
    .A2(net6665),
    .B(_03101_),
    .Y(_03102_));
 XOR2x2_ASAP7_75t_R _25488_ (.A(_03102_),
    .B(_00876_),
    .Y(_03103_));
 NAND2x2_ASAP7_75t_R _25490_ (.A(net5400),
    .B(net5690),
    .Y(_03105_));
 NAND2x1_ASAP7_75t_R _25491_ (.A(net4740),
    .B(_03105_),
    .Y(_03106_));
 OAI21x1_ASAP7_75t_R _25492_ (.A1(net5689),
    .A2(net6157),
    .B(_01255_),
    .Y(_03107_));
 AO21x1_ASAP7_75t_R _25495_ (.A1(net4739),
    .A2(net6149),
    .B(net6145),
    .Y(_03110_));
 AOI21x1_ASAP7_75t_R _25496_ (.A1(net6155),
    .A2(_03106_),
    .B(_03110_),
    .Y(_03111_));
 INVx1_ASAP7_75t_R _25497_ (.A(_01258_),
    .Y(_03112_));
 AOI21x1_ASAP7_75t_R _25498_ (.A1(_03072_),
    .A2(_03073_),
    .B(_03112_),
    .Y(_03113_));
 OAI21x1_ASAP7_75t_R _25499_ (.A1(net5692),
    .A2(net6158),
    .B(_01254_),
    .Y(_03114_));
 INVx1_ASAP7_75t_R _25500_ (.A(_03114_),
    .Y(_03115_));
 OAI21x1_ASAP7_75t_R _25501_ (.A1(net4657),
    .A2(_03115_),
    .B(net6153),
    .Y(_03116_));
 INVx1_ASAP7_75t_R _25502_ (.A(_01255_),
    .Y(_03117_));
 OA21x2_ASAP7_75t_R _25503_ (.A1(net6158),
    .A2(net5692),
    .B(_03117_),
    .Y(_03118_));
 OAI21x1_ASAP7_75t_R _25506_ (.A1(_03075_),
    .A2(_03118_),
    .B(net6146),
    .Y(_03121_));
 AOI21x1_ASAP7_75t_R _25508_ (.A1(_03116_),
    .A2(_03121_),
    .B(net5686),
    .Y(_03123_));
 OAI21x1_ASAP7_75t_R _25510_ (.A1(_03111_),
    .A2(_03123_),
    .B(net5681),
    .Y(_03125_));
 NAND2x1_ASAP7_75t_R _25511_ (.A(net6142),
    .B(_03125_),
    .Y(_03126_));
 NOR2x1_ASAP7_75t_R _25512_ (.A(_03098_),
    .B(_03126_),
    .Y(_03127_));
 NAND3x1_ASAP7_75t_R _25513_ (.A(_03022_),
    .B(_03023_),
    .C(_03013_),
    .Y(_03128_));
 INVx2_ASAP7_75t_R _25514_ (.A(net5692),
    .Y(_03129_));
 AO21x1_ASAP7_75t_R _25515_ (.A1(_03128_),
    .A2(_03129_),
    .B(net5057),
    .Y(_03130_));
 AOI21x1_ASAP7_75t_R _25516_ (.A1(net5399),
    .A2(net5395),
    .B(net6155),
    .Y(_03131_));
 NAND2x1_ASAP7_75t_R _25517_ (.A(_03130_),
    .B(_03131_),
    .Y(_03132_));
 INVx1_ASAP7_75t_R _25518_ (.A(net5056),
    .Y(_03133_));
 OAI21x1_ASAP7_75t_R _25519_ (.A1(net5689),
    .A2(net6157),
    .B(_03133_),
    .Y(_03134_));
 OA21x2_ASAP7_75t_R _25521_ (.A1(_03134_),
    .A2(net6147),
    .B(net6144),
    .Y(_03136_));
 INVx1_ASAP7_75t_R _25522_ (.A(_01262_),
    .Y(_03137_));
 OAI21x1_ASAP7_75t_R _25523_ (.A1(net5689),
    .A2(net6157),
    .B(_03137_),
    .Y(_03138_));
 OAI21x1_ASAP7_75t_R _25524_ (.A1(net5692),
    .A2(net6158),
    .B(net5053),
    .Y(_03139_));
 AO21x1_ASAP7_75t_R _25525_ (.A1(net4655),
    .A2(_03139_),
    .B(net6147),
    .Y(_03140_));
 AND2x2_ASAP7_75t_R _25526_ (.A(_03136_),
    .B(_03140_),
    .Y(_03141_));
 AOI21x1_ASAP7_75t_R _25527_ (.A1(_03072_),
    .A2(_03073_),
    .B(_01255_),
    .Y(_03142_));
 NOR2x1_ASAP7_75t_R _25529_ (.A(_01272_),
    .B(net6154),
    .Y(_03144_));
 AO21x1_ASAP7_75t_R _25530_ (.A1(net4738),
    .A2(net6154),
    .B(_03144_),
    .Y(_03145_));
 OAI21x1_ASAP7_75t_R _25531_ (.A1(net6144),
    .A2(_03145_),
    .B(net5681),
    .Y(_03146_));
 AOI21x1_ASAP7_75t_R _25532_ (.A1(_03132_),
    .A2(_03141_),
    .B(_03146_),
    .Y(_03147_));
 INVx1_ASAP7_75t_R _25533_ (.A(_01261_),
    .Y(_03148_));
 AOI21x1_ASAP7_75t_R _25535_ (.A1(_03148_),
    .A2(net5396),
    .B(net6155),
    .Y(_03150_));
 INVx1_ASAP7_75t_R _25536_ (.A(_01259_),
    .Y(_03151_));
 AO21x1_ASAP7_75t_R _25537_ (.A1(net5682),
    .A2(_03072_),
    .B(_03151_),
    .Y(_03152_));
 AOI21x1_ASAP7_75t_R _25539_ (.A1(_03129_),
    .A2(_03128_),
    .B(net5056),
    .Y(_03154_));
 NAND2x1_ASAP7_75t_R _25540_ (.A(net6154),
    .B(net4876),
    .Y(_03155_));
 INVx1_ASAP7_75t_R _25541_ (.A(_03155_),
    .Y(_03156_));
 AOI211x1_ASAP7_75t_R _25542_ (.A1(_03150_),
    .A2(_03152_),
    .B(_03156_),
    .C(net5686),
    .Y(_03157_));
 OA21x2_ASAP7_75t_R _25543_ (.A1(_03139_),
    .A2(net6148),
    .B(_03066_),
    .Y(_03158_));
 INVx1_ASAP7_75t_R _25544_ (.A(_03158_),
    .Y(_03159_));
 INVx1_ASAP7_75t_R _25545_ (.A(_03154_),
    .Y(_03160_));
 NAND2x1_ASAP7_75t_R _25546_ (.A(net6153),
    .B(net4656),
    .Y(_03161_));
 OAI21x1_ASAP7_75t_R _25547_ (.A1(net6154),
    .A2(net4654),
    .B(_03161_),
    .Y(_03162_));
 INVx1_ASAP7_75t_R _25548_ (.A(_03095_),
    .Y(_03163_));
 OAI21x1_ASAP7_75t_R _25550_ (.A1(_03159_),
    .A2(_03162_),
    .B(net5393),
    .Y(_03165_));
 INVx1_ASAP7_75t_R _25551_ (.A(_03103_),
    .Y(_03166_));
 OAI21x1_ASAP7_75t_R _25553_ (.A1(_03157_),
    .A2(_03165_),
    .B(net5680),
    .Y(_03168_));
 XOR2x2_ASAP7_75t_R _25554_ (.A(net6555),
    .B(_00685_),
    .Y(_03169_));
 XOR2x2_ASAP7_75t_R _25555_ (.A(_03169_),
    .B(net6588),
    .Y(_03170_));
 XOR2x2_ASAP7_75t_R _25556_ (.A(_03170_),
    .B(_11564_),
    .Y(_03171_));
 NOR2x1_ASAP7_75t_R _25557_ (.A(net6665),
    .B(_00502_),
    .Y(_03172_));
 AO21x1_ASAP7_75t_R _25558_ (.A1(_03171_),
    .A2(net6665),
    .B(_03172_),
    .Y(_03173_));
 XOR2x2_ASAP7_75t_R _25559_ (.A(_03173_),
    .B(_00875_),
    .Y(_03174_));
 OAI21x1_ASAP7_75t_R _25561_ (.A1(_03147_),
    .A2(_03168_),
    .B(net6141),
    .Y(_03176_));
 AOI21x1_ASAP7_75t_R _25562_ (.A1(_03160_),
    .A2(_03105_),
    .B(net6148),
    .Y(_03177_));
 AO21x1_ASAP7_75t_R _25563_ (.A1(_03128_),
    .A2(_03129_),
    .B(_01263_),
    .Y(_03178_));
 INVx1_ASAP7_75t_R _25564_ (.A(_03178_),
    .Y(_03179_));
 OAI21x1_ASAP7_75t_R _25566_ (.A1(net5398),
    .A2(net5402),
    .B(net6152),
    .Y(_03181_));
 OAI21x1_ASAP7_75t_R _25568_ (.A1(net4653),
    .A2(_03181_),
    .B(net6144),
    .Y(_03183_));
 OAI21x1_ASAP7_75t_R _25569_ (.A1(net4507),
    .A2(_03183_),
    .B(net5681),
    .Y(_03184_));
 INVx1_ASAP7_75t_R _25570_ (.A(_01264_),
    .Y(_03185_));
 AO21x1_ASAP7_75t_R _25571_ (.A1(_03128_),
    .A2(_03129_),
    .B(_03185_),
    .Y(_03186_));
 INVx1_ASAP7_75t_R _25572_ (.A(_03186_),
    .Y(_03187_));
 OAI21x1_ASAP7_75t_R _25574_ (.A1(_03187_),
    .A2(_03181_),
    .B(net5687),
    .Y(_03189_));
 NOR2x2_ASAP7_75t_R _25575_ (.A(net5694),
    .B(net5400),
    .Y(_03190_));
 NOR2x1_ASAP7_75t_R _25576_ (.A(net5053),
    .B(net5398),
    .Y(_03191_));
 NOR3x1_ASAP7_75t_R _25578_ (.A(_03190_),
    .B(_03191_),
    .C(net6148),
    .Y(_03193_));
 NOR2x1_ASAP7_75t_R _25579_ (.A(_03189_),
    .B(_03193_),
    .Y(_03194_));
 OAI21x1_ASAP7_75t_R _25580_ (.A1(_03184_),
    .A2(_03194_),
    .B(net6142),
    .Y(_03195_));
 AOI21x1_ASAP7_75t_R _25581_ (.A1(net5399),
    .A2(net5395),
    .B(net6152),
    .Y(_03196_));
 AOI21x1_ASAP7_75t_R _25582_ (.A1(net5051),
    .A2(_03035_),
    .B(net6155),
    .Y(_03197_));
 INVx1_ASAP7_75t_R _25583_ (.A(_03197_),
    .Y(_03198_));
 NOR2x1_ASAP7_75t_R _25584_ (.A(_03191_),
    .B(_03198_),
    .Y(_03199_));
 OAI21x1_ASAP7_75t_R _25585_ (.A1(_03196_),
    .A2(_03199_),
    .B(net6144),
    .Y(_03200_));
 NAND2x1_ASAP7_75t_R _25586_ (.A(net5396),
    .B(net5395),
    .Y(_03201_));
 AOI21x1_ASAP7_75t_R _25587_ (.A1(_03148_),
    .A2(net5399),
    .B(net6150),
    .Y(_03202_));
 NAND2x1_ASAP7_75t_R _25588_ (.A(_03201_),
    .B(_03202_),
    .Y(_03203_));
 AOI21x1_ASAP7_75t_R _25589_ (.A1(net5049),
    .A2(net5399),
    .B(net6155),
    .Y(_03204_));
 NAND2x1_ASAP7_75t_R _25590_ (.A(net4740),
    .B(_03204_),
    .Y(_03205_));
 AO21x1_ASAP7_75t_R _25591_ (.A1(_03203_),
    .A2(_03205_),
    .B(net6143),
    .Y(_03206_));
 AOI21x1_ASAP7_75t_R _25592_ (.A1(_03200_),
    .A2(_03206_),
    .B(net5681),
    .Y(_03207_));
 INVx1_ASAP7_75t_R _25593_ (.A(_03174_),
    .Y(_03208_));
 OAI21x1_ASAP7_75t_R _25595_ (.A1(_03195_),
    .A2(_03207_),
    .B(net5679),
    .Y(_03210_));
 OA21x2_ASAP7_75t_R _25596_ (.A1(net4876),
    .A2(_03075_),
    .B(net6154),
    .Y(_03211_));
 NAND2x1_ASAP7_75t_R _25598_ (.A(net5687),
    .B(_03198_),
    .Y(_03213_));
 NOR2x1_ASAP7_75t_R _25599_ (.A(_03211_),
    .B(_03213_),
    .Y(_03214_));
 AOI21x1_ASAP7_75t_R _25600_ (.A1(net5694),
    .A2(net5398),
    .B(net6152),
    .Y(_03215_));
 INVx2_ASAP7_75t_R _25601_ (.A(_03142_),
    .Y(_03216_));
 AND2x4_ASAP7_75t_R _25602_ (.A(_03215_),
    .B(_03216_),
    .Y(_03217_));
 NOR2x1_ASAP7_75t_R _25603_ (.A(net5055),
    .B(_03035_),
    .Y(_03218_));
 OAI21x1_ASAP7_75t_R _25604_ (.A1(net5400),
    .A2(net5402),
    .B(net6152),
    .Y(_03219_));
 OAI21x1_ASAP7_75t_R _25606_ (.A1(_03218_),
    .A2(_03219_),
    .B(net6144),
    .Y(_03221_));
 NOR2x1p5_ASAP7_75t_R _25607_ (.A(net4463),
    .B(_03221_),
    .Y(_03222_));
 OAI21x1_ASAP7_75t_R _25608_ (.A1(_03222_),
    .A2(_03214_),
    .B(net5394),
    .Y(_03223_));
 AOI21x1_ASAP7_75t_R _25609_ (.A1(net4875),
    .A2(_03131_),
    .B(net5686),
    .Y(_03224_));
 OAI21x1_ASAP7_75t_R _25610_ (.A1(net5692),
    .A2(net6158),
    .B(_03151_),
    .Y(_03225_));
 INVx1_ASAP7_75t_R _25611_ (.A(_03225_),
    .Y(_03226_));
 NAND2x1_ASAP7_75t_R _25612_ (.A(net6153),
    .B(net4506),
    .Y(_03227_));
 NAND2x1p5_ASAP7_75t_R _25613_ (.A(net6150),
    .B(_03080_),
    .Y(_03228_));
 AND3x1_ASAP7_75t_R _25614_ (.A(_03227_),
    .B(net5685),
    .C(net4557),
    .Y(_03229_));
 OA21x2_ASAP7_75t_R _25616_ (.A1(net4655),
    .A2(net6147),
    .B(net5681),
    .Y(_03231_));
 OAI21x1_ASAP7_75t_R _25617_ (.A1(_03224_),
    .A2(_03229_),
    .B(_03231_),
    .Y(_03232_));
 AOI21x1_ASAP7_75t_R _25618_ (.A1(_03232_),
    .A2(_03223_),
    .B(net6142),
    .Y(_03233_));
 OAI22x1_ASAP7_75t_R _25619_ (.A1(_03127_),
    .A2(_03176_),
    .B1(_03210_),
    .B2(_03233_),
    .Y(_00104_));
 AO21x1_ASAP7_75t_R _25620_ (.A1(net5400),
    .A2(net5056),
    .B(net6152),
    .Y(_03234_));
 NOR2x1_ASAP7_75t_R _25621_ (.A(_03187_),
    .B(_03234_),
    .Y(_03235_));
 INVx2_ASAP7_75t_R _25622_ (.A(_03080_),
    .Y(_03236_));
 OA21x2_ASAP7_75t_R _25623_ (.A1(net6157),
    .A2(net5689),
    .B(net5050),
    .Y(_03237_));
 OAI21x1_ASAP7_75t_R _25624_ (.A1(_03236_),
    .A2(_03237_),
    .B(net6149),
    .Y(_03238_));
 NAND2x1_ASAP7_75t_R _25625_ (.A(net5686),
    .B(_03238_),
    .Y(_03239_));
 NOR2x1_ASAP7_75t_R _25626_ (.A(_03235_),
    .B(_03239_),
    .Y(_03240_));
 AO21x1_ASAP7_75t_R _25627_ (.A1(net4740),
    .A2(net6151),
    .B(net5687),
    .Y(_03241_));
 AND2x2_ASAP7_75t_R _25628_ (.A(_03196_),
    .B(net4875),
    .Y(_03242_));
 OAI21x1_ASAP7_75t_R _25629_ (.A1(_03241_),
    .A2(_03242_),
    .B(net5681),
    .Y(_03243_));
 NOR2x1_ASAP7_75t_R _25630_ (.A(net5057),
    .B(net5398),
    .Y(_03244_));
 OAI21x1_ASAP7_75t_R _25631_ (.A1(_03244_),
    .A2(_03052_),
    .B(net6144),
    .Y(_03245_));
 AOI21x1_ASAP7_75t_R _25632_ (.A1(_03197_),
    .A2(_03105_),
    .B(_03245_),
    .Y(_03246_));
 NAND2x1_ASAP7_75t_R _25633_ (.A(net5399),
    .B(net5401),
    .Y(_03247_));
 OAI21x1_ASAP7_75t_R _25634_ (.A1(net6147),
    .A2(_03247_),
    .B(net5686),
    .Y(_03248_));
 NAND2x1p5_ASAP7_75t_R _25635_ (.A(_03107_),
    .B(net6150),
    .Y(_03249_));
 INVx1_ASAP7_75t_R _25636_ (.A(_03130_),
    .Y(_03250_));
 OAI21x1_ASAP7_75t_R _25637_ (.A1(net4556),
    .A2(_03250_),
    .B(_03155_),
    .Y(_03251_));
 OAI21x1_ASAP7_75t_R _25638_ (.A1(_03248_),
    .A2(_03251_),
    .B(net5394),
    .Y(_03252_));
 OAI22x1_ASAP7_75t_R _25639_ (.A1(_03240_),
    .A2(_03243_),
    .B1(_03246_),
    .B2(_03252_),
    .Y(_03253_));
 AOI21x1_ASAP7_75t_R _25640_ (.A1(_03105_),
    .A2(_03197_),
    .B(net6144),
    .Y(_03254_));
 NOR2x1_ASAP7_75t_R _25642_ (.A(net5398),
    .B(net5690),
    .Y(_03256_));
 NOR2x1_ASAP7_75t_R _25643_ (.A(_03256_),
    .B(_03052_),
    .Y(_03257_));
 NOR2x1_ASAP7_75t_R _25644_ (.A(net5394),
    .B(_03257_),
    .Y(_03258_));
 OA21x2_ASAP7_75t_R _25645_ (.A1(net6158),
    .A2(net5692),
    .B(_01263_),
    .Y(_03259_));
 OAI21x1_ASAP7_75t_R _25646_ (.A1(_03113_),
    .A2(_03259_),
    .B(net6153),
    .Y(_03260_));
 INVx1_ASAP7_75t_R _25647_ (.A(_03260_),
    .Y(_03261_));
 INVx1_ASAP7_75t_R _25648_ (.A(_01269_),
    .Y(_03262_));
 AO21x1_ASAP7_75t_R _25650_ (.A1(_03093_),
    .A2(_03094_),
    .B(net6153),
    .Y(_03264_));
 OAI21x1_ASAP7_75t_R _25651_ (.A1(_03262_),
    .A2(_03264_),
    .B(net6144),
    .Y(_03265_));
 OAI21x1_ASAP7_75t_R _25652_ (.A1(_03261_),
    .A2(_03265_),
    .B(net6141),
    .Y(_03266_));
 AOI21x1_ASAP7_75t_R _25653_ (.A1(_03148_),
    .A2(net5399),
    .B(net6155),
    .Y(_03267_));
 NOR2x1_ASAP7_75t_R _25654_ (.A(net5400),
    .B(net5402),
    .Y(_03268_));
 OAI21x1_ASAP7_75t_R _25655_ (.A1(net5057),
    .A2(net5398),
    .B(net6155),
    .Y(_03269_));
 NOR2x1_ASAP7_75t_R _25656_ (.A(net6144),
    .B(net5681),
    .Y(_03270_));
 OAI21x1_ASAP7_75t_R _25657_ (.A1(_03268_),
    .A2(_03269_),
    .B(_03270_),
    .Y(_03271_));
 AOI21x1_ASAP7_75t_R _25658_ (.A1(net4875),
    .A2(_03267_),
    .B(_03271_),
    .Y(_03272_));
 AOI211x1_ASAP7_75t_R _25659_ (.A1(net4651),
    .A2(_03258_),
    .B(_03266_),
    .C(_03272_),
    .Y(_03273_));
 AOI21x1_ASAP7_75t_R _25660_ (.A1(net5679),
    .A2(_03253_),
    .B(_03273_),
    .Y(_03274_));
 AOI21x1_ASAP7_75t_R _25661_ (.A1(_03072_),
    .A2(_03073_),
    .B(_03148_),
    .Y(_03275_));
 AOI21x1_ASAP7_75t_R _25663_ (.A1(net6147),
    .A2(_03275_),
    .B(net5685),
    .Y(_03277_));
 INVx1_ASAP7_75t_R _25664_ (.A(net5111),
    .Y(_03278_));
 NAND2x1_ASAP7_75t_R _25665_ (.A(_03215_),
    .B(_03278_),
    .Y(_03279_));
 AOI21x1_ASAP7_75t_R _25666_ (.A1(_03277_),
    .A2(_03279_),
    .B(net5681),
    .Y(_03280_));
 NOR2x1_ASAP7_75t_R _25667_ (.A(net5396),
    .B(net5401),
    .Y(_03281_));
 AOI21x1_ASAP7_75t_R _25668_ (.A1(net5051),
    .A2(_03035_),
    .B(net6150),
    .Y(_03282_));
 AOI21x1_ASAP7_75t_R _25669_ (.A1(_03247_),
    .A2(_03282_),
    .B(net6143),
    .Y(_03283_));
 OAI21x1_ASAP7_75t_R _25670_ (.A1(_03281_),
    .A2(net4557),
    .B(_03283_),
    .Y(_03284_));
 AOI21x1_ASAP7_75t_R _25671_ (.A1(_03280_),
    .A2(_03284_),
    .B(net5679),
    .Y(_03285_));
 NAND2x1_ASAP7_75t_R _25672_ (.A(net6153),
    .B(_03190_),
    .Y(_03286_));
 NAND2x1_ASAP7_75t_R _25674_ (.A(_01273_),
    .B(net6147),
    .Y(_03288_));
 OA21x2_ASAP7_75t_R _25675_ (.A1(net6147),
    .A2(net4655),
    .B(_03288_),
    .Y(_03289_));
 AOI21x1_ASAP7_75t_R _25676_ (.A1(_03286_),
    .A2(_03289_),
    .B(net6143),
    .Y(_03290_));
 INVx2_ASAP7_75t_R _25677_ (.A(_03249_),
    .Y(_03291_));
 NAND2x1p5_ASAP7_75t_R _25678_ (.A(_03186_),
    .B(_03291_),
    .Y(_03292_));
 AOI21x1_ASAP7_75t_R _25679_ (.A1(_03140_),
    .A2(net4432),
    .B(net5686),
    .Y(_03293_));
 OAI21x1_ASAP7_75t_R _25680_ (.A1(_03290_),
    .A2(_03293_),
    .B(net5681),
    .Y(_03294_));
 NAND2x1_ASAP7_75t_R _25681_ (.A(_03285_),
    .B(_03294_),
    .Y(_03295_));
 INVx1_ASAP7_75t_R _25682_ (.A(_03138_),
    .Y(_03296_));
 NOR2x1_ASAP7_75t_R _25683_ (.A(_03296_),
    .B(_03228_),
    .Y(_03297_));
 OAI21x1_ASAP7_75t_R _25684_ (.A1(net5396),
    .A2(net5395),
    .B(net6153),
    .Y(_03298_));
 NOR2x1_ASAP7_75t_R _25685_ (.A(_03115_),
    .B(_03298_),
    .Y(_03299_));
 OAI21x1_ASAP7_75t_R _25686_ (.A1(_03297_),
    .A2(_03299_),
    .B(net5684),
    .Y(_03300_));
 INVx1_ASAP7_75t_R _25687_ (.A(net4739),
    .Y(_03301_));
 OAI21x1_ASAP7_75t_R _25688_ (.A1(_03301_),
    .A2(_03054_),
    .B(net6153),
    .Y(_03302_));
 NAND2x1_ASAP7_75t_R _25689_ (.A(net5401),
    .B(net5691),
    .Y(_03303_));
 AOI21x1_ASAP7_75t_R _25690_ (.A1(_03303_),
    .A2(_03131_),
    .B(net5683),
    .Y(_03304_));
 AOI21x1_ASAP7_75t_R _25691_ (.A1(_03302_),
    .A2(_03304_),
    .B(net5391),
    .Y(_03305_));
 NAND2x1_ASAP7_75t_R _25692_ (.A(_03300_),
    .B(_03305_),
    .Y(_03306_));
 NAND2x1_ASAP7_75t_R _25693_ (.A(net4877),
    .B(net6153),
    .Y(_03307_));
 OA21x2_ASAP7_75t_R _25694_ (.A1(_03307_),
    .A2(net5399),
    .B(net6144),
    .Y(_03308_));
 AOI21x1_ASAP7_75t_R _25695_ (.A1(_03238_),
    .A2(_03308_),
    .B(net5681),
    .Y(_03309_));
 INVx1_ASAP7_75t_R _25696_ (.A(net5050),
    .Y(_03310_));
 AO21x1_ASAP7_75t_R _25697_ (.A1(_03128_),
    .A2(_03129_),
    .B(_03310_),
    .Y(_03311_));
 NAND2x2_ASAP7_75t_R _25698_ (.A(net5398),
    .B(net5690),
    .Y(_03312_));
 AOI21x1_ASAP7_75t_R _25699_ (.A1(_03312_),
    .A2(_03204_),
    .B(net6144),
    .Y(_03313_));
 OAI21x1_ASAP7_75t_R _25700_ (.A1(net6150),
    .A2(_03311_),
    .B(_03313_),
    .Y(_03314_));
 AOI21x1_ASAP7_75t_R _25701_ (.A1(_03309_),
    .A2(_03314_),
    .B(net6141),
    .Y(_03315_));
 AOI21x1_ASAP7_75t_R _25702_ (.A1(_03306_),
    .A2(_03315_),
    .B(net6142),
    .Y(_03316_));
 NAND2x1_ASAP7_75t_R _25703_ (.A(_03316_),
    .B(_03295_),
    .Y(_03317_));
 OAI21x1_ASAP7_75t_R _25704_ (.A1(net5680),
    .A2(_03274_),
    .B(_03317_),
    .Y(_00105_));
 NOR2x1_ASAP7_75t_R _25705_ (.A(_03262_),
    .B(net6151),
    .Y(_03318_));
 AO21x1_ASAP7_75t_R _25706_ (.A1(net5398),
    .A2(net5694),
    .B(net6155),
    .Y(_03319_));
 OAI21x1_ASAP7_75t_R _25707_ (.A1(net5111),
    .A2(_03319_),
    .B(net6144),
    .Y(_03320_));
 OAI21x1_ASAP7_75t_R _25708_ (.A1(_03318_),
    .A2(_03320_),
    .B(net5681),
    .Y(_03321_));
 OA21x2_ASAP7_75t_R _25709_ (.A1(_03074_),
    .A2(net5397),
    .B(_03215_),
    .Y(_03322_));
 NAND2x1p5_ASAP7_75t_R _25710_ (.A(_03216_),
    .B(net6148),
    .Y(_03323_));
 NOR2x1_ASAP7_75t_R _25711_ (.A(_03070_),
    .B(_03323_),
    .Y(_03324_));
 OA21x2_ASAP7_75t_R _25712_ (.A1(_03322_),
    .A2(_03324_),
    .B(net5687),
    .Y(_03325_));
 OAI21x1_ASAP7_75t_R _25713_ (.A1(_03321_),
    .A2(_03325_),
    .B(net5680),
    .Y(_03326_));
 AO21x1_ASAP7_75t_R _25714_ (.A1(_03128_),
    .A2(_03129_),
    .B(net5053),
    .Y(_03327_));
 NOR2x1_ASAP7_75t_R _25715_ (.A(_01272_),
    .B(net6151),
    .Y(_03328_));
 AO21x1_ASAP7_75t_R _25716_ (.A1(_03291_),
    .A2(_03327_),
    .B(_03328_),
    .Y(_03329_));
 NAND2x1_ASAP7_75t_R _25717_ (.A(net6144),
    .B(_03329_),
    .Y(_03330_));
 AO21x1_ASAP7_75t_R _25718_ (.A1(net5690),
    .A2(net5400),
    .B(_03219_),
    .Y(_03331_));
 INVx1_ASAP7_75t_R _25719_ (.A(_03217_),
    .Y(_03332_));
 AO21x1_ASAP7_75t_R _25720_ (.A1(_03331_),
    .A2(_03332_),
    .B(net6144),
    .Y(_03333_));
 AOI21x1_ASAP7_75t_R _25721_ (.A1(_03330_),
    .A2(_03333_),
    .B(net5681),
    .Y(_03334_));
 NOR2x1_ASAP7_75t_R _25722_ (.A(_03334_),
    .B(_03326_),
    .Y(_03335_));
 AO21x1_ASAP7_75t_R _25723_ (.A1(net4652),
    .A2(_03138_),
    .B(net6147),
    .Y(_03336_));
 AOI21x1_ASAP7_75t_R _25724_ (.A1(net5052),
    .A2(net5399),
    .B(net6153),
    .Y(_03337_));
 NAND2x1_ASAP7_75t_R _25725_ (.A(_03312_),
    .B(_03337_),
    .Y(_03338_));
 AOI21x1_ASAP7_75t_R _25726_ (.A1(_03336_),
    .A2(_03338_),
    .B(net5684),
    .Y(_03339_));
 NAND2x1_ASAP7_75t_R _25727_ (.A(_03201_),
    .B(_03337_),
    .Y(_03340_));
 NOR2x1_ASAP7_75t_R _25728_ (.A(net5049),
    .B(net5396),
    .Y(_03341_));
 OAI21x1_ASAP7_75t_R _25729_ (.A1(_03226_),
    .A2(_03341_),
    .B(net6153),
    .Y(_03342_));
 AOI21x1_ASAP7_75t_R _25730_ (.A1(_03340_),
    .A2(_03342_),
    .B(net6145),
    .Y(_03343_));
 OAI21x1_ASAP7_75t_R _25731_ (.A1(_03339_),
    .A2(_03343_),
    .B(net5681),
    .Y(_03344_));
 OAI21x1_ASAP7_75t_R _25732_ (.A1(_03301_),
    .A2(net4558),
    .B(net6147),
    .Y(_03345_));
 AOI21x1_ASAP7_75t_R _25733_ (.A1(net5054),
    .A2(net5399),
    .B(net6150),
    .Y(_03346_));
 NAND2x1_ASAP7_75t_R _25734_ (.A(_03201_),
    .B(_03346_),
    .Y(_03347_));
 AOI21x1_ASAP7_75t_R _25735_ (.A1(_03345_),
    .A2(_03347_),
    .B(net5684),
    .Y(_03348_));
 AOI211x1_ASAP7_75t_R _25736_ (.A1(net5691),
    .A2(net5399),
    .B(_03226_),
    .C(net6153),
    .Y(_03349_));
 OAI21x1_ASAP7_75t_R _25737_ (.A1(_03341_),
    .A2(_03052_),
    .B(net5685),
    .Y(_03350_));
 NOR2x1_ASAP7_75t_R _25738_ (.A(_03349_),
    .B(_03350_),
    .Y(_03351_));
 OAI21x1_ASAP7_75t_R _25739_ (.A1(_03348_),
    .A2(_03351_),
    .B(net5392),
    .Y(_03352_));
 NAND2x1_ASAP7_75t_R _25740_ (.A(_03344_),
    .B(_03352_),
    .Y(_03353_));
 OAI21x1_ASAP7_75t_R _25741_ (.A1(net5680),
    .A2(_03353_),
    .B(net5679),
    .Y(_03354_));
 NAND2x1_ASAP7_75t_R _25742_ (.A(net6153),
    .B(_03115_),
    .Y(_03355_));
 OAI21x1_ASAP7_75t_R _25743_ (.A1(_03296_),
    .A2(net4558),
    .B(net6147),
    .Y(_03356_));
 AOI21x1_ASAP7_75t_R _25744_ (.A1(_03355_),
    .A2(_03356_),
    .B(net5684),
    .Y(_03357_));
 AND2x2_ASAP7_75t_R _25745_ (.A(_01256_),
    .B(_01262_),
    .Y(_03358_));
 INVx1_ASAP7_75t_R _25746_ (.A(_03358_),
    .Y(_03359_));
 OAI21x1_ASAP7_75t_R _25747_ (.A1(net5692),
    .A2(net6158),
    .B(_03359_),
    .Y(_03360_));
 INVx1_ASAP7_75t_R _25748_ (.A(_03360_),
    .Y(_03361_));
 OAI21x1_ASAP7_75t_R _25749_ (.A1(_03361_),
    .A2(_03237_),
    .B(net6146),
    .Y(_03362_));
 AOI21x1_ASAP7_75t_R _25750_ (.A1(_03260_),
    .A2(_03362_),
    .B(net6145),
    .Y(_03363_));
 OAI21x1_ASAP7_75t_R _25751_ (.A1(_03357_),
    .A2(_03363_),
    .B(net5392),
    .Y(_03364_));
 AND2x2_ASAP7_75t_R _25753_ (.A(net6150),
    .B(_01271_),
    .Y(_03366_));
 NOR2x1_ASAP7_75t_R _25754_ (.A(_03366_),
    .B(_03202_),
    .Y(_03367_));
 NAND2x1_ASAP7_75t_R _25755_ (.A(net6145),
    .B(_03367_),
    .Y(_03368_));
 OA21x2_ASAP7_75t_R _25756_ (.A1(_01274_),
    .A2(net6147),
    .B(net5684),
    .Y(_03369_));
 NAND2x1_ASAP7_75t_R _25757_ (.A(net5693),
    .B(net5396),
    .Y(_03370_));
 NAND2x1_ASAP7_75t_R _25758_ (.A(_03370_),
    .B(_03267_),
    .Y(_03371_));
 AOI21x1_ASAP7_75t_R _25759_ (.A1(_03369_),
    .A2(_03371_),
    .B(net5392),
    .Y(_03372_));
 AOI21x1_ASAP7_75t_R _25760_ (.A1(_03368_),
    .A2(_03372_),
    .B(net6142),
    .Y(_03373_));
 AOI21x1_ASAP7_75t_R _25761_ (.A1(_03364_),
    .A2(_03373_),
    .B(net5679),
    .Y(_03374_));
 AO21x1_ASAP7_75t_R _25762_ (.A1(_03073_),
    .A2(_03072_),
    .B(_03185_),
    .Y(_03375_));
 NAND2x1_ASAP7_75t_R _25763_ (.A(_03375_),
    .B(_03282_),
    .Y(_03376_));
 AOI21x1_ASAP7_75t_R _25764_ (.A1(_03371_),
    .A2(_03376_),
    .B(net6145),
    .Y(_03377_));
 NAND2x1_ASAP7_75t_R _25765_ (.A(net6147),
    .B(_03139_),
    .Y(_03378_));
 OAI21x1_ASAP7_75t_R _25766_ (.A1(_03296_),
    .A2(_03378_),
    .B(net6145),
    .Y(_03379_));
 OAI21x1_ASAP7_75t_R _25767_ (.A1(_03379_),
    .A2(_03217_),
    .B(net5681),
    .Y(_03380_));
 NOR2x1_ASAP7_75t_R _25768_ (.A(_03377_),
    .B(_03380_),
    .Y(_03381_));
 NAND2x1_ASAP7_75t_R _25769_ (.A(net6150),
    .B(_03134_),
    .Y(_03382_));
 NOR2x1_ASAP7_75t_R _25770_ (.A(_03054_),
    .B(_03382_),
    .Y(_03383_));
 OAI21x1_ASAP7_75t_R _25771_ (.A1(net5693),
    .A2(net5396),
    .B(net6153),
    .Y(_03384_));
 OAI21x1_ASAP7_75t_R _25772_ (.A1(net4558),
    .A2(_03384_),
    .B(net5684),
    .Y(_03385_));
 OAI21x1_ASAP7_75t_R _25773_ (.A1(_03383_),
    .A2(_03385_),
    .B(net5391),
    .Y(_03386_));
 INVx1_ASAP7_75t_R _25774_ (.A(_03202_),
    .Y(_03387_));
 NAND3x1_ASAP7_75t_R _25775_ (.A(_03186_),
    .B(_03077_),
    .C(net6148),
    .Y(_03388_));
 AOI21x1_ASAP7_75t_R _25776_ (.A1(_03387_),
    .A2(_03388_),
    .B(net5686),
    .Y(_03389_));
 NOR2x1_ASAP7_75t_R _25777_ (.A(_03386_),
    .B(_03389_),
    .Y(_03390_));
 OAI21x1_ASAP7_75t_R _25778_ (.A1(_03381_),
    .A2(_03390_),
    .B(net6142),
    .Y(_03391_));
 NAND2x1_ASAP7_75t_R _25779_ (.A(_03374_),
    .B(_03391_),
    .Y(_03392_));
 OAI21x1_ASAP7_75t_R _25780_ (.A1(_03354_),
    .A2(_03335_),
    .B(_03392_),
    .Y(_00106_));
 AOI21x1_ASAP7_75t_R _25781_ (.A1(net6149),
    .A2(net4876),
    .B(net6145),
    .Y(_03393_));
 OAI21x1_ASAP7_75t_R _25782_ (.A1(net4739),
    .A2(_03264_),
    .B(_03393_),
    .Y(_03394_));
 NAND2x1_ASAP7_75t_R _25783_ (.A(net5681),
    .B(_03370_),
    .Y(_03395_));
 AO21x1_ASAP7_75t_R _25784_ (.A1(net5399),
    .A2(net4878),
    .B(net6146),
    .Y(_03396_));
 NAND2x1_ASAP7_75t_R _25785_ (.A(net6153),
    .B(_03236_),
    .Y(_03397_));
 OAI22x1_ASAP7_75t_R _25786_ (.A1(_03395_),
    .A2(_03396_),
    .B1(_03397_),
    .B2(net5681),
    .Y(_03398_));
 OAI21x1_ASAP7_75t_R _25787_ (.A1(_03394_),
    .A2(_03398_),
    .B(net6141),
    .Y(_03399_));
 OA21x2_ASAP7_75t_R _25788_ (.A1(net6153),
    .A2(net4652),
    .B(_03163_),
    .Y(_03400_));
 NAND2x1_ASAP7_75t_R _25789_ (.A(_03347_),
    .B(_03400_),
    .Y(_03401_));
 INVx1_ASAP7_75t_R _25790_ (.A(_03204_),
    .Y(_03402_));
 AO21x1_ASAP7_75t_R _25791_ (.A1(_03128_),
    .A2(_03129_),
    .B(_03359_),
    .Y(_03403_));
 INVx1_ASAP7_75t_R _25792_ (.A(_03403_),
    .Y(_03404_));
 AOI21x1_ASAP7_75t_R _25793_ (.A1(net4740),
    .A2(_03196_),
    .B(_03163_),
    .Y(_03405_));
 OAI21x1_ASAP7_75t_R _25794_ (.A1(_03402_),
    .A2(_03404_),
    .B(_03405_),
    .Y(_03406_));
 AOI21x1_ASAP7_75t_R _25795_ (.A1(_03401_),
    .A2(_03406_),
    .B(net5685),
    .Y(_03407_));
 NOR2x1_ASAP7_75t_R _25796_ (.A(_03399_),
    .B(_03407_),
    .Y(_03408_));
 OAI21x1_ASAP7_75t_R _25797_ (.A1(_03118_),
    .A2(_03341_),
    .B(net6153),
    .Y(_03409_));
 OAI21x1_ASAP7_75t_R _25798_ (.A1(_03226_),
    .A2(_03281_),
    .B(net6147),
    .Y(_03410_));
 AOI21x1_ASAP7_75t_R _25799_ (.A1(_03409_),
    .A2(_03410_),
    .B(net6145),
    .Y(_03411_));
 AOI21x1_ASAP7_75t_R _25800_ (.A1(_03132_),
    .A2(_03279_),
    .B(net5686),
    .Y(_03412_));
 NOR2x1_ASAP7_75t_R _25801_ (.A(_03411_),
    .B(_03412_),
    .Y(_03413_));
 OAI21x1_ASAP7_75t_R _25802_ (.A1(net5689),
    .A2(net6157),
    .B(_03151_),
    .Y(_03414_));
 AO21x1_ASAP7_75t_R _25803_ (.A1(_03414_),
    .A2(_03360_),
    .B(net6153),
    .Y(_03415_));
 AOI21x1_ASAP7_75t_R _25804_ (.A1(_03415_),
    .A2(_03260_),
    .B(net5685),
    .Y(_03416_));
 NAND2x1_ASAP7_75t_R _25805_ (.A(net5681),
    .B(_03350_),
    .Y(_03417_));
 OAI21x1_ASAP7_75t_R _25806_ (.A1(_03416_),
    .A2(_03417_),
    .B(net5679),
    .Y(_03418_));
 AOI21x1_ASAP7_75t_R _25807_ (.A1(net5392),
    .A2(_03413_),
    .B(_03418_),
    .Y(_03419_));
 OAI21x1_ASAP7_75t_R _25808_ (.A1(_03408_),
    .A2(_03419_),
    .B(net6142),
    .Y(_03420_));
 OAI21x1_ASAP7_75t_R _25809_ (.A1(_03275_),
    .A2(_03070_),
    .B(net6149),
    .Y(_03421_));
 OAI21x1_ASAP7_75t_R _25810_ (.A1(net4738),
    .A2(_03259_),
    .B(net6153),
    .Y(_03422_));
 AOI21x1_ASAP7_75t_R _25811_ (.A1(_03421_),
    .A2(_03422_),
    .B(net5683),
    .Y(_03423_));
 OAI21x1_ASAP7_75t_R _25812_ (.A1(net4657),
    .A2(_03236_),
    .B(net6153),
    .Y(_03424_));
 AOI22x1_ASAP7_75t_R _25813_ (.A1(net6156),
    .A2(net5688),
    .B1(net6161),
    .B2(net6160),
    .Y(_03425_));
 AOI22x1_ASAP7_75t_R _25814_ (.A1(net5682),
    .A2(_03072_),
    .B1(net6159),
    .B2(_03007_),
    .Y(_03426_));
 OAI21x1_ASAP7_75t_R _25815_ (.A1(_03425_),
    .A2(_03426_),
    .B(net6149),
    .Y(_03427_));
 AOI21x1_ASAP7_75t_R _25816_ (.A1(_03424_),
    .A2(_03427_),
    .B(net6145),
    .Y(_03428_));
 OAI21x1_ASAP7_75t_R _25817_ (.A1(_03423_),
    .A2(_03428_),
    .B(net5391),
    .Y(_03429_));
 AO21x1_ASAP7_75t_R _25818_ (.A1(net4740),
    .A2(_03414_),
    .B(net6149),
    .Y(_03430_));
 NAND2x1_ASAP7_75t_R _25819_ (.A(_03312_),
    .B(_03204_),
    .Y(_03431_));
 AOI21x1_ASAP7_75t_R _25820_ (.A1(_03430_),
    .A2(_03431_),
    .B(net6144),
    .Y(_03432_));
 INVx1_ASAP7_75t_R _25821_ (.A(_03267_),
    .Y(_03433_));
 OAI21x1_ASAP7_75t_R _25822_ (.A1(_03426_),
    .A2(net5110),
    .B(net6153),
    .Y(_03434_));
 AOI21x1_ASAP7_75t_R _25823_ (.A1(_03433_),
    .A2(_03434_),
    .B(net5683),
    .Y(_03435_));
 OAI21x1_ASAP7_75t_R _25824_ (.A1(_03432_),
    .A2(_03435_),
    .B(net5681),
    .Y(_03436_));
 AOI21x1_ASAP7_75t_R _25825_ (.A1(_03429_),
    .A2(_03436_),
    .B(net6141),
    .Y(_03437_));
 NOR2x1_ASAP7_75t_R _25826_ (.A(_03115_),
    .B(net4556),
    .Y(_03438_));
 NOR2x1_ASAP7_75t_R _25827_ (.A(_03070_),
    .B(_03298_),
    .Y(_03439_));
 OAI21x1_ASAP7_75t_R _25828_ (.A1(_03439_),
    .A2(_03438_),
    .B(net5684),
    .Y(_03440_));
 NAND2x1_ASAP7_75t_R _25829_ (.A(_03186_),
    .B(_03337_),
    .Y(_03441_));
 INVx1_ASAP7_75t_R _25830_ (.A(_03118_),
    .Y(_03442_));
 AOI21x1_ASAP7_75t_R _25831_ (.A1(net5399),
    .A2(net5691),
    .B(net6147),
    .Y(_03443_));
 AOI21x1_ASAP7_75t_R _25832_ (.A1(_03442_),
    .A2(_03443_),
    .B(net5685),
    .Y(_03444_));
 AOI21x1_ASAP7_75t_R _25833_ (.A1(_03441_),
    .A2(_03444_),
    .B(net5681),
    .Y(_03445_));
 NAND2x1_ASAP7_75t_R _25834_ (.A(_03440_),
    .B(_03445_),
    .Y(_03446_));
 NAND2x1_ASAP7_75t_R _25835_ (.A(_03201_),
    .B(_03443_),
    .Y(_03447_));
 AOI21x1_ASAP7_75t_R _25836_ (.A1(net4556),
    .A2(_03447_),
    .B(net6145),
    .Y(_03448_));
 OAI21x1_ASAP7_75t_R _25837_ (.A1(_03118_),
    .A2(_03256_),
    .B(net6150),
    .Y(_03449_));
 AOI21x1_ASAP7_75t_R _25838_ (.A1(_03434_),
    .A2(_03449_),
    .B(net5683),
    .Y(_03450_));
 OAI21x1_ASAP7_75t_R _25839_ (.A1(_03448_),
    .A2(_03450_),
    .B(net5681),
    .Y(_03451_));
 AOI21x1_ASAP7_75t_R _25840_ (.A1(_03446_),
    .A2(_03451_),
    .B(net5679),
    .Y(_03452_));
 OAI21x1_ASAP7_75t_R _25841_ (.A1(_03437_),
    .A2(_03452_),
    .B(net5680),
    .Y(_03453_));
 NAND2x1_ASAP7_75t_R _25842_ (.A(_03420_),
    .B(_03453_),
    .Y(_00107_));
 OA21x2_ASAP7_75t_R _25843_ (.A1(_03320_),
    .A2(_03257_),
    .B(net5681),
    .Y(_03454_));
 NAND2x1_ASAP7_75t_R _25844_ (.A(net5694),
    .B(net5402),
    .Y(_03455_));
 AOI21x1_ASAP7_75t_R _25845_ (.A1(_03455_),
    .A2(_03312_),
    .B(net6151),
    .Y(_03456_));
 NOR2x1_ASAP7_75t_R _25846_ (.A(_03075_),
    .B(_03319_),
    .Y(_03457_));
 OAI21x1_ASAP7_75t_R _25847_ (.A1(_03456_),
    .A2(_03457_),
    .B(net5687),
    .Y(_03458_));
 AOI21x1_ASAP7_75t_R _25848_ (.A1(net5054),
    .A2(net5400),
    .B(net6155),
    .Y(_03459_));
 OAI21x1_ASAP7_75t_R _25849_ (.A1(net4876),
    .A2(net4873),
    .B(net5687),
    .Y(_03460_));
 NOR2x1_ASAP7_75t_R _25850_ (.A(_03268_),
    .B(_03269_),
    .Y(_03461_));
 NOR2x1_ASAP7_75t_R _25851_ (.A(_03256_),
    .B(_03219_),
    .Y(_03462_));
 OAI21x1_ASAP7_75t_R _25852_ (.A1(_03461_),
    .A2(_03462_),
    .B(net6144),
    .Y(_03463_));
 AOI21x1_ASAP7_75t_R _25853_ (.A1(_03460_),
    .A2(_03463_),
    .B(net5681),
    .Y(_03464_));
 AOI211x1_ASAP7_75t_R _25854_ (.A1(_03454_),
    .A2(_03458_),
    .B(_03464_),
    .C(net6141),
    .Y(_03465_));
 NAND2x1_ASAP7_75t_R _25855_ (.A(_03105_),
    .B(_03150_),
    .Y(_03466_));
 AND3x1_ASAP7_75t_R _25856_ (.A(_03376_),
    .B(_03466_),
    .C(net5686),
    .Y(_03467_));
 NAND2x1_ASAP7_75t_R _25857_ (.A(net6143),
    .B(_03140_),
    .Y(_03468_));
 AND3x1_ASAP7_75t_R _25858_ (.A(_03105_),
    .B(net6148),
    .C(_03130_),
    .Y(_03469_));
 OAI21x1_ASAP7_75t_R _25859_ (.A1(_03468_),
    .A2(_03469_),
    .B(net5681),
    .Y(_03470_));
 OAI21x1_ASAP7_75t_R _25860_ (.A1(net4738),
    .A2(_03226_),
    .B(net6147),
    .Y(_03471_));
 AOI21x1_ASAP7_75t_R _25861_ (.A1(_03471_),
    .A2(_03336_),
    .B(net6145),
    .Y(_03472_));
 AO21x1_ASAP7_75t_R _25862_ (.A1(_03139_),
    .A2(_03414_),
    .B(net6153),
    .Y(_03473_));
 AOI21x1_ASAP7_75t_R _25863_ (.A1(net5049),
    .A2(net5396),
    .B(net6152),
    .Y(_03474_));
 NAND2x1_ASAP7_75t_R _25864_ (.A(net4739),
    .B(_03474_),
    .Y(_03475_));
 AOI21x1_ASAP7_75t_R _25865_ (.A1(_03473_),
    .A2(_03475_),
    .B(net5685),
    .Y(_03476_));
 OAI21x1_ASAP7_75t_R _25866_ (.A1(_03472_),
    .A2(_03476_),
    .B(net5392),
    .Y(_03477_));
 OAI21x1_ASAP7_75t_R _25867_ (.A1(_03467_),
    .A2(_03470_),
    .B(_03477_),
    .Y(_03478_));
 OAI21x1_ASAP7_75t_R _25868_ (.A1(net5679),
    .A2(_03478_),
    .B(net5680),
    .Y(_03479_));
 AOI21x1_ASAP7_75t_R _25869_ (.A1(net5397),
    .A2(net5402),
    .B(net6151),
    .Y(_03480_));
 NOR2x1_ASAP7_75t_R _25870_ (.A(net6154),
    .B(net5397),
    .Y(_03481_));
 AOI21x1_ASAP7_75t_R _25871_ (.A1(net4650),
    .A2(_03480_),
    .B(_03481_),
    .Y(_03482_));
 AOI21x1_ASAP7_75t_R _25872_ (.A1(net6144),
    .A2(_03482_),
    .B(net6141),
    .Y(_03483_));
 AO21x1_ASAP7_75t_R _25873_ (.A1(_03105_),
    .A2(_03114_),
    .B(net6148),
    .Y(_03484_));
 NAND2x1_ASAP7_75t_R _25874_ (.A(_03254_),
    .B(_03484_),
    .Y(_03485_));
 AO21x1_ASAP7_75t_R _25875_ (.A1(_03483_),
    .A2(_03485_),
    .B(net5394),
    .Y(_03486_));
 OAI21x1_ASAP7_75t_R _25876_ (.A1(_03211_),
    .A2(_03058_),
    .B(net6144),
    .Y(_03487_));
 INVx1_ASAP7_75t_R _25877_ (.A(_03456_),
    .Y(_03488_));
 NAND2x1_ASAP7_75t_R _25878_ (.A(net5397),
    .B(net5402),
    .Y(_03489_));
 NAND2x1_ASAP7_75t_R _25879_ (.A(_03489_),
    .B(net4873),
    .Y(_03490_));
 AO21x1_ASAP7_75t_R _25880_ (.A1(_03488_),
    .A2(_03490_),
    .B(net6144),
    .Y(_03491_));
 AOI21x1_ASAP7_75t_R _25881_ (.A1(_03487_),
    .A2(_03491_),
    .B(_03208_),
    .Y(_03492_));
 OA21x2_ASAP7_75t_R _25882_ (.A1(_03310_),
    .A2(net6148),
    .B(net6144),
    .Y(_03493_));
 AOI21x1_ASAP7_75t_R _25883_ (.A1(_03493_),
    .A2(_03323_),
    .B(net5679),
    .Y(_03494_));
 NAND2x1_ASAP7_75t_R _25884_ (.A(_03312_),
    .B(_03459_),
    .Y(_03495_));
 NAND2x1_ASAP7_75t_R _25885_ (.A(_03158_),
    .B(_03495_),
    .Y(_03496_));
 AOI21x1_ASAP7_75t_R _25886_ (.A1(_03494_),
    .A2(_03496_),
    .B(net5681),
    .Y(_03497_));
 AND2x2_ASAP7_75t_R _25887_ (.A(_03282_),
    .B(_03216_),
    .Y(_03498_));
 AOI21x1_ASAP7_75t_R _25888_ (.A1(net6152),
    .A2(_03077_),
    .B(net6144),
    .Y(_03499_));
 AOI21x1_ASAP7_75t_R _25889_ (.A1(_03234_),
    .A2(_03499_),
    .B(net6141),
    .Y(_03500_));
 OAI21x1_ASAP7_75t_R _25890_ (.A1(_03183_),
    .A2(_03498_),
    .B(_03500_),
    .Y(_03501_));
 AOI21x1_ASAP7_75t_R _25891_ (.A1(_03501_),
    .A2(_03497_),
    .B(net5680),
    .Y(_03502_));
 OAI21x1_ASAP7_75t_R _25892_ (.A1(_03486_),
    .A2(_03492_),
    .B(_03502_),
    .Y(_03503_));
 OAI21x1_ASAP7_75t_R _25893_ (.A1(_03465_),
    .A2(_03479_),
    .B(_03503_),
    .Y(_00108_));
 OAI21x1_ASAP7_75t_R _25894_ (.A1(_03275_),
    .A2(_03282_),
    .B(net5685),
    .Y(_03504_));
 NAND2x1_ASAP7_75t_R _25895_ (.A(net5681),
    .B(_03504_),
    .Y(_03505_));
 NAND2x1_ASAP7_75t_R _25896_ (.A(net6153),
    .B(net4740),
    .Y(_03506_));
 AOI21x1_ASAP7_75t_R _25897_ (.A1(_03506_),
    .A2(_03410_),
    .B(net5685),
    .Y(_03507_));
 OAI21x1_ASAP7_75t_R _25898_ (.A1(_03505_),
    .A2(_03507_),
    .B(net5679),
    .Y(_03508_));
 AOI21x1_ASAP7_75t_R _25899_ (.A1(_03138_),
    .A2(_03360_),
    .B(net6153),
    .Y(_03509_));
 AOI21x1_ASAP7_75t_R _25900_ (.A1(_03139_),
    .A2(_03414_),
    .B(net6146),
    .Y(_03510_));
 OAI21x1_ASAP7_75t_R _25901_ (.A1(_03509_),
    .A2(_03510_),
    .B(net5685),
    .Y(_03511_));
 NAND2x1_ASAP7_75t_R _25902_ (.A(_03163_),
    .B(_03511_),
    .Y(_03512_));
 NAND2x1_ASAP7_75t_R _25903_ (.A(_03375_),
    .B(_03197_),
    .Y(_03513_));
 INVx1_ASAP7_75t_R _25904_ (.A(_03177_),
    .Y(_03514_));
 AOI21x1_ASAP7_75t_R _25905_ (.A1(_03513_),
    .A2(_03514_),
    .B(_03066_),
    .Y(_03515_));
 NOR2x1_ASAP7_75t_R _25906_ (.A(_03512_),
    .B(_03515_),
    .Y(_03516_));
 OAI21x1_ASAP7_75t_R _25907_ (.A1(_03508_),
    .A2(_03516_),
    .B(net5680),
    .Y(_03517_));
 NAND2x1_ASAP7_75t_R _25908_ (.A(net6147),
    .B(net4738),
    .Y(_03518_));
 AO21x1_ASAP7_75t_R _25909_ (.A1(_03312_),
    .A2(_03134_),
    .B(net6147),
    .Y(_03519_));
 NAND2x1_ASAP7_75t_R _25910_ (.A(_03518_),
    .B(_03519_),
    .Y(_03520_));
 NOR2x1_ASAP7_75t_R _25911_ (.A(_03075_),
    .B(_03228_),
    .Y(_03521_));
 OAI21x1_ASAP7_75t_R _25912_ (.A1(net6147),
    .A2(_03341_),
    .B(net6143),
    .Y(_03522_));
 OAI21x1_ASAP7_75t_R _25913_ (.A1(_03521_),
    .A2(_03522_),
    .B(net5681),
    .Y(_03523_));
 AOI21x1_ASAP7_75t_R _25914_ (.A1(net5685),
    .A2(_03520_),
    .B(_03523_),
    .Y(_03524_));
 AO21x1_ASAP7_75t_R _25915_ (.A1(net5690),
    .A2(net6151),
    .B(net5687),
    .Y(_03525_));
 OAI21x1_ASAP7_75t_R _25916_ (.A1(_03525_),
    .A2(_03456_),
    .B(net5394),
    .Y(_03526_));
 OA21x2_ASAP7_75t_R _25917_ (.A1(_03218_),
    .A2(_03179_),
    .B(net6151),
    .Y(_03527_));
 AO21x1_ASAP7_75t_R _25918_ (.A1(_03196_),
    .A2(_03455_),
    .B(net6144),
    .Y(_03528_));
 NOR2x1_ASAP7_75t_R _25919_ (.A(_03527_),
    .B(_03528_),
    .Y(_03529_));
 OAI21x1_ASAP7_75t_R _25920_ (.A1(_03526_),
    .A2(_03529_),
    .B(net6141),
    .Y(_03530_));
 NOR2x1_ASAP7_75t_R _25921_ (.A(_03524_),
    .B(_03530_),
    .Y(_03531_));
 NOR2x1_ASAP7_75t_R _25922_ (.A(_03517_),
    .B(_03531_),
    .Y(_03532_));
 NOR2x1_ASAP7_75t_R _25923_ (.A(net4878),
    .B(net6155),
    .Y(_03533_));
 AOI21x1_ASAP7_75t_R _25924_ (.A1(net6155),
    .A2(net4875),
    .B(_03533_),
    .Y(_03534_));
 OAI21x1_ASAP7_75t_R _25925_ (.A1(net5686),
    .A2(_03534_),
    .B(net5681),
    .Y(_03535_));
 OAI21x1_ASAP7_75t_R _25926_ (.A1(net4656),
    .A2(_03118_),
    .B(net6146),
    .Y(_03536_));
 OAI21x1_ASAP7_75t_R _25927_ (.A1(_03236_),
    .A2(_03341_),
    .B(net6153),
    .Y(_03537_));
 AOI21x1_ASAP7_75t_R _25928_ (.A1(_03536_),
    .A2(_03537_),
    .B(net6144),
    .Y(_03538_));
 NOR2x1_ASAP7_75t_R _25929_ (.A(_03535_),
    .B(_03538_),
    .Y(_03539_));
 OA21x2_ASAP7_75t_R _25930_ (.A1(net4655),
    .A2(net6150),
    .B(net5686),
    .Y(_03540_));
 NAND2x1_ASAP7_75t_R _25931_ (.A(_03402_),
    .B(_03540_),
    .Y(_03541_));
 AOI21x1_ASAP7_75t_R _25932_ (.A1(net6146),
    .A2(_03403_),
    .B(net5686),
    .Y(_03542_));
 OAI21x1_ASAP7_75t_R _25933_ (.A1(net4653),
    .A2(_03387_),
    .B(_03542_),
    .Y(_03543_));
 AOI21x1_ASAP7_75t_R _25934_ (.A1(_03541_),
    .A2(_03543_),
    .B(net5681),
    .Y(_03544_));
 OAI21x1_ASAP7_75t_R _25935_ (.A1(_03539_),
    .A2(_03544_),
    .B(net6141),
    .Y(_03545_));
 NAND2x1_ASAP7_75t_R _25936_ (.A(_03312_),
    .B(_03346_),
    .Y(_03546_));
 NAND2x1_ASAP7_75t_R _25937_ (.A(net4740),
    .B(_03267_),
    .Y(_03547_));
 AND3x1_ASAP7_75t_R _25938_ (.A(_03546_),
    .B(_03547_),
    .C(net5686),
    .Y(_03548_));
 NAND2x1_ASAP7_75t_R _25939_ (.A(net6151),
    .B(net5402),
    .Y(_03549_));
 OA21x2_ASAP7_75t_R _25940_ (.A1(_03052_),
    .A2(net5111),
    .B(_03549_),
    .Y(_03550_));
 AO21x1_ASAP7_75t_R _25941_ (.A1(_03550_),
    .A2(net6144),
    .B(net5681),
    .Y(_03551_));
 AOI21x1_ASAP7_75t_R _25942_ (.A1(net6148),
    .A2(net4656),
    .B(net6144),
    .Y(_03552_));
 OAI21x1_ASAP7_75t_R _25943_ (.A1(_03259_),
    .A2(_03341_),
    .B(net6153),
    .Y(_03553_));
 AOI21x1_ASAP7_75t_R _25944_ (.A1(_03552_),
    .A2(_03553_),
    .B(net5393),
    .Y(_03554_));
 AO21x1_ASAP7_75t_R _25945_ (.A1(_03489_),
    .A2(net4655),
    .B(net6148),
    .Y(_03555_));
 NAND2x1_ASAP7_75t_R _25946_ (.A(_03224_),
    .B(_03555_),
    .Y(_03556_));
 AOI21x1_ASAP7_75t_R _25947_ (.A1(_03554_),
    .A2(_03556_),
    .B(net6141),
    .Y(_03557_));
 OAI21x1_ASAP7_75t_R _25948_ (.A1(_03548_),
    .A2(_03551_),
    .B(_03557_),
    .Y(_03558_));
 AOI21x1_ASAP7_75t_R _25949_ (.A1(_03545_),
    .A2(_03558_),
    .B(net5680),
    .Y(_03559_));
 NOR2x1_ASAP7_75t_R _25950_ (.A(_03532_),
    .B(_03559_),
    .Y(_00109_));
 AND3x1_ASAP7_75t_R _25951_ (.A(_03403_),
    .B(_03216_),
    .C(net6153),
    .Y(_03560_));
 AO21x1_ASAP7_75t_R _25952_ (.A1(_03150_),
    .A2(_03247_),
    .B(net5685),
    .Y(_03561_));
 AOI21x1_ASAP7_75t_R _25953_ (.A1(net6153),
    .A2(net4657),
    .B(net6145),
    .Y(_03562_));
 INVx1_ASAP7_75t_R _25954_ (.A(_03139_),
    .Y(_03563_));
 NOR2x1_ASAP7_75t_R _25955_ (.A(net5693),
    .B(net5396),
    .Y(_03564_));
 OAI21x1_ASAP7_75t_R _25956_ (.A1(_03563_),
    .A2(_03564_),
    .B(net6150),
    .Y(_03565_));
 AOI21x1_ASAP7_75t_R _25957_ (.A1(_03562_),
    .A2(_03565_),
    .B(net5391),
    .Y(_03566_));
 OAI21x1_ASAP7_75t_R _25958_ (.A1(_03560_),
    .A2(_03561_),
    .B(_03566_),
    .Y(_03567_));
 AO21x1_ASAP7_75t_R _25959_ (.A1(_03236_),
    .A2(net6153),
    .B(net6145),
    .Y(_03568_));
 NOR2x1_ASAP7_75t_R _25960_ (.A(_03367_),
    .B(_03568_),
    .Y(_03569_));
 AO21x1_ASAP7_75t_R _25961_ (.A1(net4740),
    .A2(_03134_),
    .B(net6150),
    .Y(_03570_));
 NAND2x1_ASAP7_75t_R _25962_ (.A(_03312_),
    .B(_03267_),
    .Y(_03571_));
 AOI21x1_ASAP7_75t_R _25963_ (.A1(_03570_),
    .A2(_03571_),
    .B(net5684),
    .Y(_03572_));
 OAI21x1_ASAP7_75t_R _25964_ (.A1(_03572_),
    .A2(_03569_),
    .B(net5392),
    .Y(_03573_));
 AOI21x1_ASAP7_75t_R _25965_ (.A1(_03573_),
    .A2(_03567_),
    .B(net5679),
    .Y(_03574_));
 NAND2x1p5_ASAP7_75t_R _25966_ (.A(_03216_),
    .B(_03480_),
    .Y(_03575_));
 OAI21x1_ASAP7_75t_R _25967_ (.A1(net6153),
    .A2(net4652),
    .B(net5683),
    .Y(_03576_));
 NOR3x1_ASAP7_75t_R _25968_ (.A(net5396),
    .B(net6153),
    .C(net4874),
    .Y(_03577_));
 NOR2x1_ASAP7_75t_R _25969_ (.A(_03576_),
    .B(_03577_),
    .Y(_03578_));
 NAND2x1_ASAP7_75t_R _25970_ (.A(_03575_),
    .B(_03578_),
    .Y(_03579_));
 OAI21x1_ASAP7_75t_R _25971_ (.A1(net4876),
    .A2(_03237_),
    .B(net6149),
    .Y(_03580_));
 AOI21x1_ASAP7_75t_R _25972_ (.A1(_03186_),
    .A2(_03346_),
    .B(net5686),
    .Y(_03581_));
 AOI21x1_ASAP7_75t_R _25973_ (.A1(_03580_),
    .A2(_03581_),
    .B(net5391),
    .Y(_03582_));
 NAND2x1_ASAP7_75t_R _25974_ (.A(_03579_),
    .B(_03582_),
    .Y(_03583_));
 AO21x1_ASAP7_75t_R _25975_ (.A1(net4652),
    .A2(_03134_),
    .B(net6153),
    .Y(_03584_));
 AOI21x1_ASAP7_75t_R _25976_ (.A1(_03355_),
    .A2(_03584_),
    .B(net6145),
    .Y(_03585_));
 AO21x1_ASAP7_75t_R _25977_ (.A1(_01266_),
    .A2(_01270_),
    .B(net6150),
    .Y(_03586_));
 NOR2x1_ASAP7_75t_R _25978_ (.A(net5395),
    .B(net5691),
    .Y(_03587_));
 OAI21x1_ASAP7_75t_R _25979_ (.A1(_03190_),
    .A2(_03587_),
    .B(net6149),
    .Y(_03588_));
 AOI21x1_ASAP7_75t_R _25980_ (.A1(_03586_),
    .A2(_03588_),
    .B(net5684),
    .Y(_03589_));
 OAI21x1_ASAP7_75t_R _25981_ (.A1(_03585_),
    .A2(_03589_),
    .B(net5392),
    .Y(_03590_));
 AOI21x1_ASAP7_75t_R _25982_ (.A1(_03583_),
    .A2(_03590_),
    .B(net6141),
    .Y(_03591_));
 OAI21x1_ASAP7_75t_R _25983_ (.A1(_03574_),
    .A2(_03591_),
    .B(net5680),
    .Y(_03592_));
 AND3x1_ASAP7_75t_R _25984_ (.A(_03442_),
    .B(net6147),
    .C(_03375_),
    .Y(_03593_));
 AOI21x1_ASAP7_75t_R _25985_ (.A1(_01267_),
    .A2(net6147),
    .B(net5685),
    .Y(_03594_));
 AOI21x1_ASAP7_75t_R _25986_ (.A1(_03594_),
    .A2(_03546_),
    .B(net5681),
    .Y(_03595_));
 OAI21x1_ASAP7_75t_R _25987_ (.A1(_03248_),
    .A2(_03593_),
    .B(_03595_),
    .Y(_03596_));
 INVx1_ASAP7_75t_R _25988_ (.A(_03379_),
    .Y(_03597_));
 AOI21x1_ASAP7_75t_R _25989_ (.A1(_03396_),
    .A2(_03495_),
    .B(net6144),
    .Y(_03598_));
 OAI21x1_ASAP7_75t_R _25990_ (.A1(_03597_),
    .A2(_03598_),
    .B(net5681),
    .Y(_03599_));
 AOI21x1_ASAP7_75t_R _25991_ (.A1(_03596_),
    .A2(_03599_),
    .B(net5679),
    .Y(_03600_));
 AOI21x1_ASAP7_75t_R _25992_ (.A1(_03288_),
    .A2(_03203_),
    .B(net6145),
    .Y(_03601_));
 NAND2x1_ASAP7_75t_R _25993_ (.A(net6153),
    .B(_03118_),
    .Y(_03602_));
 AOI21x1_ASAP7_75t_R _25994_ (.A1(_03602_),
    .A2(_03410_),
    .B(net5685),
    .Y(_03603_));
 OAI21x1_ASAP7_75t_R _25995_ (.A1(_03601_),
    .A2(_03603_),
    .B(net5681),
    .Y(_03604_));
 NAND2x1_ASAP7_75t_R _25996_ (.A(_03247_),
    .B(_03474_),
    .Y(_03605_));
 OAI21x1_ASAP7_75t_R _25997_ (.A1(_03425_),
    .A2(_03054_),
    .B(net6149),
    .Y(_03606_));
 AOI21x1_ASAP7_75t_R _25998_ (.A1(_03605_),
    .A2(_03606_),
    .B(net6144),
    .Y(_03607_));
 OAI21x1_ASAP7_75t_R _25999_ (.A1(_03275_),
    .A2(_03190_),
    .B(net6153),
    .Y(_03608_));
 OAI21x1_ASAP7_75t_R _26000_ (.A1(_03426_),
    .A2(net5110),
    .B(net6149),
    .Y(_03609_));
 AOI21x1_ASAP7_75t_R _26001_ (.A1(_03608_),
    .A2(_03609_),
    .B(net5683),
    .Y(_03610_));
 OAI21x1_ASAP7_75t_R _26002_ (.A1(_03607_),
    .A2(_03610_),
    .B(net5391),
    .Y(_03611_));
 AOI21x1_ASAP7_75t_R _26003_ (.A1(_03604_),
    .A2(_03611_),
    .B(net6141),
    .Y(_03612_));
 OAI21x1_ASAP7_75t_R _26004_ (.A1(_03600_),
    .A2(_03612_),
    .B(net6142),
    .Y(_03613_));
 NAND2x1_ASAP7_75t_R _26005_ (.A(_03613_),
    .B(_03592_),
    .Y(_00110_));
 NAND2x1_ASAP7_75t_R _26006_ (.A(net4740),
    .B(_03196_),
    .Y(_03614_));
 AND3x1_ASAP7_75t_R _26007_ (.A(_03614_),
    .B(_03292_),
    .C(net5687),
    .Y(_03615_));
 AO21x1_ASAP7_75t_R _26008_ (.A1(_03331_),
    .A2(_03581_),
    .B(net5394),
    .Y(_03616_));
 NOR2x1_ASAP7_75t_R _26009_ (.A(net5686),
    .B(_03474_),
    .Y(_03617_));
 AOI21x1_ASAP7_75t_R _26010_ (.A1(_03495_),
    .A2(_03617_),
    .B(net5681),
    .Y(_03618_));
 AO21x1_ASAP7_75t_R _26011_ (.A1(net5400),
    .A2(_03310_),
    .B(net6155),
    .Y(_03619_));
 AOI21x1_ASAP7_75t_R _26012_ (.A1(_03327_),
    .A2(_03196_),
    .B(net6144),
    .Y(_03620_));
 OAI21x1_ASAP7_75t_R _26013_ (.A1(_03250_),
    .A2(_03619_),
    .B(_03620_),
    .Y(_03621_));
 AOI21x1_ASAP7_75t_R _26014_ (.A1(_03618_),
    .A2(_03621_),
    .B(net6141),
    .Y(_03622_));
 OAI21x1_ASAP7_75t_R _26015_ (.A1(_03616_),
    .A2(_03615_),
    .B(_03622_),
    .Y(_03623_));
 OAI21x1_ASAP7_75t_R _26016_ (.A1(_03236_),
    .A2(_03237_),
    .B(net6153),
    .Y(_03624_));
 NOR2x1_ASAP7_75t_R _26017_ (.A(net6144),
    .B(_03150_),
    .Y(_03625_));
 NAND2x1_ASAP7_75t_R _26018_ (.A(_03624_),
    .B(_03625_),
    .Y(_03626_));
 NAND2x1_ASAP7_75t_R _26019_ (.A(net6147),
    .B(_03259_),
    .Y(_03627_));
 OA21x2_ASAP7_75t_R _26020_ (.A1(net4740),
    .A2(net6147),
    .B(net6144),
    .Y(_03628_));
 AOI21x1_ASAP7_75t_R _26021_ (.A1(_03627_),
    .A2(_03628_),
    .B(net5393),
    .Y(_03629_));
 AOI21x1_ASAP7_75t_R _26022_ (.A1(_03626_),
    .A2(_03629_),
    .B(net5679),
    .Y(_03630_));
 AND3x1_ASAP7_75t_R _26023_ (.A(_03312_),
    .B(net6154),
    .C(_03077_),
    .Y(_03631_));
 NAND2x1_ASAP7_75t_R _26024_ (.A(net6155),
    .B(net5395),
    .Y(_03632_));
 OAI21x1_ASAP7_75t_R _26025_ (.A1(_03256_),
    .A2(_03219_),
    .B(_03632_),
    .Y(_03633_));
 AOI21x1_ASAP7_75t_R _26026_ (.A1(net5687),
    .A2(_03633_),
    .B(net5681),
    .Y(_03634_));
 OAI21x1_ASAP7_75t_R _26027_ (.A1(_03320_),
    .A2(_03631_),
    .B(_03634_),
    .Y(_03635_));
 AOI21x1_ASAP7_75t_R _26028_ (.A1(_03630_),
    .A2(_03635_),
    .B(net5680),
    .Y(_03636_));
 NAND2x1_ASAP7_75t_R _26029_ (.A(_03636_),
    .B(_03623_),
    .Y(_03637_));
 OAI21x1_ASAP7_75t_R _26030_ (.A1(_03310_),
    .A2(net6153),
    .B(_03136_),
    .Y(_03638_));
 AO21x1_ASAP7_75t_R _26031_ (.A1(_03105_),
    .A2(_03139_),
    .B(net6148),
    .Y(_03639_));
 NAND2x1_ASAP7_75t_R _26032_ (.A(_03254_),
    .B(_03639_),
    .Y(_03640_));
 AOI21x1_ASAP7_75t_R _26033_ (.A1(_03638_),
    .A2(_03640_),
    .B(net5681),
    .Y(_03641_));
 OR2x2_ASAP7_75t_R _26034_ (.A(_01270_),
    .B(net6153),
    .Y(_03642_));
 AO21x1_ASAP7_75t_R _26035_ (.A1(net4739),
    .A2(net4652),
    .B(net6150),
    .Y(_03643_));
 AOI21x1_ASAP7_75t_R _26036_ (.A1(_03642_),
    .A2(_03643_),
    .B(net5684),
    .Y(_03644_));
 INVx1_ASAP7_75t_R _26037_ (.A(_03370_),
    .Y(_03645_));
 NOR2x1_ASAP7_75t_R _26038_ (.A(_03645_),
    .B(_03298_),
    .Y(_03646_));
 OAI21x1_ASAP7_75t_R _26039_ (.A1(net4738),
    .A2(_03228_),
    .B(net5684),
    .Y(_03647_));
 OAI21x1_ASAP7_75t_R _26040_ (.A1(_03646_),
    .A2(_03647_),
    .B(net5681),
    .Y(_03648_));
 OAI21x1_ASAP7_75t_R _26041_ (.A1(_03644_),
    .A2(_03648_),
    .B(net6141),
    .Y(_03649_));
 NOR2x1_ASAP7_75t_R _26042_ (.A(_03641_),
    .B(_03649_),
    .Y(_03650_));
 NAND2x1_ASAP7_75t_R _26043_ (.A(_03077_),
    .B(_03215_),
    .Y(_03651_));
 AOI21x1_ASAP7_75t_R _26044_ (.A1(_03415_),
    .A2(_03651_),
    .B(net6145),
    .Y(_03652_));
 AOI21x1_ASAP7_75t_R _26045_ (.A1(_03077_),
    .A2(_03130_),
    .B(net6148),
    .Y(_03653_));
 OAI21x1_ASAP7_75t_R _26046_ (.A1(net4656),
    .A2(_03228_),
    .B(net6144),
    .Y(_03654_));
 NOR2x1_ASAP7_75t_R _26047_ (.A(_03653_),
    .B(_03654_),
    .Y(_03655_));
 OAI21x1_ASAP7_75t_R _26048_ (.A1(_03652_),
    .A2(_03655_),
    .B(net5392),
    .Y(_03656_));
 AO21x1_ASAP7_75t_R _26049_ (.A1(_03114_),
    .A2(_03134_),
    .B(net6150),
    .Y(_03657_));
 OAI21x1_ASAP7_75t_R _26050_ (.A1(_03115_),
    .A2(_03564_),
    .B(net6150),
    .Y(_03658_));
 AOI21x1_ASAP7_75t_R _26051_ (.A1(_03657_),
    .A2(_03658_),
    .B(net5684),
    .Y(_03659_));
 AOI21x1_ASAP7_75t_R _26052_ (.A1(_03307_),
    .A2(_03588_),
    .B(net6145),
    .Y(_03660_));
 OAI21x1_ASAP7_75t_R _26053_ (.A1(_03659_),
    .A2(_03660_),
    .B(net5681),
    .Y(_03661_));
 AOI21x1_ASAP7_75t_R _26054_ (.A1(_03656_),
    .A2(_03661_),
    .B(net6141),
    .Y(_03662_));
 OAI21x1_ASAP7_75t_R _26055_ (.A1(_03650_),
    .A2(_03662_),
    .B(net5680),
    .Y(_03663_));
 NAND2x1_ASAP7_75t_R _26056_ (.A(_03663_),
    .B(_03637_),
    .Y(_00111_));
 NOR2x1_ASAP7_75t_R _26057_ (.A(net6654),
    .B(_00474_),
    .Y(_03664_));
 XOR2x2_ASAP7_75t_R _26058_ (.A(_00694_),
    .B(_00687_),
    .Y(_03665_));
 XOR2x2_ASAP7_75t_R _26059_ (.A(_03665_),
    .B(net6436),
    .Y(_03666_));
 XOR2x2_ASAP7_75t_R _26060_ (.A(net6430),
    .B(net6410),
    .Y(_03667_));
 NAND2x1_ASAP7_75t_R _26061_ (.A(_03666_),
    .B(_03667_),
    .Y(_03668_));
 XOR2x2_ASAP7_75t_R _26062_ (.A(_03665_),
    .B(net6552),
    .Y(_03669_));
 XOR2x2_ASAP7_75t_R _26063_ (.A(_12160_),
    .B(net6410),
    .Y(_03670_));
 NAND2x1_ASAP7_75t_R _26064_ (.A(_03669_),
    .B(_03670_),
    .Y(_03671_));
 AOI21x1_ASAP7_75t_R _26065_ (.A1(_03668_),
    .A2(_03671_),
    .B(net6454),
    .Y(_03672_));
 OAI21x1_ASAP7_75t_R _26066_ (.A1(_03664_),
    .A2(net6350),
    .B(net6478),
    .Y(_03673_));
 AND2x2_ASAP7_75t_R _26067_ (.A(net6454),
    .B(_00474_),
    .Y(_03674_));
 NAND2x1_ASAP7_75t_R _26068_ (.A(_03669_),
    .B(_03667_),
    .Y(_03675_));
 NAND2x1_ASAP7_75t_R _26069_ (.A(_03666_),
    .B(_03670_),
    .Y(_03676_));
 AOI21x1_ASAP7_75t_R _26070_ (.A1(_03675_),
    .A2(_03676_),
    .B(net6454),
    .Y(_03677_));
 INVx1_ASAP7_75t_R _26071_ (.A(net6478),
    .Y(_03678_));
 OAI21x1_ASAP7_75t_R _26072_ (.A1(_03674_),
    .A2(net6349),
    .B(_03678_),
    .Y(_03679_));
 NAND2x2_ASAP7_75t_R _26073_ (.A(_03673_),
    .B(_03679_),
    .Y(_01283_));
 NOR2x1_ASAP7_75t_R _26074_ (.A(net6657),
    .B(_00475_),
    .Y(_03680_));
 XOR2x2_ASAP7_75t_R _26075_ (.A(net6612),
    .B(net6580),
    .Y(_03681_));
 XOR2x2_ASAP7_75t_R _26076_ (.A(_03681_),
    .B(net6638),
    .Y(_03682_));
 NAND2x1_ASAP7_75t_R _26077_ (.A(_03665_),
    .B(_03682_),
    .Y(_03683_));
 NOR2x1_ASAP7_75t_R _26078_ (.A(_03665_),
    .B(_03682_),
    .Y(_03684_));
 INVx1_ASAP7_75t_R _26079_ (.A(_03684_),
    .Y(_03685_));
 AOI21x1_ASAP7_75t_R _26080_ (.A1(_03683_),
    .A2(_03685_),
    .B(net6454),
    .Y(_03686_));
 OAI21x1_ASAP7_75t_R _26081_ (.A1(net6398),
    .A2(_03686_),
    .B(net6479),
    .Y(_03687_));
 INVx1_ASAP7_75t_R _26082_ (.A(_03665_),
    .Y(_03688_));
 XOR2x2_ASAP7_75t_R _26083_ (.A(_03681_),
    .B(net6408),
    .Y(_03689_));
 NOR2x1_ASAP7_75t_R _26084_ (.A(_03688_),
    .B(_03689_),
    .Y(_03690_));
 OAI21x1_ASAP7_75t_R _26085_ (.A1(_03690_),
    .A2(_03684_),
    .B(net6654),
    .Y(_03691_));
 INVx1_ASAP7_75t_R _26086_ (.A(net6479),
    .Y(_03692_));
 INVx1_ASAP7_75t_R _26087_ (.A(_03680_),
    .Y(_03693_));
 NAND3x1_ASAP7_75t_R _26088_ (.A(_03691_),
    .B(_03692_),
    .C(net6386),
    .Y(_03694_));
 NAND2x1_ASAP7_75t_R _26089_ (.A(_03687_),
    .B(_03694_),
    .Y(_01280_));
 NOR2x1_ASAP7_75t_R _26090_ (.A(net6656),
    .B(_00476_),
    .Y(_03695_));
 INVx1_ASAP7_75t_R _26091_ (.A(_03695_),
    .Y(_03696_));
 XOR2x2_ASAP7_75t_R _26092_ (.A(_00593_),
    .B(net6610),
    .Y(_03697_));
 XOR2x2_ASAP7_75t_R _26093_ (.A(net6411),
    .B(net6551),
    .Y(_03698_));
 NOR2x1_ASAP7_75t_R _26094_ (.A(_03697_),
    .B(_03698_),
    .Y(_03699_));
 INVx1_ASAP7_75t_R _26095_ (.A(net6551),
    .Y(_03700_));
 NOR2x1_ASAP7_75t_R _26096_ (.A(_03700_),
    .B(net6411),
    .Y(_03701_));
 AND2x2_ASAP7_75t_R _26097_ (.A(net6411),
    .B(_03700_),
    .Y(_03702_));
 OAI21x1_ASAP7_75t_R _26098_ (.A1(_03701_),
    .A2(_03702_),
    .B(_03697_),
    .Y(_03703_));
 INVx1_ASAP7_75t_R _26099_ (.A(_03703_),
    .Y(_03704_));
 OAI21x1_ASAP7_75t_R _26100_ (.A1(_03699_),
    .A2(_03704_),
    .B(net6656),
    .Y(_03705_));
 AOI21x1_ASAP7_75t_R _26101_ (.A1(_03696_),
    .A2(_03705_),
    .B(_08844_),
    .Y(_03706_));
 NAND2x1_ASAP7_75t_R _26102_ (.A(_00476_),
    .B(net6454),
    .Y(_03707_));
 INVx1_ASAP7_75t_R _26103_ (.A(_03697_),
    .Y(_03708_));
 XOR2x2_ASAP7_75t_R _26104_ (.A(net6411),
    .B(_03700_),
    .Y(_03709_));
 NAND2x1_ASAP7_75t_R _26105_ (.A(_03708_),
    .B(_03709_),
    .Y(_03710_));
 NAND3x1_ASAP7_75t_R _26106_ (.A(_03710_),
    .B(_03703_),
    .C(net6656),
    .Y(_03711_));
 AOI21x1_ASAP7_75t_R _26107_ (.A1(_03707_),
    .A2(_03711_),
    .B(net6491),
    .Y(_03712_));
 NOR2x1_ASAP7_75t_R _26108_ (.A(_03706_),
    .B(_03712_),
    .Y(_03713_));
 OAI21x1_ASAP7_75t_R _26110_ (.A1(_03664_),
    .A2(_03672_),
    .B(_03678_),
    .Y(_03714_));
 OAI21x1_ASAP7_75t_R _26111_ (.A1(_03674_),
    .A2(_03677_),
    .B(net6478),
    .Y(_03715_));
 NAND2x2_ASAP7_75t_R _26112_ (.A(_03715_),
    .B(_03714_),
    .Y(_01275_));
 AOI21x1_ASAP7_75t_R _26113_ (.A1(_03703_),
    .A2(_03710_),
    .B(net6454),
    .Y(_03716_));
 OAI21x1_ASAP7_75t_R _26114_ (.A1(_03695_),
    .A2(_03716_),
    .B(_08844_),
    .Y(_03717_));
 INVx2_ASAP7_75t_R _26115_ (.A(_03717_),
    .Y(_03718_));
 AOI21x1_ASAP7_75t_R _26116_ (.A1(_03707_),
    .A2(_03711_),
    .B(_08844_),
    .Y(_03719_));
 NOR2x2_ASAP7_75t_R _26117_ (.A(_03718_),
    .B(_03719_),
    .Y(_03720_));
 INVx1_ASAP7_75t_R _26119_ (.A(_00690_),
    .Y(_03721_));
 XOR2x2_ASAP7_75t_R _26120_ (.A(_14978_),
    .B(_03721_),
    .Y(_03722_));
 XNOR2x2_ASAP7_75t_R _26121_ (.A(_00689_),
    .B(net6549),
    .Y(_03723_));
 XOR2x2_ASAP7_75t_R _26122_ (.A(_00594_),
    .B(_00626_),
    .Y(_03724_));
 XOR2x2_ASAP7_75t_R _26123_ (.A(_03723_),
    .B(_03724_),
    .Y(_03725_));
 NOR2x1_ASAP7_75t_R _26124_ (.A(_03722_),
    .B(_03725_),
    .Y(_03726_));
 AO21x1_ASAP7_75t_R _26125_ (.A1(_03725_),
    .A2(_03722_),
    .B(net6454),
    .Y(_03727_));
 AND2x2_ASAP7_75t_R _26126_ (.A(net6454),
    .B(_00528_),
    .Y(_03728_));
 INVx1_ASAP7_75t_R _26127_ (.A(_03728_),
    .Y(_03729_));
 OAI21x1_ASAP7_75t_R _26128_ (.A1(_03726_),
    .A2(_03727_),
    .B(_03729_),
    .Y(_03730_));
 XOR2x2_ASAP7_75t_R _26129_ (.A(_03730_),
    .B(net6490),
    .Y(_03731_));
 OAI21x1_ASAP7_75t_R _26130_ (.A1(net5676),
    .A2(net6139),
    .B(net4987),
    .Y(_03732_));
 NAND2x1p5_ASAP7_75t_R _26131_ (.A(_03732_),
    .B(net6136),
    .Y(_03733_));
 INVx2_ASAP7_75t_R _26132_ (.A(_03733_),
    .Y(_03734_));
 NAND3x1_ASAP7_75t_R _26133_ (.A(_03705_),
    .B(net6491),
    .C(_03696_),
    .Y(_03735_));
 INVx1_ASAP7_75t_R _26137_ (.A(net5041),
    .Y(_03739_));
 AO21x1_ASAP7_75t_R _26138_ (.A1(net5674),
    .A2(net6138),
    .B(_03739_),
    .Y(_03740_));
 INVx1_ASAP7_75t_R _26139_ (.A(_01284_),
    .Y(_03741_));
 AO21x1_ASAP7_75t_R _26140_ (.A1(net5674),
    .A2(net6138),
    .B(_03741_),
    .Y(_03742_));
 NAND2x1_ASAP7_75t_R _26141_ (.A(net5387),
    .B(net5389),
    .Y(_03743_));
 AOI21x1_ASAP7_75t_R _26144_ (.A1(_03742_),
    .A2(net5109),
    .B(net6135),
    .Y(_03746_));
 XNOR2x2_ASAP7_75t_R _26145_ (.A(_00690_),
    .B(net6549),
    .Y(_03747_));
 XOR2x2_ASAP7_75t_R _26146_ (.A(_03747_),
    .B(_12235_),
    .Y(_03748_));
 XNOR2x2_ASAP7_75t_R _26147_ (.A(_15010_),
    .B(_03748_),
    .Y(_03749_));
 NOR2x1_ASAP7_75t_R _26148_ (.A(net6655),
    .B(_00527_),
    .Y(_03750_));
 AO21x1_ASAP7_75t_R _26149_ (.A1(_03749_),
    .A2(net6654),
    .B(_03750_),
    .Y(_03751_));
 XOR2x2_ASAP7_75t_R _26150_ (.A(_03751_),
    .B(_00905_),
    .Y(_03752_));
 AOI211x1_ASAP7_75t_R _26153_ (.A1(net4462),
    .A2(net4649),
    .B(_03746_),
    .C(net6126),
    .Y(_03755_));
 XNOR2x2_ASAP7_75t_R _26154_ (.A(_00905_),
    .B(_03751_),
    .Y(_03756_));
 INVx1_ASAP7_75t_R _26157_ (.A(_01285_),
    .Y(_03759_));
 OAI21x1_ASAP7_75t_R _26158_ (.A1(net4871),
    .A2(net5388),
    .B(net6132),
    .Y(_03760_));
 NOR2x1_ASAP7_75t_R _26159_ (.A(net5046),
    .B(net5387),
    .Y(_03761_));
 NAND3x1_ASAP7_75t_R _26162_ (.A(_03691_),
    .B(net6479),
    .C(_03693_),
    .Y(_03764_));
 OAI21x1_ASAP7_75t_R _26163_ (.A1(net6398),
    .A2(_03686_),
    .B(_03692_),
    .Y(_03765_));
 AOI22x1_ASAP7_75t_R _26164_ (.A1(net5674),
    .A2(net6138),
    .B1(net6117),
    .B2(net5673),
    .Y(_03766_));
 OAI22x1_ASAP7_75t_R _26165_ (.A1(_03760_),
    .A2(_03761_),
    .B1(net6132),
    .B2(_03766_),
    .Y(_03767_));
 INVx1_ASAP7_75t_R _26166_ (.A(_12213_),
    .Y(_03768_));
 XOR2x2_ASAP7_75t_R _26167_ (.A(_12272_),
    .B(_12236_),
    .Y(_03769_));
 NOR2x1_ASAP7_75t_R _26168_ (.A(_03768_),
    .B(_03769_),
    .Y(_03770_));
 XOR2x2_ASAP7_75t_R _26169_ (.A(_12272_),
    .B(_00692_),
    .Y(_03771_));
 NOR2x1_ASAP7_75t_R _26170_ (.A(_12213_),
    .B(_03771_),
    .Y(_03772_));
 OAI21x1_ASAP7_75t_R _26171_ (.A1(_03770_),
    .A2(_03772_),
    .B(net6653),
    .Y(_03773_));
 INVx1_ASAP7_75t_R _26172_ (.A(_00906_),
    .Y(_03774_));
 NOR2x1_ASAP7_75t_R _26173_ (.A(net6655),
    .B(_00526_),
    .Y(_03775_));
 INVx1_ASAP7_75t_R _26174_ (.A(_03775_),
    .Y(_03776_));
 NAND3x1_ASAP7_75t_R _26175_ (.A(_03773_),
    .B(_03774_),
    .C(_03776_),
    .Y(_03777_));
 AO21x1_ASAP7_75t_R _26176_ (.A1(_03773_),
    .A2(_03776_),
    .B(_03774_),
    .Y(_03778_));
 NAND2x1_ASAP7_75t_R _26177_ (.A(_03777_),
    .B(_03778_),
    .Y(_03779_));
 OAI21x1_ASAP7_75t_R _26180_ (.A1(net6121),
    .A2(_03767_),
    .B(net5671),
    .Y(_03782_));
 XOR2x2_ASAP7_75t_R _26181_ (.A(_00692_),
    .B(_00693_),
    .Y(_03783_));
 XOR2x2_ASAP7_75t_R _26182_ (.A(_03783_),
    .B(_00660_),
    .Y(_03784_));
 XOR2x2_ASAP7_75t_R _26183_ (.A(_03784_),
    .B(_12318_),
    .Y(_03785_));
 NOR2x1_ASAP7_75t_R _26184_ (.A(net6655),
    .B(_00525_),
    .Y(_03786_));
 AO21x1_ASAP7_75t_R _26185_ (.A1(_03785_),
    .A2(net6657),
    .B(_03786_),
    .Y(_03787_));
 XOR2x2_ASAP7_75t_R _26186_ (.A(_03787_),
    .B(_00907_),
    .Y(_03788_));
 INVx1_ASAP7_75t_R _26187_ (.A(_03788_),
    .Y(_03789_));
 OAI21x1_ASAP7_75t_R _26189_ (.A1(_03755_),
    .A2(_03782_),
    .B(_03789_),
    .Y(_03791_));
 INVx1_ASAP7_75t_R _26191_ (.A(_01286_),
    .Y(_03793_));
 NAND2x1_ASAP7_75t_R _26193_ (.A(_03793_),
    .B(net5387),
    .Y(_03795_));
 NAND2x1p5_ASAP7_75t_R _26194_ (.A(_03765_),
    .B(_03764_),
    .Y(_03796_));
 INVx1_ASAP7_75t_R _26195_ (.A(net6490),
    .Y(_03797_));
 XOR2x2_ASAP7_75t_R _26196_ (.A(_03730_),
    .B(_03797_),
    .Y(_03798_));
 AOI21x1_ASAP7_75t_R _26198_ (.A1(net5388),
    .A2(net5384),
    .B(net6115),
    .Y(_03800_));
 NAND2x1_ASAP7_75t_R _26199_ (.A(net4648),
    .B(net5108),
    .Y(_03801_));
 INVx1_ASAP7_75t_R _26200_ (.A(_01279_),
    .Y(_03802_));
 OAI21x1_ASAP7_75t_R _26201_ (.A1(net5676),
    .A2(net6139),
    .B(_03802_),
    .Y(_03803_));
 INVx1_ASAP7_75t_R _26202_ (.A(_03803_),
    .Y(_03804_));
 NOR2x1_ASAP7_75t_R _26203_ (.A(net5677),
    .B(net5387),
    .Y(_03805_));
 OAI21x1_ASAP7_75t_R _26205_ (.A1(_03804_),
    .A2(_03805_),
    .B(net6115),
    .Y(_03807_));
 AO21x1_ASAP7_75t_R _26207_ (.A1(_03801_),
    .A2(_03807_),
    .B(net6121),
    .Y(_03809_));
 NAND2x1_ASAP7_75t_R _26208_ (.A(net5677),
    .B(net5387),
    .Y(_03810_));
 AO21x1_ASAP7_75t_R _26211_ (.A1(_03810_),
    .A2(_03742_),
    .B(net6135),
    .Y(_03813_));
 NAND2x1_ASAP7_75t_R _26212_ (.A(net5041),
    .B(net5386),
    .Y(_03814_));
 NAND2x1_ASAP7_75t_R _26213_ (.A(_03814_),
    .B(net5108),
    .Y(_03815_));
 AO21x1_ASAP7_75t_R _26214_ (.A1(_03813_),
    .A2(_03815_),
    .B(net6126),
    .Y(_03816_));
 AOI21x1_ASAP7_75t_R _26216_ (.A1(_03809_),
    .A2(_03816_),
    .B(net5670),
    .Y(_03818_));
 XOR2x2_ASAP7_75t_R _26217_ (.A(_15074_),
    .B(net6427),
    .Y(_03819_));
 XOR2x2_ASAP7_75t_R _26218_ (.A(_03819_),
    .B(net6433),
    .Y(_03820_));
 NOR2x1_ASAP7_75t_R _26219_ (.A(net6655),
    .B(_00524_),
    .Y(_03821_));
 AO21x1_ASAP7_75t_R _26220_ (.A1(_03820_),
    .A2(net6657),
    .B(_03821_),
    .Y(_03822_));
 XOR2x2_ASAP7_75t_R _26221_ (.A(_03822_),
    .B(_00908_),
    .Y(_03823_));
 OAI21x1_ASAP7_75t_R _26223_ (.A1(_03791_),
    .A2(_03818_),
    .B(net6108),
    .Y(_03825_));
 INVx2_ASAP7_75t_R _26224_ (.A(_03732_),
    .Y(_03826_));
 AO21x1_ASAP7_75t_R _26226_ (.A1(_03826_),
    .A2(net6112),
    .B(net6126),
    .Y(_03828_));
 INVx1_ASAP7_75t_R _26227_ (.A(_03828_),
    .Y(_03829_));
 OAI21x1_ASAP7_75t_R _26228_ (.A1(_03718_),
    .A2(net6137),
    .B(net4986),
    .Y(_03830_));
 INVx2_ASAP7_75t_R _26229_ (.A(_03830_),
    .Y(_03831_));
 NOR2x1_ASAP7_75t_R _26230_ (.A(net6111),
    .B(_03831_),
    .Y(_03832_));
 NAND2x1_ASAP7_75t_R _26231_ (.A(net5675),
    .B(net5388),
    .Y(_03833_));
 NOR2x1_ASAP7_75t_R _26232_ (.A(net6132),
    .B(_03833_),
    .Y(_03834_));
 NOR2x1_ASAP7_75t_R _26233_ (.A(_03832_),
    .B(_03834_),
    .Y(_03835_));
 AOI21x1_ASAP7_75t_R _26235_ (.A1(_03829_),
    .A2(_03835_),
    .B(net5671),
    .Y(_03837_));
 INVx1_ASAP7_75t_R _26236_ (.A(_01281_),
    .Y(_03838_));
 AO21x1_ASAP7_75t_R _26237_ (.A1(net5674),
    .A2(net6138),
    .B(_03838_),
    .Y(_03839_));
 OAI21x1_ASAP7_75t_R _26238_ (.A1(net5676),
    .A2(net6139),
    .B(_01277_),
    .Y(_03840_));
 AO21x1_ASAP7_75t_R _26239_ (.A1(_03839_),
    .A2(net4866),
    .B(net6134),
    .Y(_03841_));
 AO21x1_ASAP7_75t_R _26240_ (.A1(net5674),
    .A2(net6138),
    .B(_01277_),
    .Y(_03842_));
 NAND2x1_ASAP7_75t_R _26241_ (.A(_03842_),
    .B(net4462),
    .Y(_03843_));
 AO21x1_ASAP7_75t_R _26242_ (.A1(_03841_),
    .A2(_03843_),
    .B(net6122),
    .Y(_03844_));
 NAND2x1_ASAP7_75t_R _26243_ (.A(_03837_),
    .B(_03844_),
    .Y(_03845_));
 NAND2x1_ASAP7_75t_R _26244_ (.A(net5675),
    .B(net5384),
    .Y(_03846_));
 AOI21x1_ASAP7_75t_R _26246_ (.A1(_03846_),
    .A2(net5109),
    .B(net6112),
    .Y(_03848_));
 AOI21x1_ASAP7_75t_R _26247_ (.A1(net5387),
    .A2(net5390),
    .B(net6132),
    .Y(_03849_));
 AND2x2_ASAP7_75t_R _26248_ (.A(_03849_),
    .B(_03846_),
    .Y(_03850_));
 OAI21x1_ASAP7_75t_R _26249_ (.A1(_03848_),
    .A2(_03850_),
    .B(net6122),
    .Y(_03851_));
 AO21x1_ASAP7_75t_R _26250_ (.A1(net5674),
    .A2(net6138),
    .B(net4869),
    .Y(_03852_));
 INVx1_ASAP7_75t_R _26251_ (.A(net4987),
    .Y(_03853_));
 OA21x2_ASAP7_75t_R _26252_ (.A1(net6139),
    .A2(net5676),
    .B(_03853_),
    .Y(_03854_));
 INVx4_ASAP7_75t_R _26253_ (.A(_03854_),
    .Y(_03855_));
 AOI21x1_ASAP7_75t_R _26254_ (.A1(net4646),
    .A2(_03855_),
    .B(net6134),
    .Y(_03856_));
 OA21x2_ASAP7_75t_R _26255_ (.A1(net6139),
    .A2(net5676),
    .B(net5048),
    .Y(_03857_));
 INVx1_ASAP7_75t_R _26256_ (.A(_03857_),
    .Y(_03858_));
 INVx1_ASAP7_75t_R _26257_ (.A(_01277_),
    .Y(_03859_));
 NOR2x1_ASAP7_75t_R _26259_ (.A(_03859_),
    .B(net5387),
    .Y(_03861_));
 INVx1_ASAP7_75t_R _26260_ (.A(_03861_),
    .Y(_03862_));
 AOI21x1_ASAP7_75t_R _26262_ (.A1(_03858_),
    .A2(_03862_),
    .B(net6113),
    .Y(_03864_));
 OAI21x1_ASAP7_75t_R _26263_ (.A1(_03856_),
    .A2(_03864_),
    .B(net6126),
    .Y(_03865_));
 NAND3x1_ASAP7_75t_R _26264_ (.A(_03851_),
    .B(_03865_),
    .C(net5671),
    .Y(_03866_));
 AOI21x1_ASAP7_75t_R _26265_ (.A1(_03845_),
    .A2(_03866_),
    .B(net5669),
    .Y(_03867_));
 NAND2x1_ASAP7_75t_R _26267_ (.A(net5046),
    .B(net5386),
    .Y(_03869_));
 OAI21x1_ASAP7_75t_R _26268_ (.A1(net6133),
    .A2(_03869_),
    .B(net6120),
    .Y(_03870_));
 OA21x2_ASAP7_75t_R _26269_ (.A1(net6137),
    .A2(_03718_),
    .B(net5048),
    .Y(_03871_));
 NOR2x1_ASAP7_75t_R _26271_ (.A(net6110),
    .B(net4647),
    .Y(_03873_));
 AO21x1_ASAP7_75t_R _26272_ (.A1(net6110),
    .A2(_03871_),
    .B(_03873_),
    .Y(_03874_));
 OA21x2_ASAP7_75t_R _26273_ (.A1(_03731_),
    .A2(net4647),
    .B(net6123),
    .Y(_03875_));
 NAND2x1_ASAP7_75t_R _26274_ (.A(_03741_),
    .B(net5386),
    .Y(_03876_));
 AOI21x1_ASAP7_75t_R _26275_ (.A1(net5047),
    .A2(net5388),
    .B(net6110),
    .Y(_03877_));
 NAND2x1_ASAP7_75t_R _26276_ (.A(_03876_),
    .B(_03877_),
    .Y(_03878_));
 NAND2x1_ASAP7_75t_R _26277_ (.A(_03776_),
    .B(_03773_),
    .Y(_03879_));
 XOR2x2_ASAP7_75t_R _26278_ (.A(_03879_),
    .B(_00906_),
    .Y(_03880_));
 AOI21x1_ASAP7_75t_R _26280_ (.A1(_03875_),
    .A2(_03878_),
    .B(net5667),
    .Y(_03882_));
 OAI21x1_ASAP7_75t_R _26281_ (.A1(_03870_),
    .A2(_03874_),
    .B(_03882_),
    .Y(_03883_));
 OAI21x1_ASAP7_75t_R _26283_ (.A1(net5384),
    .A2(net5386),
    .B(_03840_),
    .Y(_03884_));
 OAI21x1_ASAP7_75t_R _26284_ (.A1(_03718_),
    .A2(net6137),
    .B(_03802_),
    .Y(_03885_));
 NOR2x1_ASAP7_75t_R _26285_ (.A(_03731_),
    .B(_03885_),
    .Y(_03886_));
 AOI21x1_ASAP7_75t_R _26286_ (.A1(net6136),
    .A2(_03884_),
    .B(_03886_),
    .Y(_03887_));
 OAI21x1_ASAP7_75t_R _26287_ (.A1(_03718_),
    .A2(net6137),
    .B(_03759_),
    .Y(_03888_));
 OAI21x1_ASAP7_75t_R _26288_ (.A1(net6133),
    .A2(net4644),
    .B(_03752_),
    .Y(_03889_));
 NOR2x1_ASAP7_75t_R _26289_ (.A(net6133),
    .B(_03869_),
    .Y(_03890_));
 NOR2x1_ASAP7_75t_R _26290_ (.A(_03889_),
    .B(_03890_),
    .Y(_03891_));
 NAND2x1_ASAP7_75t_R _26291_ (.A(_03887_),
    .B(_03891_),
    .Y(_03892_));
 AO21x1_ASAP7_75t_R _26293_ (.A1(_03735_),
    .A2(net6138),
    .B(net4987),
    .Y(_03894_));
 INVx1_ASAP7_75t_R _26295_ (.A(_01295_),
    .Y(_03896_));
 NOR2x1_ASAP7_75t_R _26296_ (.A(_03896_),
    .B(net6114),
    .Y(_03897_));
 AO21x1_ASAP7_75t_R _26297_ (.A1(net6114),
    .A2(net4733),
    .B(_03897_),
    .Y(_03898_));
 AOI21x1_ASAP7_75t_R _26298_ (.A1(net6122),
    .A2(_03898_),
    .B(net5670),
    .Y(_03899_));
 AOI21x1_ASAP7_75t_R _26299_ (.A1(_03892_),
    .A2(_03899_),
    .B(_03789_),
    .Y(_03900_));
 NAND2x1_ASAP7_75t_R _26300_ (.A(_03883_),
    .B(_03900_),
    .Y(_03901_));
 AOI21x1_ASAP7_75t_R _26301_ (.A1(_03795_),
    .A2(_03800_),
    .B(_03756_),
    .Y(_03902_));
 OAI21x1_ASAP7_75t_R _26302_ (.A1(net6135),
    .A2(net4643),
    .B(_03902_),
    .Y(_03903_));
 OA21x2_ASAP7_75t_R _26303_ (.A1(net6136),
    .A2(net4643),
    .B(net6122),
    .Y(_03904_));
 INVx1_ASAP7_75t_R _26304_ (.A(_01282_),
    .Y(_03905_));
 OAI21x1_ASAP7_75t_R _26305_ (.A1(net5676),
    .A2(net6139),
    .B(_03905_),
    .Y(_03906_));
 NOR2x1_ASAP7_75t_R _26306_ (.A(net6136),
    .B(net4642),
    .Y(_03907_));
 NOR2x1_ASAP7_75t_R _26307_ (.A(_03907_),
    .B(_03734_),
    .Y(_03908_));
 AOI21x1_ASAP7_75t_R _26308_ (.A1(_03904_),
    .A2(_03908_),
    .B(net5670),
    .Y(_03909_));
 NAND2x1_ASAP7_75t_R _26309_ (.A(_03903_),
    .B(_03909_),
    .Y(_03910_));
 NAND2x1_ASAP7_75t_R _26310_ (.A(net5043),
    .B(net5387),
    .Y(_03911_));
 AOI21x1_ASAP7_75t_R _26312_ (.A1(net6134),
    .A2(_03911_),
    .B(net6126),
    .Y(_03913_));
 OAI21x1_ASAP7_75t_R _26313_ (.A1(_03804_),
    .A2(_03861_),
    .B(net6112),
    .Y(_03914_));
 AOI21x1_ASAP7_75t_R _26314_ (.A1(_03913_),
    .A2(_03914_),
    .B(net5667),
    .Y(_03915_));
 AOI21x1_ASAP7_75t_R _26315_ (.A1(net5677),
    .A2(net5387),
    .B(net6136),
    .Y(_03916_));
 NAND2x1_ASAP7_75t_R _26316_ (.A(_03894_),
    .B(_03916_),
    .Y(_03917_));
 AO21x1_ASAP7_75t_R _26317_ (.A1(net5674),
    .A2(net6138),
    .B(net5048),
    .Y(_03918_));
 AOI21x1_ASAP7_75t_R _26318_ (.A1(net5387),
    .A2(net5384),
    .B(net6115),
    .Y(_03919_));
 AOI21x1_ASAP7_75t_R _26319_ (.A1(_03918_),
    .A2(_03919_),
    .B(net6120),
    .Y(_03920_));
 NAND2x1_ASAP7_75t_R _26320_ (.A(_03917_),
    .B(_03920_),
    .Y(_03921_));
 AOI21x1_ASAP7_75t_R _26321_ (.A1(_03915_),
    .A2(_03921_),
    .B(net6116),
    .Y(_03922_));
 AOI21x1_ASAP7_75t_R _26322_ (.A1(_03910_),
    .A2(_03922_),
    .B(net6108),
    .Y(_03923_));
 NAND2x1_ASAP7_75t_R _26323_ (.A(_03901_),
    .B(_03923_),
    .Y(_03924_));
 OAI21x1_ASAP7_75t_R _26324_ (.A1(_03825_),
    .A2(_03867_),
    .B(_03924_),
    .Y(_00112_));
 INVx1_ASAP7_75t_R _26325_ (.A(_03823_),
    .Y(_03925_));
 NOR2x1_ASAP7_75t_R _26326_ (.A(_03805_),
    .B(_03760_),
    .Y(_03926_));
 AO21x1_ASAP7_75t_R _26328_ (.A1(_03849_),
    .A2(_03842_),
    .B(net6122),
    .Y(_03928_));
 OAI21x1_ASAP7_75t_R _26329_ (.A1(_03926_),
    .A2(_03928_),
    .B(net5671),
    .Y(_03929_));
 NAND2x1_ASAP7_75t_R _26331_ (.A(net6109),
    .B(_03804_),
    .Y(_03931_));
 OAI21x1_ASAP7_75t_R _26332_ (.A1(net6109),
    .A2(net4866),
    .B(_03931_),
    .Y(_03932_));
 AOI22x1_ASAP7_75t_R _26333_ (.A1(net5674),
    .A2(net6138),
    .B1(net6140),
    .B2(_03687_),
    .Y(_03933_));
 AO21x1_ASAP7_75t_R _26334_ (.A1(_03933_),
    .A2(net6109),
    .B(net6123),
    .Y(_03934_));
 NOR2x1_ASAP7_75t_R _26335_ (.A(net6109),
    .B(net4732),
    .Y(_03935_));
 NOR3x1_ASAP7_75t_R _26336_ (.A(_03932_),
    .B(_03934_),
    .C(_03935_),
    .Y(_03936_));
 NOR2x1_ASAP7_75t_R _26337_ (.A(net4868),
    .B(net5386),
    .Y(_03937_));
 AO21x1_ASAP7_75t_R _26338_ (.A1(net5386),
    .A2(net5041),
    .B(net6136),
    .Y(_03938_));
 NOR2x1_ASAP7_75t_R _26339_ (.A(_03937_),
    .B(_03938_),
    .Y(_03939_));
 AOI21x1_ASAP7_75t_R _26340_ (.A1(net4870),
    .A2(net5388),
    .B(net6111),
    .Y(_03940_));
 AO21x1_ASAP7_75t_R _26342_ (.A1(_03940_),
    .A2(_03855_),
    .B(net6125),
    .Y(_03942_));
 AOI21x1_ASAP7_75t_R _26343_ (.A1(net6133),
    .A2(net4737),
    .B(net6120),
    .Y(_03943_));
 AOI21x1_ASAP7_75t_R _26345_ (.A1(net5388),
    .A2(net5384),
    .B(net6136),
    .Y(_03945_));
 NAND2x1_ASAP7_75t_R _26346_ (.A(net4648),
    .B(_03945_),
    .Y(_03946_));
 AOI21x1_ASAP7_75t_R _26347_ (.A1(_03943_),
    .A2(_03946_),
    .B(net5672),
    .Y(_03947_));
 OAI21x1_ASAP7_75t_R _26348_ (.A1(_03939_),
    .A2(_03942_),
    .B(_03947_),
    .Y(_03948_));
 OAI21x1_ASAP7_75t_R _26349_ (.A1(_03929_),
    .A2(_03936_),
    .B(_03948_),
    .Y(_03949_));
 INVx1_ASAP7_75t_R _26350_ (.A(net4648),
    .Y(_03950_));
 AO21x1_ASAP7_75t_R _26351_ (.A1(net5388),
    .A2(_03741_),
    .B(net6115),
    .Y(_03951_));
 NOR2x1_ASAP7_75t_R _26352_ (.A(_03950_),
    .B(_03951_),
    .Y(_03952_));
 INVx1_ASAP7_75t_R _26353_ (.A(_03842_),
    .Y(_03953_));
 AO21x1_ASAP7_75t_R _26354_ (.A1(net5384),
    .A2(net5387),
    .B(net6131),
    .Y(_03954_));
 NOR2x1_ASAP7_75t_R _26355_ (.A(net5668),
    .B(net6127),
    .Y(_03955_));
 OAI21x1_ASAP7_75t_R _26356_ (.A1(_03953_),
    .A2(_03954_),
    .B(_03955_),
    .Y(_03956_));
 NOR2x1_ASAP7_75t_R _26357_ (.A(_03952_),
    .B(_03956_),
    .Y(_03957_));
 NAND2x1_ASAP7_75t_R _26358_ (.A(net5677),
    .B(net5388),
    .Y(_03958_));
 AND2x2_ASAP7_75t_R _26359_ (.A(_03849_),
    .B(_03958_),
    .Y(_03959_));
 NOR2x1_ASAP7_75t_R _26360_ (.A(net5672),
    .B(net6127),
    .Y(_03960_));
 OAI21x1_ASAP7_75t_R _26361_ (.A1(net5107),
    .A2(_03760_),
    .B(_03960_),
    .Y(_03961_));
 NOR2x1_ASAP7_75t_R _26362_ (.A(_03959_),
    .B(_03961_),
    .Y(_03962_));
 NAND2x1_ASAP7_75t_R _26363_ (.A(net5042),
    .B(net5387),
    .Y(_03963_));
 AOI21x1_ASAP7_75t_R _26364_ (.A1(_03839_),
    .A2(_03963_),
    .B(net6131),
    .Y(_03964_));
 INVx1_ASAP7_75t_R _26365_ (.A(_01292_),
    .Y(_03965_));
 NAND2x1_ASAP7_75t_R _26367_ (.A(net6131),
    .B(net5668),
    .Y(_03967_));
 OAI21x1_ASAP7_75t_R _26368_ (.A1(_03965_),
    .A2(_03967_),
    .B(net6127),
    .Y(_03968_));
 OAI21x1_ASAP7_75t_R _26369_ (.A1(_03964_),
    .A2(_03968_),
    .B(net6116),
    .Y(_03969_));
 NOR3x1_ASAP7_75t_R _26370_ (.A(_03957_),
    .B(_03962_),
    .C(_03969_),
    .Y(_03970_));
 AOI21x1_ASAP7_75t_R _26371_ (.A1(net5669),
    .A2(_03949_),
    .B(_03970_),
    .Y(_03971_));
 NAND2x1_ASAP7_75t_R _26372_ (.A(net6490),
    .B(_03730_),
    .Y(_03972_));
 INVx1_ASAP7_75t_R _26373_ (.A(_03730_),
    .Y(_03973_));
 NAND2x1_ASAP7_75t_R _26374_ (.A(_03797_),
    .B(_03973_),
    .Y(_03974_));
 AOI21x1_ASAP7_75t_R _26375_ (.A1(_03972_),
    .A2(_03974_),
    .B(net5044),
    .Y(_03975_));
 AOI21x1_ASAP7_75t_R _26377_ (.A1(net5387),
    .A2(_03975_),
    .B(net6122),
    .Y(_03977_));
 NAND2x1_ASAP7_75t_R _26378_ (.A(_03855_),
    .B(_03940_),
    .Y(_03978_));
 AOI21x1_ASAP7_75t_R _26379_ (.A1(_03977_),
    .A2(_03978_),
    .B(net5667),
    .Y(_03979_));
 NAND2x1_ASAP7_75t_R _26380_ (.A(net5675),
    .B(net5386),
    .Y(_03980_));
 AOI21x1_ASAP7_75t_R _26382_ (.A1(net5040),
    .A2(net5388),
    .B(net6115),
    .Y(_03982_));
 AOI21x1_ASAP7_75t_R _26383_ (.A1(net5106),
    .A2(_03982_),
    .B(net6124),
    .Y(_03983_));
 OAI21x1_ASAP7_75t_R _26384_ (.A1(net6132),
    .A2(_03963_),
    .B(_03983_),
    .Y(_03984_));
 AOI21x1_ASAP7_75t_R _26385_ (.A1(_03979_),
    .A2(_03984_),
    .B(net6116),
    .Y(_03985_));
 AOI21x1_ASAP7_75t_R _26386_ (.A1(net5388),
    .A2(net5389),
    .B(net6132),
    .Y(_03986_));
 INVx1_ASAP7_75t_R _26387_ (.A(_03888_),
    .Y(_03987_));
 OAI21x1_ASAP7_75t_R _26388_ (.A1(net4502),
    .A2(net4555),
    .B(net6120),
    .Y(_03988_));
 AOI21x1_ASAP7_75t_R _26389_ (.A1(net4866),
    .A2(_03986_),
    .B(_03988_),
    .Y(_03989_));
 NAND2x1_ASAP7_75t_R _26390_ (.A(net5675),
    .B(net5390),
    .Y(_03990_));
 NAND2x1_ASAP7_75t_R _26391_ (.A(_03990_),
    .B(net5108),
    .Y(_03991_));
 AO21x1_ASAP7_75t_R _26392_ (.A1(net5109),
    .A2(net4736),
    .B(net6136),
    .Y(_03992_));
 AOI21x1_ASAP7_75t_R _26393_ (.A1(_03991_),
    .A2(_03992_),
    .B(net6120),
    .Y(_03993_));
 OAI21x1_ASAP7_75t_R _26395_ (.A1(_03989_),
    .A2(_03993_),
    .B(net5667),
    .Y(_03995_));
 NAND2x1_ASAP7_75t_R _26396_ (.A(_03985_),
    .B(_03995_),
    .Y(_03996_));
 NAND2x1_ASAP7_75t_R _26397_ (.A(_03911_),
    .B(_03986_),
    .Y(_03997_));
 AOI21x1_ASAP7_75t_R _26398_ (.A1(net4737),
    .A2(net5108),
    .B(net6125),
    .Y(_03998_));
 NAND2x1_ASAP7_75t_R _26399_ (.A(_03997_),
    .B(_03998_),
    .Y(_03999_));
 OA21x2_ASAP7_75t_R _26400_ (.A1(net6137),
    .A2(_03718_),
    .B(net5046),
    .Y(_04000_));
 AOI21x1_ASAP7_75t_R _26401_ (.A1(net6130),
    .A2(_04000_),
    .B(net6119),
    .Y(_04001_));
 NAND2x1_ASAP7_75t_R _26402_ (.A(_03846_),
    .B(_03916_),
    .Y(_04002_));
 AOI21x1_ASAP7_75t_R _26403_ (.A1(_04001_),
    .A2(_04002_),
    .B(net5667),
    .Y(_04003_));
 AOI21x1_ASAP7_75t_R _26404_ (.A1(_03999_),
    .A2(_04003_),
    .B(_03789_),
    .Y(_04004_));
 NOR2x1_ASAP7_75t_R _26405_ (.A(_03741_),
    .B(net5388),
    .Y(_04005_));
 OAI21x1_ASAP7_75t_R _26406_ (.A1(net4503),
    .A2(_04005_),
    .B(net6114),
    .Y(_04006_));
 NOR2x1_ASAP7_75t_R _26407_ (.A(net5041),
    .B(net5388),
    .Y(_04007_));
 NOR2x1_ASAP7_75t_R _26408_ (.A(net5387),
    .B(net4987),
    .Y(_04008_));
 OAI21x1_ASAP7_75t_R _26409_ (.A1(_04007_),
    .A2(_04008_),
    .B(net6136),
    .Y(_04009_));
 AOI21x1_ASAP7_75t_R _26410_ (.A1(_04006_),
    .A2(_04009_),
    .B(net6120),
    .Y(_04010_));
 INVx1_ASAP7_75t_R _26412_ (.A(net5105),
    .Y(_04012_));
 NAND2x1_ASAP7_75t_R _26413_ (.A(net6114),
    .B(_04012_),
    .Y(_04013_));
 INVx1_ASAP7_75t_R _26414_ (.A(_01296_),
    .Y(_04014_));
 NOR2x1_ASAP7_75t_R _26415_ (.A(_04014_),
    .B(net6114),
    .Y(_04015_));
 AOI21x1_ASAP7_75t_R _26416_ (.A1(net6113),
    .A2(net4503),
    .B(_04015_),
    .Y(_04016_));
 AOI21x1_ASAP7_75t_R _26418_ (.A1(_04013_),
    .A2(_04016_),
    .B(net6126),
    .Y(_04018_));
 OAI21x1_ASAP7_75t_R _26419_ (.A1(_04010_),
    .A2(_04018_),
    .B(net5667),
    .Y(_04019_));
 AOI21x1_ASAP7_75t_R _26420_ (.A1(_04004_),
    .A2(_04019_),
    .B(net6108),
    .Y(_04020_));
 NAND2x1_ASAP7_75t_R _26421_ (.A(_03996_),
    .B(_04020_),
    .Y(_04021_));
 OAI21x1_ASAP7_75t_R _26422_ (.A1(_03925_),
    .A2(_03971_),
    .B(_04021_),
    .Y(_00113_));
 NOR2x1_ASAP7_75t_R _26423_ (.A(_03965_),
    .B(net6134),
    .Y(_04022_));
 AOI21x1_ASAP7_75t_R _26424_ (.A1(_03958_),
    .A2(_03990_),
    .B(net6112),
    .Y(_04023_));
 OAI21x1_ASAP7_75t_R _26425_ (.A1(_04022_),
    .A2(_04023_),
    .B(net6127),
    .Y(_04024_));
 AOI21x1_ASAP7_75t_R _26426_ (.A1(net4734),
    .A2(_03858_),
    .B(net6113),
    .Y(_04025_));
 AOI21x1_ASAP7_75t_R _26427_ (.A1(_03810_),
    .A2(_03862_),
    .B(net6135),
    .Y(_04026_));
 OAI21x1_ASAP7_75t_R _26428_ (.A1(_04025_),
    .A2(_04026_),
    .B(net6121),
    .Y(_04027_));
 AOI21x1_ASAP7_75t_R _26429_ (.A1(_04024_),
    .A2(_04027_),
    .B(net5670),
    .Y(_04028_));
 AOI21x1_ASAP7_75t_R _26430_ (.A1(net4733),
    .A2(_03869_),
    .B(net6114),
    .Y(_04029_));
 AO21x1_ASAP7_75t_R _26431_ (.A1(_03896_),
    .A2(net6114),
    .B(net6122),
    .Y(_04030_));
 OAI21x1_ASAP7_75t_R _26432_ (.A1(_04029_),
    .A2(_04030_),
    .B(net5670),
    .Y(_04031_));
 AND2x2_ASAP7_75t_R _26433_ (.A(_03919_),
    .B(_03833_),
    .Y(_04032_));
 AO21x1_ASAP7_75t_R _26434_ (.A1(_03916_),
    .A2(net4733),
    .B(net6126),
    .Y(_04033_));
 NOR2x1_ASAP7_75t_R _26435_ (.A(_04032_),
    .B(_04033_),
    .Y(_04034_));
 OAI21x1_ASAP7_75t_R _26436_ (.A1(_04031_),
    .A2(_04034_),
    .B(_03789_),
    .Y(_04035_));
 OAI21x1_ASAP7_75t_R _26437_ (.A1(_04028_),
    .A2(_04035_),
    .B(_03925_),
    .Y(_04036_));
 AO21x1_ASAP7_75t_R _26438_ (.A1(net5388),
    .A2(_03741_),
    .B(net6136),
    .Y(_04037_));
 NAND2x1_ASAP7_75t_R _26439_ (.A(_01294_),
    .B(net6134),
    .Y(_04038_));
 AO21x1_ASAP7_75t_R _26440_ (.A1(_04037_),
    .A2(_04038_),
    .B(net6121),
    .Y(_04039_));
 NOR2x1_ASAP7_75t_R _26441_ (.A(_01297_),
    .B(net6134),
    .Y(_04040_));
 INVx1_ASAP7_75t_R _26442_ (.A(_03810_),
    .Y(_04041_));
 NOR2x1_ASAP7_75t_R _26443_ (.A(_04041_),
    .B(_03951_),
    .Y(_04042_));
 OAI21x1_ASAP7_75t_R _26444_ (.A1(_04040_),
    .A2(_04042_),
    .B(net6121),
    .Y(_04043_));
 AOI21x1_ASAP7_75t_R _26445_ (.A1(_04039_),
    .A2(_04043_),
    .B(net5670),
    .Y(_04044_));
 INVx1_ASAP7_75t_R _26446_ (.A(_03840_),
    .Y(_04045_));
 AO21x1_ASAP7_75t_R _26447_ (.A1(_04045_),
    .A2(net6115),
    .B(net6122),
    .Y(_04046_));
 OA21x2_ASAP7_75t_R _26448_ (.A1(net4553),
    .A2(_03987_),
    .B(net6130),
    .Y(_04047_));
 OAI21x1_ASAP7_75t_R _26449_ (.A1(_04046_),
    .A2(_04047_),
    .B(net5670),
    .Y(_04048_));
 AND2x2_ASAP7_75t_R _26450_ (.A(_01279_),
    .B(net5045),
    .Y(_04049_));
 AOI21x1_ASAP7_75t_R _26451_ (.A1(net5387),
    .A2(_04049_),
    .B(_03798_),
    .Y(_04050_));
 AO21x1_ASAP7_75t_R _26452_ (.A1(net5674),
    .A2(net6138),
    .B(net5042),
    .Y(_04051_));
 AOI211x1_ASAP7_75t_R _26453_ (.A1(_04050_),
    .A2(_04051_),
    .B(_03964_),
    .C(net6124),
    .Y(_04052_));
 OAI21x1_ASAP7_75t_R _26454_ (.A1(_04048_),
    .A2(_04052_),
    .B(net6116),
    .Y(_04053_));
 NOR2x1_ASAP7_75t_R _26455_ (.A(_04044_),
    .B(_04053_),
    .Y(_04054_));
 NOR2x1_ASAP7_75t_R _26456_ (.A(_04008_),
    .B(net4555),
    .Y(_04055_));
 OA21x2_ASAP7_75t_R _26457_ (.A1(net6137),
    .A2(_03718_),
    .B(_03905_),
    .Y(_04056_));
 INVx1_ASAP7_75t_R _26458_ (.A(_04056_),
    .Y(_04057_));
 AOI21x1_ASAP7_75t_R _26459_ (.A1(net5109),
    .A2(_04057_),
    .B(net6129),
    .Y(_04058_));
 OAI21x1_ASAP7_75t_R _26460_ (.A1(_04058_),
    .A2(_04055_),
    .B(net6123),
    .Y(_04059_));
 INVx1_ASAP7_75t_R _26461_ (.A(_03906_),
    .Y(_04060_));
 AO21x1_ASAP7_75t_R _26462_ (.A1(net5388),
    .A2(net5675),
    .B(net6109),
    .Y(_04061_));
 AO21x1_ASAP7_75t_R _26463_ (.A1(net5674),
    .A2(net6138),
    .B(net5040),
    .Y(_04062_));
 AOI21x1_ASAP7_75t_R _26464_ (.A1(_04062_),
    .A2(_03849_),
    .B(net6124),
    .Y(_04063_));
 OAI21x1_ASAP7_75t_R _26465_ (.A1(_04060_),
    .A2(_04061_),
    .B(_04063_),
    .Y(_04064_));
 AOI21x1_ASAP7_75t_R _26467_ (.A1(_04064_),
    .A2(_04059_),
    .B(net6116),
    .Y(_04066_));
 INVx1_ASAP7_75t_R _26468_ (.A(_04007_),
    .Y(_04067_));
 AOI21x1_ASAP7_75t_R _26469_ (.A1(net4646),
    .A2(_04067_),
    .B(net6113),
    .Y(_04068_));
 NAND2x1_ASAP7_75t_R _26470_ (.A(net6126),
    .B(_04037_),
    .Y(_04069_));
 OAI21x1_ASAP7_75t_R _26471_ (.A1(_04068_),
    .A2(_04069_),
    .B(net6116),
    .Y(_04070_));
 AOI21x1_ASAP7_75t_R _26472_ (.A1(net5675),
    .A2(net5388),
    .B(_03731_),
    .Y(_04071_));
 NAND2x1_ASAP7_75t_R _26473_ (.A(_03855_),
    .B(_04071_),
    .Y(_04072_));
 NAND3x1_ASAP7_75t_R _26474_ (.A(net5109),
    .B(net6129),
    .C(net4645),
    .Y(_04073_));
 AOI21x1_ASAP7_75t_R _26475_ (.A1(_04072_),
    .A2(_04073_),
    .B(net6123),
    .Y(_04074_));
 OAI21x1_ASAP7_75t_R _26476_ (.A1(_04070_),
    .A2(_04074_),
    .B(net5670),
    .Y(_04075_));
 OAI21x1_ASAP7_75t_R _26477_ (.A1(_04075_),
    .A2(_04066_),
    .B(net6108),
    .Y(_04076_));
 INVx1_ASAP7_75t_R _26478_ (.A(_03740_),
    .Y(_04077_));
 AO21x1_ASAP7_75t_R _26479_ (.A1(net5387),
    .A2(net5043),
    .B(net6132),
    .Y(_04078_));
 NOR2x1_ASAP7_75t_R _26480_ (.A(_04077_),
    .B(_04078_),
    .Y(_04079_));
 OAI21x1_ASAP7_75t_R _26481_ (.A1(_04042_),
    .A2(_04079_),
    .B(net6121),
    .Y(_04080_));
 NAND2x1_ASAP7_75t_R _26482_ (.A(net6136),
    .B(net4643),
    .Y(_04081_));
 OAI21x1_ASAP7_75t_R _26483_ (.A1(_04005_),
    .A2(_04081_),
    .B(net6126),
    .Y(_04082_));
 INVx1_ASAP7_75t_R _26484_ (.A(_04082_),
    .Y(_04083_));
 AOI21x1_ASAP7_75t_R _26485_ (.A1(_03917_),
    .A2(_04083_),
    .B(_03789_),
    .Y(_04084_));
 NAND2x1_ASAP7_75t_R _26486_ (.A(_04080_),
    .B(_04084_),
    .Y(_04085_));
 OA211x2_ASAP7_75t_R _26487_ (.A1(_03810_),
    .A2(net6113),
    .B(net6126),
    .C(net4643),
    .Y(_04086_));
 AO21x1_ASAP7_75t_R _26488_ (.A1(net5388),
    .A2(net4872),
    .B(net6133),
    .Y(_04087_));
 INVx1_ASAP7_75t_R _26489_ (.A(_04081_),
    .Y(_04088_));
 NAND2x1_ASAP7_75t_R _26490_ (.A(net5109),
    .B(_04088_),
    .Y(_04089_));
 AOI21x1_ASAP7_75t_R _26491_ (.A1(_04087_),
    .A2(_04089_),
    .B(net6126),
    .Y(_04090_));
 NOR2x1_ASAP7_75t_R _26492_ (.A(net6116),
    .B(net4504),
    .Y(_04091_));
 OAI21x1_ASAP7_75t_R _26493_ (.A1(_04086_),
    .A2(_04090_),
    .B(_04091_),
    .Y(_04092_));
 AOI21x1_ASAP7_75t_R _26494_ (.A1(_04085_),
    .A2(_04092_),
    .B(net5670),
    .Y(_04093_));
 OAI22x1_ASAP7_75t_R _26495_ (.A1(_04036_),
    .A2(_04054_),
    .B1(_04076_),
    .B2(_04093_),
    .Y(_00114_));
 NAND2x1_ASAP7_75t_R _26496_ (.A(_03740_),
    .B(_04050_),
    .Y(_04094_));
 AOI21x1_ASAP7_75t_R _26497_ (.A1(net4737),
    .A2(_03945_),
    .B(net5672),
    .Y(_04095_));
 NAND2x1_ASAP7_75t_R _26498_ (.A(_04094_),
    .B(_04095_),
    .Y(_04096_));
 OA21x2_ASAP7_75t_R _26499_ (.A1(net4642),
    .A2(net6110),
    .B(net5672),
    .Y(_04097_));
 NAND2x1_ASAP7_75t_R _26500_ (.A(net5386),
    .B(net5384),
    .Y(_04098_));
 AOI21x1_ASAP7_75t_R _26501_ (.A1(net5047),
    .A2(net5388),
    .B(_03731_),
    .Y(_04099_));
 NAND2x1_ASAP7_75t_R _26502_ (.A(_04098_),
    .B(_04099_),
    .Y(_04100_));
 AOI21x1_ASAP7_75t_R _26503_ (.A1(_04097_),
    .A2(_04100_),
    .B(net6118),
    .Y(_04101_));
 NAND2x1_ASAP7_75t_R _26504_ (.A(_04096_),
    .B(_04101_),
    .Y(_04102_));
 AND3x1_ASAP7_75t_R _26505_ (.A(net6110),
    .B(net5672),
    .C(_03826_),
    .Y(_04103_));
 AOI21x1_ASAP7_75t_R _26506_ (.A1(net4867),
    .A2(net5388),
    .B(net5672),
    .Y(_04104_));
 NAND2x1_ASAP7_75t_R _26507_ (.A(_03916_),
    .B(_04104_),
    .Y(_04105_));
 NOR2x1_ASAP7_75t_R _26508_ (.A(net6110),
    .B(net5672),
    .Y(_04106_));
 AOI21x1_ASAP7_75t_R _26509_ (.A1(_03831_),
    .A2(_04106_),
    .B(_03873_),
    .Y(_04107_));
 NAND2x1_ASAP7_75t_R _26510_ (.A(_04105_),
    .B(_04107_),
    .Y(_04108_));
 OAI21x1_ASAP7_75t_R _26511_ (.A1(_04103_),
    .A2(_04108_),
    .B(net6118),
    .Y(_04109_));
 AOI21x1_ASAP7_75t_R _26512_ (.A1(_04109_),
    .A2(_04102_),
    .B(_03789_),
    .Y(_04110_));
 OA21x2_ASAP7_75t_R _26513_ (.A1(net6139),
    .A2(net5676),
    .B(net5042),
    .Y(_04111_));
 OAI21x1_ASAP7_75t_R _26514_ (.A1(_03871_),
    .A2(_04111_),
    .B(net6109),
    .Y(_04112_));
 NOR2x1_ASAP7_75t_R _26515_ (.A(_04049_),
    .B(net5388),
    .Y(_04113_));
 OAI21x1_ASAP7_75t_R _26516_ (.A1(_04056_),
    .A2(_04113_),
    .B(net6129),
    .Y(_04114_));
 AOI21x1_ASAP7_75t_R _26517_ (.A1(_04112_),
    .A2(_04114_),
    .B(net6118),
    .Y(_04115_));
 OAI21x1_ASAP7_75t_R _26518_ (.A1(_04063_),
    .A2(_04115_),
    .B(net5667),
    .Y(_04116_));
 OA21x2_ASAP7_75t_R _26519_ (.A1(net6137),
    .A2(_03718_),
    .B(net4872),
    .Y(_04117_));
 OAI21x1_ASAP7_75t_R _26520_ (.A1(net4553),
    .A2(_04117_),
    .B(net6109),
    .Y(_04118_));
 OAI21x1_ASAP7_75t_R _26521_ (.A1(_04060_),
    .A2(_03766_),
    .B(net6132),
    .Y(_04119_));
 AOI21x1_ASAP7_75t_R _26522_ (.A1(_04118_),
    .A2(_04119_),
    .B(net6124),
    .Y(_04120_));
 OAI21x1_ASAP7_75t_R _26523_ (.A1(_04045_),
    .A2(_03933_),
    .B(net6132),
    .Y(_04121_));
 AOI21x1_ASAP7_75t_R _26524_ (.A1(_04121_),
    .A2(_04002_),
    .B(net6119),
    .Y(_04122_));
 OAI21x1_ASAP7_75t_R _26525_ (.A1(_04120_),
    .A2(_04122_),
    .B(net5672),
    .Y(_04123_));
 AOI21x1_ASAP7_75t_R _26526_ (.A1(_04116_),
    .A2(_04123_),
    .B(net6116),
    .Y(_04124_));
 OAI21x1_ASAP7_75t_R _26527_ (.A1(_04110_),
    .A2(_04124_),
    .B(net6108),
    .Y(_04125_));
 NOR2x1_ASAP7_75t_R _26528_ (.A(net5677),
    .B(net5390),
    .Y(_04126_));
 OAI21x1_ASAP7_75t_R _26529_ (.A1(_03933_),
    .A2(_04126_),
    .B(net6109),
    .Y(_04127_));
 OAI21x1_ASAP7_75t_R _26530_ (.A1(_03826_),
    .A2(_04061_),
    .B(_04127_),
    .Y(_04128_));
 AOI21x1_ASAP7_75t_R _26531_ (.A1(net6128),
    .A2(net4736),
    .B(net6123),
    .Y(_04129_));
 NAND2x1_ASAP7_75t_R _26532_ (.A(_04098_),
    .B(_04071_),
    .Y(_04130_));
 AOI21x1_ASAP7_75t_R _26533_ (.A1(_04129_),
    .A2(_04130_),
    .B(net5672),
    .Y(_04131_));
 OAI21x1_ASAP7_75t_R _26534_ (.A1(net6118),
    .A2(_04128_),
    .B(_04131_),
    .Y(_04132_));
 OAI21x1_ASAP7_75t_R _26535_ (.A1(net5386),
    .A2(net5384),
    .B(net6110),
    .Y(_04133_));
 NOR2x1_ASAP7_75t_R _26536_ (.A(_03857_),
    .B(_04133_),
    .Y(_04134_));
 AND3x1_ASAP7_75t_R _26537_ (.A(net4736),
    .B(_03840_),
    .C(net6136),
    .Y(_04135_));
 OAI21x1_ASAP7_75t_R _26538_ (.A1(_04134_),
    .A2(_04135_),
    .B(net6118),
    .Y(_04136_));
 OAI21x1_ASAP7_75t_R _26539_ (.A1(net4502),
    .A2(_04007_),
    .B(net6136),
    .Y(_04137_));
 AOI21x1_ASAP7_75t_R _26540_ (.A1(_03855_),
    .A2(_04071_),
    .B(net6118),
    .Y(_04138_));
 AOI21x1_ASAP7_75t_R _26541_ (.A1(_04137_),
    .A2(_04138_),
    .B(net5667),
    .Y(_04139_));
 NAND2x1_ASAP7_75t_R _26542_ (.A(_04136_),
    .B(_04139_),
    .Y(_04140_));
 AOI21x1_ASAP7_75t_R _26543_ (.A1(_04132_),
    .A2(_04140_),
    .B(_03789_),
    .Y(_04141_));
 OAI21x1_ASAP7_75t_R _26544_ (.A1(_03857_),
    .A2(_04000_),
    .B(net6128),
    .Y(_04142_));
 OAI21x1_ASAP7_75t_R _26545_ (.A1(_04111_),
    .A2(_04008_),
    .B(net6109),
    .Y(_04143_));
 AOI21x1_ASAP7_75t_R _26546_ (.A1(_04142_),
    .A2(_04143_),
    .B(net6118),
    .Y(_04144_));
 OAI21x1_ASAP7_75t_R _26547_ (.A1(net4554),
    .A2(_03871_),
    .B(net6109),
    .Y(_04145_));
 NOR2x1_ASAP7_75t_R _26548_ (.A(net5675),
    .B(net5390),
    .Y(_04146_));
 OAI21x1_ASAP7_75t_R _26549_ (.A1(_03933_),
    .A2(_04146_),
    .B(net6128),
    .Y(_04147_));
 AOI21x1_ASAP7_75t_R _26550_ (.A1(_04145_),
    .A2(_04147_),
    .B(net6123),
    .Y(_04148_));
 OAI21x1_ASAP7_75t_R _26551_ (.A1(_04144_),
    .A2(_04148_),
    .B(net5672),
    .Y(_04149_));
 OAI21x1_ASAP7_75t_R _26552_ (.A1(_03826_),
    .A2(_04056_),
    .B(net6109),
    .Y(_04150_));
 NAND2x1_ASAP7_75t_R _26553_ (.A(net5106),
    .B(_03982_),
    .Y(_04151_));
 AOI21x1_ASAP7_75t_R _26554_ (.A1(_04150_),
    .A2(_04151_),
    .B(net6123),
    .Y(_04152_));
 AOI21x1_ASAP7_75t_R _26555_ (.A1(_03951_),
    .A2(_04127_),
    .B(net6118),
    .Y(_04153_));
 OAI21x1_ASAP7_75t_R _26556_ (.A1(_04152_),
    .A2(_04153_),
    .B(net5667),
    .Y(_04154_));
 AOI21x1_ASAP7_75t_R _26557_ (.A1(_04149_),
    .A2(_04154_),
    .B(net6116),
    .Y(_04155_));
 OAI21x1_ASAP7_75t_R _26558_ (.A1(_04141_),
    .A2(_04155_),
    .B(_03925_),
    .Y(_04156_));
 NAND2x1_ASAP7_75t_R _26559_ (.A(_04156_),
    .B(_04125_),
    .Y(_00115_));
 AOI21x1_ASAP7_75t_R _26560_ (.A1(_03741_),
    .A2(net5387),
    .B(net6115),
    .Y(_04157_));
 INVx1_ASAP7_75t_R _26561_ (.A(_04157_),
    .Y(_04158_));
 NOR2x1_ASAP7_75t_R _26562_ (.A(_03805_),
    .B(_04158_),
    .Y(_04159_));
 OAI21x1_ASAP7_75t_R _26563_ (.A1(_04077_),
    .A2(_04078_),
    .B(net6122),
    .Y(_04160_));
 NOR2x1_ASAP7_75t_R _26564_ (.A(_04159_),
    .B(_04160_),
    .Y(_04161_));
 AOI21x1_ASAP7_75t_R _26565_ (.A1(net4866),
    .A2(_03958_),
    .B(net6112),
    .Y(_04162_));
 NAND2x1_ASAP7_75t_R _26566_ (.A(net6114),
    .B(_04005_),
    .Y(_04163_));
 AOI21x1_ASAP7_75t_R _26567_ (.A1(net5388),
    .A2(_03975_),
    .B(net6119),
    .Y(_04164_));
 NAND2x1_ASAP7_75t_R _26568_ (.A(_04163_),
    .B(_04164_),
    .Y(_04165_));
 OAI21x1_ASAP7_75t_R _26569_ (.A1(_04162_),
    .A2(_04165_),
    .B(net5667),
    .Y(_04166_));
 NOR2x1_ASAP7_75t_R _26570_ (.A(_04161_),
    .B(_04166_),
    .Y(_04167_));
 AO21x1_ASAP7_75t_R _26571_ (.A1(_03987_),
    .A2(net6115),
    .B(net6126),
    .Y(_04168_));
 AO21x1_ASAP7_75t_R _26572_ (.A1(_04008_),
    .A2(net6132),
    .B(_04060_),
    .Y(_04169_));
 OAI21x1_ASAP7_75t_R _26573_ (.A1(_04168_),
    .A2(_04169_),
    .B(net5670),
    .Y(_04170_));
 NOR2x1_ASAP7_75t_R _26574_ (.A(_03831_),
    .B(_03938_),
    .Y(_04171_));
 AO21x1_ASAP7_75t_R _26575_ (.A1(_03877_),
    .A2(_03876_),
    .B(net6118),
    .Y(_04172_));
 NOR2x1_ASAP7_75t_R _26576_ (.A(_04171_),
    .B(_04172_),
    .Y(_04173_));
 OAI21x1_ASAP7_75t_R _26577_ (.A1(_04170_),
    .A2(_04173_),
    .B(net6116),
    .Y(_04174_));
 OAI21x1_ASAP7_75t_R _26578_ (.A1(_04167_),
    .A2(_04174_),
    .B(_03925_),
    .Y(_04175_));
 AO21x1_ASAP7_75t_R _26579_ (.A1(net5106),
    .A2(_03842_),
    .B(net6109),
    .Y(_04176_));
 NAND2x1_ASAP7_75t_R _26580_ (.A(net5677),
    .B(net5390),
    .Y(_04177_));
 AO21x1_ASAP7_75t_R _26581_ (.A1(_04177_),
    .A2(net5106),
    .B(net6131),
    .Y(_04178_));
 AOI21x1_ASAP7_75t_R _26582_ (.A1(_04176_),
    .A2(_04178_),
    .B(net6127),
    .Y(_04179_));
 AO21x1_ASAP7_75t_R _26583_ (.A1(net5387),
    .A2(net5677),
    .B(net6109),
    .Y(_04180_));
 OAI21x1_ASAP7_75t_R _26584_ (.A1(_04126_),
    .A2(_04180_),
    .B(net6127),
    .Y(_04181_));
 OAI21x1_ASAP7_75t_R _26585_ (.A1(_03959_),
    .A2(_04181_),
    .B(net5668),
    .Y(_04182_));
 NOR2x1_ASAP7_75t_R _26586_ (.A(_04179_),
    .B(_04182_),
    .Y(_04183_));
 AND2x2_ASAP7_75t_R _26587_ (.A(_03919_),
    .B(_03958_),
    .Y(_04184_));
 OAI21x1_ASAP7_75t_R _26588_ (.A1(_03953_),
    .A2(_03954_),
    .B(net6127),
    .Y(_04185_));
 NOR2x1_ASAP7_75t_R _26589_ (.A(_04184_),
    .B(_04185_),
    .Y(_04186_));
 NOR2x1_ASAP7_75t_R _26590_ (.A(net4505),
    .B(net4865),
    .Y(_04187_));
 AO21x1_ASAP7_75t_R _26591_ (.A1(_04187_),
    .A2(net6122),
    .B(net5668),
    .Y(_04188_));
 OAI21x1_ASAP7_75t_R _26592_ (.A1(_04186_),
    .A2(_04188_),
    .B(net5669),
    .Y(_04189_));
 NOR2x1_ASAP7_75t_R _26593_ (.A(_04183_),
    .B(_04189_),
    .Y(_04190_));
 AO21x1_ASAP7_75t_R _26594_ (.A1(net4735),
    .A2(net5388),
    .B(_04078_),
    .Y(_04191_));
 OAI21x1_ASAP7_75t_R _26595_ (.A1(net6136),
    .A2(_03937_),
    .B(net6118),
    .Y(_04192_));
 OAI21x1_ASAP7_75t_R _26596_ (.A1(_03940_),
    .A2(_04192_),
    .B(net5672),
    .Y(_04193_));
 AOI21x1_ASAP7_75t_R _26597_ (.A1(_03902_),
    .A2(_04191_),
    .B(_04193_),
    .Y(_04194_));
 NAND2x1_ASAP7_75t_R _26598_ (.A(net6109),
    .B(_04045_),
    .Y(_04195_));
 OAI21x1_ASAP7_75t_R _26599_ (.A1(net5107),
    .A2(_03760_),
    .B(_04195_),
    .Y(_04196_));
 AO21x1_ASAP7_75t_R _26600_ (.A1(net5107),
    .A2(net6109),
    .B(net6127),
    .Y(_04197_));
 NOR2x1_ASAP7_75t_R _26601_ (.A(_04196_),
    .B(_04197_),
    .Y(_04198_));
 NAND2x1_ASAP7_75t_R _26602_ (.A(net4649),
    .B(_03849_),
    .Y(_04199_));
 OA21x2_ASAP7_75t_R _26603_ (.A1(net5387),
    .A2(net6109),
    .B(net6127),
    .Y(_04200_));
 AO21x1_ASAP7_75t_R _26604_ (.A1(_04199_),
    .A2(_04200_),
    .B(net5671),
    .Y(_04201_));
 OAI21x1_ASAP7_75t_R _26605_ (.A1(_04198_),
    .A2(_04201_),
    .B(net5669),
    .Y(_04202_));
 OAI21x1_ASAP7_75t_R _26606_ (.A1(_04194_),
    .A2(_04202_),
    .B(net6108),
    .Y(_04203_));
 NOR2x1_ASAP7_75t_R _26607_ (.A(net6122),
    .B(_03848_),
    .Y(_04204_));
 NAND2x1_ASAP7_75t_R _26608_ (.A(net4441),
    .B(_04204_),
    .Y(_04205_));
 NAND2x1_ASAP7_75t_R _26609_ (.A(net5109),
    .B(net4865),
    .Y(_04206_));
 NAND2x1_ASAP7_75t_R _26610_ (.A(net5677),
    .B(net5384),
    .Y(_04207_));
 NAND2x1_ASAP7_75t_R _26611_ (.A(_03833_),
    .B(_04207_),
    .Y(_04208_));
 OA21x2_ASAP7_75t_R _26612_ (.A1(_04208_),
    .A2(net6134),
    .B(net6122),
    .Y(_04209_));
 AOI21x1_ASAP7_75t_R _26613_ (.A1(_04206_),
    .A2(_04209_),
    .B(net5671),
    .Y(_04210_));
 AOI21x1_ASAP7_75t_R _26614_ (.A1(net5106),
    .A2(net4865),
    .B(_03870_),
    .Y(_04211_));
 NOR2x1_ASAP7_75t_R _26615_ (.A(net6109),
    .B(_04008_),
    .Y(_04212_));
 AO21x1_ASAP7_75t_R _26616_ (.A1(net5042),
    .A2(net6109),
    .B(net6119),
    .Y(_04213_));
 OAI21x1_ASAP7_75t_R _26617_ (.A1(_04212_),
    .A2(_04213_),
    .B(net5672),
    .Y(_04214_));
 OAI21x1_ASAP7_75t_R _26618_ (.A1(_04211_),
    .A2(_04214_),
    .B(net6116),
    .Y(_04215_));
 AOI21x1_ASAP7_75t_R _26619_ (.A1(_04205_),
    .A2(_04210_),
    .B(_04215_),
    .Y(_04216_));
 OAI22x1_ASAP7_75t_R _26620_ (.A1(_04175_),
    .A2(_04190_),
    .B1(_04203_),
    .B2(_04216_),
    .Y(_00116_));
 AND3x1_ASAP7_75t_R _26621_ (.A(_03855_),
    .B(_03740_),
    .C(net6114),
    .Y(_04217_));
 AO21x1_ASAP7_75t_R _26622_ (.A1(_03734_),
    .A2(_03918_),
    .B(net6126),
    .Y(_04218_));
 AO21x1_ASAP7_75t_R _26623_ (.A1(net5386),
    .A2(net4870),
    .B(net6133),
    .Y(_04219_));
 OA21x2_ASAP7_75t_R _26624_ (.A1(net4867),
    .A2(net6111),
    .B(net6125),
    .Y(_04220_));
 AOI21x1_ASAP7_75t_R _26625_ (.A1(_04219_),
    .A2(_04220_),
    .B(net5672),
    .Y(_04221_));
 OA21x2_ASAP7_75t_R _26626_ (.A1(_04217_),
    .A2(_04218_),
    .B(_04221_),
    .Y(_04222_));
 OA21x2_ASAP7_75t_R _26627_ (.A1(_04168_),
    .A2(_03982_),
    .B(net5670),
    .Y(_04223_));
 NOR2x1_ASAP7_75t_R _26628_ (.A(net6119),
    .B(_04050_),
    .Y(_04224_));
 OAI21x1_ASAP7_75t_R _26629_ (.A1(_04037_),
    .A2(_03950_),
    .B(_04224_),
    .Y(_04225_));
 AO21x1_ASAP7_75t_R _26630_ (.A1(_04223_),
    .A2(_04225_),
    .B(_03925_),
    .Y(_04226_));
 NOR2x1_ASAP7_75t_R _26631_ (.A(_04222_),
    .B(_04226_),
    .Y(_04227_));
 AOI22x1_ASAP7_75t_R _26632_ (.A1(net5106),
    .A2(net4645),
    .B1(_03972_),
    .B2(_03974_),
    .Y(_04228_));
 OAI21x1_ASAP7_75t_R _26633_ (.A1(_03935_),
    .A2(_04228_),
    .B(net6119),
    .Y(_04229_));
 NAND2x1p5_ASAP7_75t_R _26634_ (.A(_03862_),
    .B(net4462),
    .Y(_04230_));
 OA21x2_ASAP7_75t_R _26635_ (.A1(_04117_),
    .A2(net6130),
    .B(net6124),
    .Y(_04231_));
 AOI21x1_ASAP7_75t_R _26636_ (.A1(_04230_),
    .A2(_04231_),
    .B(net5670),
    .Y(_04232_));
 NOR2x1_ASAP7_75t_R _26637_ (.A(net5677),
    .B(net6109),
    .Y(_04233_));
 NOR2x1_ASAP7_75t_R _26638_ (.A(net6122),
    .B(_04233_),
    .Y(_04234_));
 AOI21x1_ASAP7_75t_R _26639_ (.A1(_04234_),
    .A2(_04178_),
    .B(_03880_),
    .Y(_04235_));
 AOI21x1_ASAP7_75t_R _26640_ (.A1(_03839_),
    .A2(_03963_),
    .B(net6109),
    .Y(_04236_));
 INVx1_ASAP7_75t_R _26641_ (.A(_03766_),
    .Y(_04237_));
 AOI21x1_ASAP7_75t_R _26642_ (.A1(_04177_),
    .A2(_04237_),
    .B(net6131),
    .Y(_04238_));
 OAI21x1_ASAP7_75t_R _26643_ (.A1(_04236_),
    .A2(_04238_),
    .B(net6122),
    .Y(_04239_));
 AOI22x1_ASAP7_75t_R _26644_ (.A1(_04229_),
    .A2(_04232_),
    .B1(_04235_),
    .B2(_04239_),
    .Y(_04240_));
 OAI21x1_ASAP7_75t_R _26645_ (.A1(net6108),
    .A2(_04240_),
    .B(net6116),
    .Y(_04241_));
 NOR2x1_ASAP7_75t_R _26646_ (.A(net6124),
    .B(_04000_),
    .Y(_04242_));
 AOI21x1_ASAP7_75t_R _26647_ (.A1(_04078_),
    .A2(_04242_),
    .B(net5670),
    .Y(_04243_));
 OA21x2_ASAP7_75t_R _26648_ (.A1(net6132),
    .A2(_03826_),
    .B(net6124),
    .Y(_04244_));
 NAND2x1_ASAP7_75t_R _26649_ (.A(_04119_),
    .B(_04244_),
    .Y(_04245_));
 AOI21x1_ASAP7_75t_R _26650_ (.A1(_04243_),
    .A2(_04245_),
    .B(net6108),
    .Y(_04246_));
 OAI21x1_ASAP7_75t_R _26651_ (.A1(net4502),
    .A2(_04113_),
    .B(net6136),
    .Y(_04247_));
 NAND2x1_ASAP7_75t_R _26652_ (.A(_03876_),
    .B(_04099_),
    .Y(_04248_));
 AOI21x1_ASAP7_75t_R _26653_ (.A1(_04247_),
    .A2(_04248_),
    .B(net6125),
    .Y(_04249_));
 NAND2x1_ASAP7_75t_R _26654_ (.A(_03911_),
    .B(_03982_),
    .Y(_04250_));
 AOI21x1_ASAP7_75t_R _26655_ (.A1(_03807_),
    .A2(_04250_),
    .B(net6119),
    .Y(_04251_));
 OAI21x1_ASAP7_75t_R _26656_ (.A1(_04249_),
    .A2(_04251_),
    .B(net5670),
    .Y(_04252_));
 AOI21x1_ASAP7_75t_R _26657_ (.A1(_04246_),
    .A2(_04252_),
    .B(net6116),
    .Y(_04253_));
 OAI21x1_ASAP7_75t_R _26658_ (.A1(net4553),
    .A2(_04000_),
    .B(net6130),
    .Y(_04254_));
 NAND2x1_ASAP7_75t_R _26659_ (.A(net5105),
    .B(_04099_),
    .Y(_04255_));
 AOI21x1_ASAP7_75t_R _26660_ (.A1(_04254_),
    .A2(_04255_),
    .B(net6124),
    .Y(_04256_));
 NOR2x1_ASAP7_75t_R _26661_ (.A(net6109),
    .B(net5384),
    .Y(_04257_));
 AOI21x1_ASAP7_75t_R _26662_ (.A1(_03846_),
    .A2(_03849_),
    .B(_04257_),
    .Y(_04258_));
 NOR2x1_ASAP7_75t_R _26663_ (.A(net6122),
    .B(_04258_),
    .Y(_04259_));
 OAI21x1_ASAP7_75t_R _26664_ (.A1(_04256_),
    .A2(_04259_),
    .B(net5670),
    .Y(_04260_));
 AO21x1_ASAP7_75t_R _26665_ (.A1(net5109),
    .A2(net4643),
    .B(net6136),
    .Y(_04261_));
 NAND2x1_ASAP7_75t_R _26666_ (.A(_03902_),
    .B(_04261_),
    .Y(_04262_));
 OA21x2_ASAP7_75t_R _26667_ (.A1(_03839_),
    .A2(net6109),
    .B(net6122),
    .Y(_04263_));
 AO21x1_ASAP7_75t_R _26668_ (.A1(_03963_),
    .A2(_04062_),
    .B(net6131),
    .Y(_04264_));
 AOI21x1_ASAP7_75t_R _26669_ (.A1(_04263_),
    .A2(_04264_),
    .B(net5671),
    .Y(_04265_));
 AOI21x1_ASAP7_75t_R _26670_ (.A1(_04262_),
    .A2(_04265_),
    .B(_03925_),
    .Y(_04266_));
 NAND2x1_ASAP7_75t_R _26671_ (.A(_04260_),
    .B(_04266_),
    .Y(_04267_));
 NAND2x1_ASAP7_75t_R _26672_ (.A(_04253_),
    .B(_04267_),
    .Y(_04268_));
 OAI21x1_ASAP7_75t_R _26673_ (.A1(_04227_),
    .A2(_04241_),
    .B(_04268_),
    .Y(_00117_));
 AOI21x1_ASAP7_75t_R _26674_ (.A1(_04207_),
    .A2(net5109),
    .B(net6112),
    .Y(_04269_));
 AOI21x1_ASAP7_75t_R _26675_ (.A1(_04067_),
    .A2(_04237_),
    .B(net6134),
    .Y(_04270_));
 OAI21x1_ASAP7_75t_R _26676_ (.A1(_04269_),
    .A2(_04270_),
    .B(net6122),
    .Y(_04271_));
 INVx1_ASAP7_75t_R _26677_ (.A(_03933_),
    .Y(_04272_));
 AOI21x1_ASAP7_75t_R _26678_ (.A1(_03846_),
    .A2(_04272_),
    .B(net6112),
    .Y(_04273_));
 NOR2x1_ASAP7_75t_R _26679_ (.A(_04041_),
    .B(_04037_),
    .Y(_04274_));
 OAI21x1_ASAP7_75t_R _26680_ (.A1(_04273_),
    .A2(_04274_),
    .B(net6127),
    .Y(_04275_));
 AOI21x1_ASAP7_75t_R _26681_ (.A1(_04271_),
    .A2(_04275_),
    .B(net5668),
    .Y(_04276_));
 OAI21x1_ASAP7_75t_R _26682_ (.A1(_04015_),
    .A2(_03746_),
    .B(net6121),
    .Y(_04277_));
 NOR2x1_ASAP7_75t_R _26683_ (.A(net6134),
    .B(_03855_),
    .Y(_04278_));
 INVx1_ASAP7_75t_R _26684_ (.A(_04119_),
    .Y(_04279_));
 OAI21x1_ASAP7_75t_R _26685_ (.A1(_04278_),
    .A2(_04279_),
    .B(net6124),
    .Y(_04280_));
 AOI21x1_ASAP7_75t_R _26686_ (.A1(_04277_),
    .A2(_04280_),
    .B(net5671),
    .Y(_04281_));
 NOR3x1_ASAP7_75t_R _26687_ (.A(_04276_),
    .B(_04281_),
    .C(net6116),
    .Y(_04282_));
 NAND2x1_ASAP7_75t_R _26688_ (.A(net5667),
    .B(_04082_),
    .Y(_04283_));
 AO21x1_ASAP7_75t_R _26689_ (.A1(net5388),
    .A2(net4867),
    .B(net6133),
    .Y(_04284_));
 NAND2x1_ASAP7_75t_R _26690_ (.A(net5105),
    .B(_03877_),
    .Y(_04285_));
 AOI21x1_ASAP7_75t_R _26691_ (.A1(_04284_),
    .A2(_04285_),
    .B(net6125),
    .Y(_04286_));
 NOR2x1_ASAP7_75t_R _26692_ (.A(_04283_),
    .B(_04286_),
    .Y(_04287_));
 AOI21x1_ASAP7_75t_R _26693_ (.A1(_01290_),
    .A2(net6128),
    .B(net6118),
    .Y(_04288_));
 NAND2x1_ASAP7_75t_R _26694_ (.A(_04288_),
    .B(_04255_),
    .Y(_04289_));
 AOI21x1_ASAP7_75t_R _26695_ (.A1(_03740_),
    .A2(_03855_),
    .B(net6115),
    .Y(_04290_));
 OAI21x1_ASAP7_75t_R _26696_ (.A1(_03986_),
    .A2(_04290_),
    .B(net6119),
    .Y(_04291_));
 AOI21x1_ASAP7_75t_R _26697_ (.A1(_04289_),
    .A2(_04291_),
    .B(net5667),
    .Y(_04292_));
 OAI21x1_ASAP7_75t_R _26698_ (.A1(_04287_),
    .A2(_04292_),
    .B(net6116),
    .Y(_04293_));
 NAND2x1_ASAP7_75t_R _26699_ (.A(net6108),
    .B(_04293_),
    .Y(_04294_));
 AOI21x1_ASAP7_75t_R _26700_ (.A1(net6109),
    .A2(_04045_),
    .B(net6123),
    .Y(_04295_));
 AO21x1_ASAP7_75t_R _26701_ (.A1(net4645),
    .A2(_03906_),
    .B(net6109),
    .Y(_04296_));
 AOI21x1_ASAP7_75t_R _26702_ (.A1(_04295_),
    .A2(_04296_),
    .B(net5667),
    .Y(_04297_));
 AND2x2_ASAP7_75t_R _26703_ (.A(_01289_),
    .B(_01293_),
    .Y(_04298_));
 OA21x2_ASAP7_75t_R _26704_ (.A1(net6128),
    .A2(_04298_),
    .B(net6123),
    .Y(_04299_));
 OAI21x1_ASAP7_75t_R _26705_ (.A1(net6109),
    .A2(_04208_),
    .B(_04299_),
    .Y(_04300_));
 AOI21x1_ASAP7_75t_R _26706_ (.A1(_04297_),
    .A2(_04300_),
    .B(net6116),
    .Y(_04301_));
 NOR2x1_ASAP7_75t_R _26707_ (.A(_04049_),
    .B(net5387),
    .Y(_04302_));
 OAI21x1_ASAP7_75t_R _26708_ (.A1(_04060_),
    .A2(_04302_),
    .B(net6132),
    .Y(_04303_));
 NAND2x1_ASAP7_75t_R _26709_ (.A(net4732),
    .B(_03849_),
    .Y(_04304_));
 AOI21x1_ASAP7_75t_R _26710_ (.A1(_04303_),
    .A2(_04304_),
    .B(net6123),
    .Y(_04305_));
 NOR2x1_ASAP7_75t_R _26711_ (.A(net4869),
    .B(net5387),
    .Y(_04306_));
 OAI21x1_ASAP7_75t_R _26712_ (.A1(_03804_),
    .A2(_04306_),
    .B(net6129),
    .Y(_04307_));
 NAND2x1_ASAP7_75t_R _26713_ (.A(_03814_),
    .B(_04099_),
    .Y(_04308_));
 AOI21x1_ASAP7_75t_R _26714_ (.A1(_04307_),
    .A2(_04308_),
    .B(net6119),
    .Y(_04309_));
 OAI21x1_ASAP7_75t_R _26715_ (.A1(_04305_),
    .A2(_04309_),
    .B(net5667),
    .Y(_04310_));
 AOI21x1_ASAP7_75t_R _26716_ (.A1(_04301_),
    .A2(_04310_),
    .B(net6108),
    .Y(_04311_));
 OAI21x1_ASAP7_75t_R _26717_ (.A1(_03831_),
    .A2(_04113_),
    .B(net6111),
    .Y(_04312_));
 AOI21x1_ASAP7_75t_R _26718_ (.A1(_04272_),
    .A2(_04157_),
    .B(net6122),
    .Y(_04313_));
 NAND2x1_ASAP7_75t_R _26719_ (.A(_04312_),
    .B(_04313_),
    .Y(_04314_));
 NAND2x1_ASAP7_75t_R _26720_ (.A(_03958_),
    .B(_04157_),
    .Y(_04315_));
 OA21x2_ASAP7_75t_R _26721_ (.A1(_03839_),
    .A2(net6134),
    .B(net6122),
    .Y(_04316_));
 AOI21x1_ASAP7_75t_R _26722_ (.A1(_04315_),
    .A2(_04316_),
    .B(net5671),
    .Y(_04317_));
 AOI21x1_ASAP7_75t_R _26723_ (.A1(_04314_),
    .A2(_04317_),
    .B(_03789_),
    .Y(_04318_));
 AOI21x1_ASAP7_75t_R _26724_ (.A1(_04037_),
    .A2(_04038_),
    .B(_03828_),
    .Y(_04319_));
 AO21x1_ASAP7_75t_R _26725_ (.A1(net4645),
    .A2(net4737),
    .B(net6136),
    .Y(_04320_));
 AO21x1_ASAP7_75t_R _26726_ (.A1(_03810_),
    .A2(_03742_),
    .B(net6113),
    .Y(_04321_));
 AOI21x1_ASAP7_75t_R _26727_ (.A1(_04320_),
    .A2(_04321_),
    .B(net6122),
    .Y(_04322_));
 OAI21x1_ASAP7_75t_R _26728_ (.A1(_04319_),
    .A2(_04322_),
    .B(net5671),
    .Y(_04323_));
 NAND2x1_ASAP7_75t_R _26729_ (.A(_04318_),
    .B(_04323_),
    .Y(_04324_));
 NAND2x1_ASAP7_75t_R _26730_ (.A(_04311_),
    .B(_04324_),
    .Y(_04325_));
 OAI21x1_ASAP7_75t_R _26731_ (.A1(_04282_),
    .A2(_04294_),
    .B(_04325_),
    .Y(_00118_));
 NOR2x1_ASAP7_75t_R _26732_ (.A(net6122),
    .B(_03886_),
    .Y(_04326_));
 NAND2x1_ASAP7_75t_R _26733_ (.A(net5042),
    .B(net6132),
    .Y(_04327_));
 AO21x1_ASAP7_75t_R _26734_ (.A1(_04326_),
    .A2(_04327_),
    .B(_03880_),
    .Y(_04328_));
 NOR3x1_ASAP7_75t_R _26735_ (.A(_03926_),
    .B(_03870_),
    .C(_03834_),
    .Y(_04329_));
 OAI21x1_ASAP7_75t_R _26736_ (.A1(_04328_),
    .A2(_04329_),
    .B(_03925_),
    .Y(_04330_));
 AO21x1_ASAP7_75t_R _26737_ (.A1(net4736),
    .A2(net4642),
    .B(net6128),
    .Y(_04331_));
 NAND2x1_ASAP7_75t_R _26738_ (.A(net6490),
    .B(_03973_),
    .Y(_04332_));
 NAND2x1_ASAP7_75t_R _26739_ (.A(_03797_),
    .B(_03730_),
    .Y(_04333_));
 AO21x1_ASAP7_75t_R _26740_ (.A1(_04332_),
    .A2(_04333_),
    .B(_01293_),
    .Y(_04334_));
 AO21x1_ASAP7_75t_R _26741_ (.A1(_04331_),
    .A2(_04334_),
    .B(net6118),
    .Y(_04335_));
 NAND2x1_ASAP7_75t_R _26742_ (.A(_03855_),
    .B(_03832_),
    .Y(_04336_));
 NAND2x1_ASAP7_75t_R _26743_ (.A(net5105),
    .B(_03945_),
    .Y(_04337_));
 AO21x1_ASAP7_75t_R _26744_ (.A1(_04336_),
    .A2(_04337_),
    .B(net6124),
    .Y(_04338_));
 AOI21x1_ASAP7_75t_R _26745_ (.A1(_04335_),
    .A2(_04338_),
    .B(net5670),
    .Y(_04339_));
 OAI21x1_ASAP7_75t_R _26746_ (.A1(_04330_),
    .A2(_04339_),
    .B(net6116),
    .Y(_04340_));
 AO21x1_ASAP7_75t_R _26747_ (.A1(net5384),
    .A2(net6109),
    .B(_04184_),
    .Y(_04341_));
 AND3x1_ASAP7_75t_R _26748_ (.A(net5106),
    .B(_04051_),
    .C(net6109),
    .Y(_04342_));
 OAI21x1_ASAP7_75t_R _26749_ (.A1(_04181_),
    .A2(_04342_),
    .B(net5672),
    .Y(_04343_));
 AOI21x1_ASAP7_75t_R _26750_ (.A1(net6122),
    .A2(_04341_),
    .B(_04343_),
    .Y(_04344_));
 AO21x1_ASAP7_75t_R _26751_ (.A1(net5387),
    .A2(net5042),
    .B(net6109),
    .Y(_04345_));
 AND2x2_ASAP7_75t_R _26752_ (.A(_04244_),
    .B(_04345_),
    .Y(_04346_));
 AO21x1_ASAP7_75t_R _26753_ (.A1(_03852_),
    .A2(net4737),
    .B(net6136),
    .Y(_04347_));
 AOI21x1_ASAP7_75t_R _26754_ (.A1(_04158_),
    .A2(_04347_),
    .B(net6124),
    .Y(_04348_));
 OAI21x1_ASAP7_75t_R _26755_ (.A1(_04346_),
    .A2(_04348_),
    .B(net5668),
    .Y(_04349_));
 NAND2x1_ASAP7_75t_R _26756_ (.A(net6108),
    .B(_04349_),
    .Y(_04350_));
 NOR2x1_ASAP7_75t_R _26757_ (.A(_04344_),
    .B(_04350_),
    .Y(_04351_));
 AND2x2_ASAP7_75t_R _26758_ (.A(_03945_),
    .B(net4737),
    .Y(_04352_));
 NAND2x1_ASAP7_75t_R _26759_ (.A(net6118),
    .B(_04009_),
    .Y(_04353_));
 AOI21x1_ASAP7_75t_R _26760_ (.A1(_03833_),
    .A2(_03919_),
    .B(net6120),
    .Y(_04354_));
 AOI21x1_ASAP7_75t_R _26761_ (.A1(_04308_),
    .A2(_04354_),
    .B(net5672),
    .Y(_04355_));
 OAI21x1_ASAP7_75t_R _26762_ (.A1(_04352_),
    .A2(_04353_),
    .B(_04355_),
    .Y(_04356_));
 AOI21x1_ASAP7_75t_R _26763_ (.A1(net6111),
    .A2(_03814_),
    .B(net6120),
    .Y(_04357_));
 AOI21x1_ASAP7_75t_R _26764_ (.A1(_04357_),
    .A2(_04285_),
    .B(net5667),
    .Y(_04358_));
 NAND2x1_ASAP7_75t_R _26765_ (.A(_03876_),
    .B(_03945_),
    .Y(_04359_));
 OAI21x1_ASAP7_75t_R _26766_ (.A1(net6111),
    .A2(_03840_),
    .B(net6118),
    .Y(_04360_));
 NOR3x1_ASAP7_75t_R _26767_ (.A(net6111),
    .B(net5386),
    .C(net4870),
    .Y(_04361_));
 NOR2x1_ASAP7_75t_R _26768_ (.A(_04360_),
    .B(_04361_),
    .Y(_04362_));
 NAND2x1_ASAP7_75t_R _26769_ (.A(_04359_),
    .B(_04362_),
    .Y(_04363_));
 AOI21x1_ASAP7_75t_R _26770_ (.A1(_04358_),
    .A2(_04363_),
    .B(_03925_),
    .Y(_04364_));
 NAND2x1_ASAP7_75t_R _26771_ (.A(_04356_),
    .B(_04364_),
    .Y(_04365_));
 OAI21x1_ASAP7_75t_R _26772_ (.A1(_03826_),
    .A2(_03871_),
    .B(net6128),
    .Y(_04366_));
 OAI21x1_ASAP7_75t_R _26773_ (.A1(_04045_),
    .A2(_04306_),
    .B(net6109),
    .Y(_04367_));
 AOI21x1_ASAP7_75t_R _26774_ (.A1(_04366_),
    .A2(_04367_),
    .B(net6119),
    .Y(_04368_));
 NAND2x1_ASAP7_75t_R _26775_ (.A(_04051_),
    .B(_03916_),
    .Y(_04369_));
 AOI21x1_ASAP7_75t_R _26776_ (.A1(_04114_),
    .A2(_04369_),
    .B(net6123),
    .Y(_04370_));
 OAI21x1_ASAP7_75t_R _26777_ (.A1(_04368_),
    .A2(_04370_),
    .B(net5672),
    .Y(_04371_));
 NOR2x1_ASAP7_75t_R _26778_ (.A(net6127),
    .B(_03975_),
    .Y(_04372_));
 OAI21x1_ASAP7_75t_R _26779_ (.A1(net6109),
    .A2(_04208_),
    .B(_04372_),
    .Y(_04373_));
 AOI21x1_ASAP7_75t_R _26780_ (.A1(net5388),
    .A2(_04233_),
    .B(_04045_),
    .Y(_04374_));
 AOI21x1_ASAP7_75t_R _26781_ (.A1(_04326_),
    .A2(_04374_),
    .B(net5672),
    .Y(_04375_));
 AOI21x1_ASAP7_75t_R _26782_ (.A1(_04373_),
    .A2(_04375_),
    .B(net6108),
    .Y(_04376_));
 AOI21x1_ASAP7_75t_R _26783_ (.A1(_04371_),
    .A2(_04376_),
    .B(net6116),
    .Y(_04377_));
 NAND2x1_ASAP7_75t_R _26784_ (.A(_04365_),
    .B(_04377_),
    .Y(_04378_));
 OAI21x1_ASAP7_75t_R _26785_ (.A1(_04340_),
    .A2(_04351_),
    .B(_04378_),
    .Y(_00119_));
 NOR2x1_ASAP7_75t_R _26786_ (.A(net6660),
    .B(_00477_),
    .Y(_04379_));
 XOR2x2_ASAP7_75t_R _26787_ (.A(_00695_),
    .B(_00569_),
    .Y(_04380_));
 XOR2x2_ASAP7_75t_R _26788_ (.A(_04380_),
    .B(_12818_),
    .Y(_04381_));
 XOR2x2_ASAP7_75t_R _26789_ (.A(_12853_),
    .B(_01589_),
    .Y(_04382_));
 NAND2x1_ASAP7_75t_R _26790_ (.A(_04381_),
    .B(_04382_),
    .Y(_04383_));
 XOR2x2_ASAP7_75t_R _26791_ (.A(_04380_),
    .B(net6545),
    .Y(_04384_));
 XOR2x2_ASAP7_75t_R _26792_ (.A(_12851_),
    .B(_01589_),
    .Y(_04385_));
 NAND2x1_ASAP7_75t_R _26793_ (.A(_04384_),
    .B(_04385_),
    .Y(_04386_));
 AOI21x1_ASAP7_75t_R _26794_ (.A1(_04383_),
    .A2(_04386_),
    .B(net6457),
    .Y(_04387_));
 OAI21x1_ASAP7_75t_R _26795_ (.A1(_04379_),
    .A2(net6348),
    .B(net6472),
    .Y(_04388_));
 AND2x2_ASAP7_75t_R _26796_ (.A(net6459),
    .B(_00477_),
    .Y(_04389_));
 NAND2x1_ASAP7_75t_R _26797_ (.A(_04384_),
    .B(_04382_),
    .Y(_04390_));
 NAND2x1_ASAP7_75t_R _26798_ (.A(_04381_),
    .B(_04385_),
    .Y(_04391_));
 AOI21x1_ASAP7_75t_R _26799_ (.A1(_04390_),
    .A2(_04391_),
    .B(net6457),
    .Y(_04392_));
 INVx1_ASAP7_75t_R _26800_ (.A(net6472),
    .Y(_04393_));
 OAI21x1_ASAP7_75t_R _26801_ (.A1(_04389_),
    .A2(net6347),
    .B(_04393_),
    .Y(_04394_));
 NAND2x1p5_ASAP7_75t_R _26802_ (.A(_04388_),
    .B(_04394_),
    .Y(_01306_));
 NOR2x1_ASAP7_75t_R _26803_ (.A(net6673),
    .B(_00478_),
    .Y(_04395_));
 XOR2x2_ASAP7_75t_R _26804_ (.A(_00631_),
    .B(_00599_),
    .Y(_04396_));
 NAND2x1_ASAP7_75t_R _26805_ (.A(_01773_),
    .B(net6396),
    .Y(_04397_));
 OR2x2_ASAP7_75t_R _26806_ (.A(_01773_),
    .B(_04396_),
    .Y(_04398_));
 INVx1_ASAP7_75t_R _26807_ (.A(_04380_),
    .Y(_04399_));
 AOI21x1_ASAP7_75t_R _26808_ (.A1(_04397_),
    .A2(_04398_),
    .B(_04399_),
    .Y(_04400_));
 XOR2x2_ASAP7_75t_R _26809_ (.A(net6571),
    .B(_04396_),
    .Y(_04401_));
 NOR2x1p5_ASAP7_75t_R _26810_ (.A(_04380_),
    .B(_04401_),
    .Y(_04402_));
 OAI21x1_ASAP7_75t_R _26811_ (.A1(_04402_),
    .A2(_04400_),
    .B(net6664),
    .Y(_04403_));
 INVx2_ASAP7_75t_R _26812_ (.A(_04403_),
    .Y(_04404_));
 OAI21x1_ASAP7_75t_R _26813_ (.A1(net6397),
    .A2(_04404_),
    .B(_00964_),
    .Y(_04405_));
 INVx1_ASAP7_75t_R _26814_ (.A(_04395_),
    .Y(_04406_));
 NAND3x1_ASAP7_75t_R _26815_ (.A(net6346),
    .B(_08947_),
    .C(_04406_),
    .Y(_04407_));
 NAND2x1_ASAP7_75t_R _26816_ (.A(_04405_),
    .B(_04407_),
    .Y(_01303_));
 NOR2x1_ASAP7_75t_R _26817_ (.A(net6660),
    .B(_00479_),
    .Y(_04408_));
 INVx1_ASAP7_75t_R _26818_ (.A(_04408_),
    .Y(_04409_));
 XOR2x2_ASAP7_75t_R _26819_ (.A(_00601_),
    .B(_00633_),
    .Y(_04410_));
 XOR2x2_ASAP7_75t_R _26820_ (.A(net6405),
    .B(net6544),
    .Y(_04411_));
 NOR2x1_ASAP7_75t_R _26821_ (.A(net6395),
    .B(_04411_),
    .Y(_04412_));
 INVx1_ASAP7_75t_R _26822_ (.A(net6544),
    .Y(_04413_));
 NOR2x1_ASAP7_75t_R _26823_ (.A(_04413_),
    .B(net6405),
    .Y(_04414_));
 INVx1_ASAP7_75t_R _26824_ (.A(net6405),
    .Y(_04415_));
 NOR2x1_ASAP7_75t_R _26825_ (.A(net6544),
    .B(_04415_),
    .Y(_04416_));
 OAI21x1_ASAP7_75t_R _26826_ (.A1(_04414_),
    .A2(_04416_),
    .B(net6395),
    .Y(_04417_));
 INVx1_ASAP7_75t_R _26827_ (.A(_04417_),
    .Y(_04418_));
 OAI21x1_ASAP7_75t_R _26828_ (.A1(_04412_),
    .A2(_04418_),
    .B(net6660),
    .Y(_04419_));
 INVx1_ASAP7_75t_R _26829_ (.A(net6476),
    .Y(_04420_));
 AOI21x1_ASAP7_75t_R _26830_ (.A1(_04409_),
    .A2(_04419_),
    .B(_04420_),
    .Y(_04421_));
 NAND2x1_ASAP7_75t_R _26831_ (.A(_00479_),
    .B(net6459),
    .Y(_04422_));
 INVx1_ASAP7_75t_R _26832_ (.A(_04410_),
    .Y(_04423_));
 XOR2x2_ASAP7_75t_R _26833_ (.A(net6405),
    .B(_04413_),
    .Y(_04424_));
 NAND2x1_ASAP7_75t_R _26834_ (.A(_04423_),
    .B(_04424_),
    .Y(_04425_));
 NAND3x1_ASAP7_75t_R _26835_ (.A(_04425_),
    .B(net6660),
    .C(_04417_),
    .Y(_04426_));
 AOI21x1_ASAP7_75t_R _26836_ (.A1(_04422_),
    .A2(_04426_),
    .B(net6476),
    .Y(_04427_));
 NOR2x2_ASAP7_75t_R _26837_ (.A(_04421_),
    .B(_04427_),
    .Y(_04428_));
 OAI21x1_ASAP7_75t_R _26839_ (.A1(_04379_),
    .A2(_04387_),
    .B(_04393_),
    .Y(_04429_));
 OAI21x1_ASAP7_75t_R _26840_ (.A1(_04389_),
    .A2(_04392_),
    .B(net6472),
    .Y(_04430_));
 NAND2x1_ASAP7_75t_R _26841_ (.A(_04429_),
    .B(_04430_),
    .Y(_04431_));
 AOI21x1_ASAP7_75t_R _26843_ (.A1(_04409_),
    .A2(_04419_),
    .B(net6476),
    .Y(_04432_));
 AOI21x1_ASAP7_75t_R _26844_ (.A1(_04422_),
    .A2(_04426_),
    .B(_04420_),
    .Y(_04433_));
 NOR2x1_ASAP7_75t_R _26845_ (.A(_04432_),
    .B(_04433_),
    .Y(_04434_));
 XNOR2x2_ASAP7_75t_R _26848_ (.A(_00698_),
    .B(_01659_),
    .Y(_04436_));
 XNOR2x2_ASAP7_75t_R _26849_ (.A(net6542),
    .B(net6544),
    .Y(_04437_));
 XOR2x2_ASAP7_75t_R _26850_ (.A(_00602_),
    .B(_00634_),
    .Y(_04438_));
 XOR2x2_ASAP7_75t_R _26851_ (.A(_04437_),
    .B(_04438_),
    .Y(_04439_));
 NOR2x1_ASAP7_75t_R _26852_ (.A(_04436_),
    .B(_04439_),
    .Y(_04440_));
 AO21x1_ASAP7_75t_R _26853_ (.A1(_04439_),
    .A2(_04436_),
    .B(net6458),
    .Y(_04441_));
 NAND2x1_ASAP7_75t_R _26854_ (.A(_00554_),
    .B(net6458),
    .Y(_04442_));
 OAI21x1_ASAP7_75t_R _26855_ (.A1(_04440_),
    .A2(_04441_),
    .B(_04442_),
    .Y(_04443_));
 XOR2x2_ASAP7_75t_R _26856_ (.A(_04443_),
    .B(_00936_),
    .Y(_04444_));
 OAI21x1_ASAP7_75t_R _26859_ (.A1(net5381),
    .A2(net5662),
    .B(_01301_),
    .Y(_04447_));
 XNOR2x2_ASAP7_75t_R _26860_ (.A(net6542),
    .B(_00698_),
    .Y(_04448_));
 XOR2x2_ASAP7_75t_R _26861_ (.A(_04448_),
    .B(_12956_),
    .Y(_04449_));
 XOR2x2_ASAP7_75t_R _26862_ (.A(_01643_),
    .B(net6543),
    .Y(_04450_));
 XOR2x2_ASAP7_75t_R _26863_ (.A(_04449_),
    .B(_04450_),
    .Y(_04451_));
 NAND2x1_ASAP7_75t_R _26864_ (.A(net6658),
    .B(_04451_),
    .Y(_04452_));
 OR2x2_ASAP7_75t_R _26865_ (.A(net6658),
    .B(_00548_),
    .Y(_04453_));
 NAND3x1_ASAP7_75t_R _26866_ (.A(_04452_),
    .B(_00937_),
    .C(_04453_),
    .Y(_04454_));
 AO21x1_ASAP7_75t_R _26867_ (.A1(_04452_),
    .A2(_04453_),
    .B(_00937_),
    .Y(_04455_));
 NAND2x1_ASAP7_75t_R _26868_ (.A(_04454_),
    .B(_04455_),
    .Y(_04456_));
 AOI21x1_ASAP7_75t_R _26870_ (.A1(net6106),
    .A2(_04447_),
    .B(net5661),
    .Y(_04458_));
 NAND2x1_ASAP7_75t_R _26871_ (.A(net5663),
    .B(net5104),
    .Y(_04459_));
 OAI21x1_ASAP7_75t_R _26872_ (.A1(net5382),
    .A2(net5664),
    .B(_01301_),
    .Y(_04460_));
 AO21x1_ASAP7_75t_R _26875_ (.A1(_04459_),
    .A2(net4730),
    .B(net6106),
    .Y(_04463_));
 XOR2x2_ASAP7_75t_R _26876_ (.A(_12928_),
    .B(_00700_),
    .Y(_04464_));
 XOR2x2_ASAP7_75t_R _26877_ (.A(_04464_),
    .B(_12907_),
    .Y(_04465_));
 NOR2x1_ASAP7_75t_R _26878_ (.A(net6658),
    .B(_00547_),
    .Y(_04466_));
 AO21x1_ASAP7_75t_R _26879_ (.A1(_04465_),
    .A2(net6658),
    .B(_04466_),
    .Y(_04467_));
 XOR2x2_ASAP7_75t_R _26880_ (.A(_04467_),
    .B(_00938_),
    .Y(_04468_));
 INVx1_ASAP7_75t_R _26881_ (.A(_04468_),
    .Y(_04469_));
 AOI21x1_ASAP7_75t_R _26883_ (.A1(net4552),
    .A2(_04463_),
    .B(net5658),
    .Y(_04471_));
 NAND3x1_ASAP7_75t_R _26884_ (.A(_04419_),
    .B(net6476),
    .C(_04409_),
    .Y(_04472_));
 AOI21x1_ASAP7_75t_R _26886_ (.A1(_04417_),
    .A2(_04425_),
    .B(net6459),
    .Y(_04474_));
 OAI21x1_ASAP7_75t_R _26887_ (.A1(_04408_),
    .A2(_04474_),
    .B(_04420_),
    .Y(_04475_));
 AO21x1_ASAP7_75t_R _26889_ (.A1(net5380),
    .A2(net5656),
    .B(_01300_),
    .Y(_04477_));
 NAND2x1p5_ASAP7_75t_R _26890_ (.A(net6105),
    .B(_04460_),
    .Y(_04478_));
 INVx1_ASAP7_75t_R _26891_ (.A(_04478_),
    .Y(_04479_));
 NAND2x1_ASAP7_75t_R _26892_ (.A(_04477_),
    .B(net4461),
    .Y(_04480_));
 OAI21x1_ASAP7_75t_R _26893_ (.A1(net5382),
    .A2(net5664),
    .B(_01300_),
    .Y(_04481_));
 INVx1_ASAP7_75t_R _26894_ (.A(_04481_),
    .Y(_04482_));
 OA21x2_ASAP7_75t_R _26895_ (.A1(net5662),
    .A2(net5381),
    .B(_01304_),
    .Y(_04483_));
 XOR2x2_ASAP7_75t_R _26897_ (.A(_04443_),
    .B(_08963_),
    .Y(_04485_));
 OAI21x1_ASAP7_75t_R _26900_ (.A1(_04482_),
    .A2(net4862),
    .B(net6092),
    .Y(_04488_));
 INVx1_ASAP7_75t_R _26901_ (.A(_00937_),
    .Y(_04489_));
 NAND3x1_ASAP7_75t_R _26902_ (.A(_04452_),
    .B(_04489_),
    .C(_04453_),
    .Y(_04490_));
 AO21x1_ASAP7_75t_R _26903_ (.A1(_04452_),
    .A2(_04453_),
    .B(_04489_),
    .Y(_04491_));
 NAND2x1_ASAP7_75t_R _26904_ (.A(_04490_),
    .B(_04491_),
    .Y(_04492_));
 AO21x1_ASAP7_75t_R _26907_ (.A1(_04480_),
    .A2(_04488_),
    .B(net5653),
    .Y(_04495_));
 NAND2x1_ASAP7_75t_R _26908_ (.A(_04471_),
    .B(_04495_),
    .Y(_04496_));
 AOI21x1_ASAP7_75t_R _26909_ (.A1(net5383),
    .A2(net5101),
    .B(net6107),
    .Y(_04497_));
 OAI21x1_ASAP7_75t_R _26910_ (.A1(_04404_),
    .A2(net6397),
    .B(_08947_),
    .Y(_04498_));
 NAND3x1_ASAP7_75t_R _26911_ (.A(_04403_),
    .B(_00964_),
    .C(_04406_),
    .Y(_04499_));
 NAND2x1p5_ASAP7_75t_R _26912_ (.A(_04499_),
    .B(_04498_),
    .Y(_04500_));
 NAND2x1_ASAP7_75t_R _26913_ (.A(net5663),
    .B(net5378),
    .Y(_04501_));
 AND2x2_ASAP7_75t_R _26914_ (.A(_04497_),
    .B(_04501_),
    .Y(_04502_));
 NOR2x1_ASAP7_75t_R _26917_ (.A(net5104),
    .B(net5378),
    .Y(_04504_));
 NOR2x1_ASAP7_75t_R _26918_ (.A(net5666),
    .B(net5383),
    .Y(_04505_));
 OA21x2_ASAP7_75t_R _26919_ (.A1(_04504_),
    .A2(_04505_),
    .B(net6107),
    .Y(_04506_));
 OAI21x1_ASAP7_75t_R _26922_ (.A1(_04502_),
    .A2(_04506_),
    .B(net5653),
    .Y(_04509_));
 INVx1_ASAP7_75t_R _26925_ (.A(_01309_),
    .Y(_04512_));
 AO21x1_ASAP7_75t_R _26926_ (.A1(net5380),
    .A2(net5656),
    .B(_04512_),
    .Y(_04513_));
 INVx1_ASAP7_75t_R _26927_ (.A(_01301_),
    .Y(_04514_));
 OA21x2_ASAP7_75t_R _26928_ (.A1(net5664),
    .A2(net5382),
    .B(_04514_),
    .Y(_04515_));
 INVx1_ASAP7_75t_R _26929_ (.A(_04515_),
    .Y(_04516_));
 AOI21x1_ASAP7_75t_R _26932_ (.A1(_04513_),
    .A2(net4459),
    .B(net6106),
    .Y(_04519_));
 INVx1_ASAP7_75t_R _26933_ (.A(_01300_),
    .Y(_04520_));
 AO21x1_ASAP7_75t_R _26934_ (.A1(net5380),
    .A2(net5656),
    .B(_04520_),
    .Y(_04521_));
 OA21x2_ASAP7_75t_R _26935_ (.A1(net5664),
    .A2(net5382),
    .B(net5038),
    .Y(_04522_));
 INVx1_ASAP7_75t_R _26936_ (.A(_04522_),
    .Y(_04523_));
 AOI21x1_ASAP7_75t_R _26939_ (.A1(_04521_),
    .A2(_04523_),
    .B(net6093),
    .Y(_04526_));
 OAI21x1_ASAP7_75t_R _26941_ (.A1(_04519_),
    .A2(_04526_),
    .B(net5661),
    .Y(_04528_));
 NAND3x1_ASAP7_75t_R _26942_ (.A(_04509_),
    .B(net5658),
    .C(_04528_),
    .Y(_04529_));
 XOR2x2_ASAP7_75t_R _26943_ (.A(_00700_),
    .B(_00701_),
    .Y(_04530_));
 XOR2x2_ASAP7_75t_R _26944_ (.A(_04530_),
    .B(_00668_),
    .Y(_04531_));
 XNOR2x2_ASAP7_75t_R _26945_ (.A(_13006_),
    .B(_04531_),
    .Y(_04532_));
 NOR2x1_ASAP7_75t_R _26946_ (.A(net6658),
    .B(_00546_),
    .Y(_04533_));
 AO21x1_ASAP7_75t_R _26947_ (.A1(_04532_),
    .A2(net6658),
    .B(_04533_),
    .Y(_04534_));
 XOR2x2_ASAP7_75t_R _26948_ (.A(_04534_),
    .B(_00939_),
    .Y(_04535_));
 INVx1_ASAP7_75t_R _26949_ (.A(_04535_),
    .Y(_04536_));
 AOI21x1_ASAP7_75t_R _26951_ (.A1(_04496_),
    .A2(_04529_),
    .B(net5644),
    .Y(_04538_));
 INVx1_ASAP7_75t_R _26952_ (.A(_01310_),
    .Y(_04539_));
 AO21x1_ASAP7_75t_R _26953_ (.A1(net5380),
    .A2(net5656),
    .B(_04539_),
    .Y(_04540_));
 NOR2x1_ASAP7_75t_R _26954_ (.A(net5103),
    .B(net5383),
    .Y(_04541_));
 INVx1_ASAP7_75t_R _26955_ (.A(_01307_),
    .Y(_04542_));
 AO21x1_ASAP7_75t_R _26956_ (.A1(net5103),
    .A2(net4861),
    .B(net6102),
    .Y(_04543_));
 OAI21x1_ASAP7_75t_R _26957_ (.A1(_04541_),
    .A2(_04543_),
    .B(net5646),
    .Y(_04544_));
 AOI21x1_ASAP7_75t_R _26958_ (.A1(net4461),
    .A2(_04540_),
    .B(_04544_),
    .Y(_04545_));
 AOI21x1_ASAP7_75t_R _26959_ (.A1(net5034),
    .A2(net5101),
    .B(net6099),
    .Y(_04546_));
 AO21x1_ASAP7_75t_R _26960_ (.A1(net5380),
    .A2(net5656),
    .B(net5036),
    .Y(_04547_));
 AOI21x1_ASAP7_75t_R _26961_ (.A1(net5379),
    .A2(net5103),
    .B(net6105),
    .Y(_04548_));
 AO21x1_ASAP7_75t_R _26962_ (.A1(net4860),
    .A2(_04547_),
    .B(_04548_),
    .Y(_04549_));
 OAI21x1_ASAP7_75t_R _26963_ (.A1(net5647),
    .A2(_04549_),
    .B(net5657),
    .Y(_04550_));
 OAI21x1_ASAP7_75t_R _26964_ (.A1(_04545_),
    .A2(_04550_),
    .B(net5644),
    .Y(_04551_));
 AOI21x1_ASAP7_75t_R _26965_ (.A1(net5379),
    .A2(net5103),
    .B(net6099),
    .Y(_04552_));
 NAND3x1_ASAP7_75t_R _26966_ (.A(_04419_),
    .B(_04420_),
    .C(_04409_),
    .Y(_04553_));
 INVx2_ASAP7_75t_R _26967_ (.A(net5382),
    .Y(_04554_));
 AO21x1_ASAP7_75t_R _26968_ (.A1(_04553_),
    .A2(_04554_),
    .B(_04539_),
    .Y(_04555_));
 NAND2x1_ASAP7_75t_R _26969_ (.A(net5663),
    .B(_04434_),
    .Y(_04556_));
 AND3x1_ASAP7_75t_R _26971_ (.A(net4858),
    .B(_04547_),
    .C(net6096),
    .Y(_04558_));
 AOI21x1_ASAP7_75t_R _26972_ (.A1(net4859),
    .A2(net4641),
    .B(_04558_),
    .Y(_04559_));
 AO21x1_ASAP7_75t_R _26973_ (.A1(_04553_),
    .A2(_04554_),
    .B(_01309_),
    .Y(_04560_));
 AND2x2_ASAP7_75t_R _26974_ (.A(net4859),
    .B(_04560_),
    .Y(_04561_));
 NOR2x1_ASAP7_75t_R _26976_ (.A(net5666),
    .B(net5102),
    .Y(_04563_));
 NAND2x1_ASAP7_75t_R _26977_ (.A(net6094),
    .B(_04563_),
    .Y(_04564_));
 INVx1_ASAP7_75t_R _26978_ (.A(_01302_),
    .Y(_04565_));
 OAI21x1_ASAP7_75t_R _26979_ (.A1(net5382),
    .A2(net5664),
    .B(_04565_),
    .Y(_04566_));
 OA21x2_ASAP7_75t_R _26980_ (.A1(net6107),
    .A2(_04566_),
    .B(net5661),
    .Y(_04567_));
 NAND2x1_ASAP7_75t_R _26981_ (.A(_04564_),
    .B(_04567_),
    .Y(_04568_));
 OAI21x1_ASAP7_75t_R _26984_ (.A1(_04561_),
    .A2(_04568_),
    .B(net6100),
    .Y(_04571_));
 AOI21x1_ASAP7_75t_R _26985_ (.A1(net5647),
    .A2(_04559_),
    .B(_04571_),
    .Y(_04572_));
 XOR2x2_ASAP7_75t_R _26986_ (.A(net6424),
    .B(_01727_),
    .Y(_04573_));
 INVx1_ASAP7_75t_R _26987_ (.A(net6542),
    .Y(_04574_));
 XOR2x2_ASAP7_75t_R _26988_ (.A(_04573_),
    .B(_04574_),
    .Y(_04575_));
 NOR2x1_ASAP7_75t_R _26989_ (.A(net6658),
    .B(_00545_),
    .Y(_04576_));
 AO21x1_ASAP7_75t_R _26990_ (.A1(_04575_),
    .A2(net6658),
    .B(_04576_),
    .Y(_04577_));
 XOR2x2_ASAP7_75t_R _26991_ (.A(_04577_),
    .B(_00940_),
    .Y(_04578_));
 OAI21x1_ASAP7_75t_R _26993_ (.A1(_04551_),
    .A2(_04572_),
    .B(net6088),
    .Y(_04580_));
 AOI21x1_ASAP7_75t_R _26995_ (.A1(_04560_),
    .A2(_04552_),
    .B(net5649),
    .Y(_04582_));
 INVx1_ASAP7_75t_R _26996_ (.A(_04582_),
    .Y(_04583_));
 AOI21x1_ASAP7_75t_R _26997_ (.A1(_04554_),
    .A2(_04553_),
    .B(_01305_),
    .Y(_04584_));
 INVx2_ASAP7_75t_R _26998_ (.A(_04584_),
    .Y(_04585_));
 OA21x2_ASAP7_75t_R _27000_ (.A1(_04585_),
    .A2(net6103),
    .B(net5649),
    .Y(_04587_));
 NAND2x1_ASAP7_75t_R _27001_ (.A(net4551),
    .B(_04587_),
    .Y(_04588_));
 INVx1_ASAP7_75t_R _27002_ (.A(_01308_),
    .Y(_04589_));
 OAI21x1_ASAP7_75t_R _27003_ (.A1(net5381),
    .A2(net5662),
    .B(_04589_),
    .Y(_04590_));
 INVx1_ASAP7_75t_R _27004_ (.A(_04590_),
    .Y(_04591_));
 AO21x1_ASAP7_75t_R _27005_ (.A1(_04591_),
    .A2(net6097),
    .B(net5657),
    .Y(_04592_));
 AOI21x1_ASAP7_75t_R _27006_ (.A1(_04583_),
    .A2(_04588_),
    .B(_04592_),
    .Y(_04593_));
 NOR2x1_ASAP7_75t_R _27007_ (.A(net5661),
    .B(net4860),
    .Y(_04594_));
 AO21x1_ASAP7_75t_R _27008_ (.A1(_04521_),
    .A2(_04566_),
    .B(net6106),
    .Y(_04595_));
 NAND2x1_ASAP7_75t_R _27009_ (.A(_04594_),
    .B(_04595_),
    .Y(_04596_));
 AOI21x1_ASAP7_75t_R _27011_ (.A1(_04447_),
    .A2(net4858),
    .B(net6107),
    .Y(_04598_));
 INVx1_ASAP7_75t_R _27012_ (.A(_04598_),
    .Y(_04599_));
 AO21x1_ASAP7_75t_R _27013_ (.A1(net5380),
    .A2(net5656),
    .B(net5038),
    .Y(_04600_));
 AOI21x1_ASAP7_75t_R _27014_ (.A1(net5378),
    .A2(net5101),
    .B(net6094),
    .Y(_04601_));
 AOI21x1_ASAP7_75t_R _27015_ (.A1(_04600_),
    .A2(_04601_),
    .B(net5652),
    .Y(_04602_));
 NAND2x1_ASAP7_75t_R _27016_ (.A(_04599_),
    .B(_04602_),
    .Y(_04603_));
 AOI21x1_ASAP7_75t_R _27017_ (.A1(_04596_),
    .A2(_04603_),
    .B(net6101),
    .Y(_04604_));
 OAI21x1_ASAP7_75t_R _27018_ (.A1(_04593_),
    .A2(_04604_),
    .B(net5644),
    .Y(_04605_));
 OAI21x1_ASAP7_75t_R _27019_ (.A1(net5382),
    .A2(net5664),
    .B(net5036),
    .Y(_04606_));
 NAND2x1_ASAP7_75t_R _27020_ (.A(_04590_),
    .B(_04606_),
    .Y(_04607_));
 AOI21x1_ASAP7_75t_R _27021_ (.A1(net6098),
    .A2(_04607_),
    .B(net5649),
    .Y(_04608_));
 INVx1_ASAP7_75t_R _27022_ (.A(_04608_),
    .Y(_04609_));
 AO21x1_ASAP7_75t_R _27023_ (.A1(net5380),
    .A2(net5656),
    .B(net5039),
    .Y(_04610_));
 AOI22x1_ASAP7_75t_R _27024_ (.A1(net5380),
    .A2(net5656),
    .B1(_04407_),
    .B2(_04405_),
    .Y(_04611_));
 OAI21x1_ASAP7_75t_R _27026_ (.A1(_04482_),
    .A2(_04611_),
    .B(net6102),
    .Y(_04613_));
 OAI21x1_ASAP7_75t_R _27027_ (.A1(net6107),
    .A2(net4853),
    .B(_04613_),
    .Y(_04614_));
 INVx1_ASAP7_75t_R _27028_ (.A(_01318_),
    .Y(_04615_));
 OAI21x1_ASAP7_75t_R _27029_ (.A1(net5381),
    .A2(net5662),
    .B(_04514_),
    .Y(_04616_));
 NAND2x1p5_ASAP7_75t_R _27030_ (.A(_04616_),
    .B(net6092),
    .Y(_04617_));
 OAI21x1_ASAP7_75t_R _27031_ (.A1(_04615_),
    .A2(net6092),
    .B(_04617_),
    .Y(_04618_));
 AOI21x1_ASAP7_75t_R _27032_ (.A1(net5653),
    .A2(_04618_),
    .B(net5658),
    .Y(_04619_));
 OAI21x1_ASAP7_75t_R _27033_ (.A1(_04609_),
    .A2(_04614_),
    .B(_04619_),
    .Y(_04620_));
 AOI21x1_ASAP7_75t_R _27034_ (.A1(_04554_),
    .A2(_04553_),
    .B(_04542_),
    .Y(_04621_));
 OAI21x1_ASAP7_75t_R _27035_ (.A1(_04621_),
    .A2(net4862),
    .B(net6094),
    .Y(_04622_));
 OA21x2_ASAP7_75t_R _27036_ (.A1(net6094),
    .A2(_04566_),
    .B(net5655),
    .Y(_04623_));
 AOI21x1_ASAP7_75t_R _27038_ (.A1(_04622_),
    .A2(_04623_),
    .B(net6101),
    .Y(_04625_));
 OR2x2_ASAP7_75t_R _27039_ (.A(net6102),
    .B(_04566_),
    .Y(_04626_));
 AOI21x1_ASAP7_75t_R _27040_ (.A1(_04475_),
    .A2(_04472_),
    .B(_01305_),
    .Y(_04627_));
 OAI21x1_ASAP7_75t_R _27041_ (.A1(net4852),
    .A2(_04621_),
    .B(net6102),
    .Y(_04628_));
 NAND3x1_ASAP7_75t_R _27043_ (.A(_04626_),
    .B(_04628_),
    .C(net5660),
    .Y(_04630_));
 AOI21x1_ASAP7_75t_R _27044_ (.A1(_04625_),
    .A2(_04630_),
    .B(_04536_),
    .Y(_04631_));
 AOI21x1_ASAP7_75t_R _27045_ (.A1(_04620_),
    .A2(_04631_),
    .B(net6088),
    .Y(_04632_));
 NAND2x1_ASAP7_75t_R _27046_ (.A(_04632_),
    .B(_04605_),
    .Y(_04633_));
 OAI21x1_ASAP7_75t_R _27047_ (.A1(_04538_),
    .A2(_04580_),
    .B(_04633_),
    .Y(_00120_));
 AOI21x1_ASAP7_75t_R _27048_ (.A1(_04512_),
    .A2(net5103),
    .B(net6099),
    .Y(_04634_));
 INVx1_ASAP7_75t_R _27049_ (.A(_04634_),
    .Y(_04635_));
 NOR2x1_ASAP7_75t_R _27051_ (.A(net5034),
    .B(net5103),
    .Y(_04637_));
 AOI21x1_ASAP7_75t_R _27052_ (.A1(net6096),
    .A2(_04637_),
    .B(net5648),
    .Y(_04638_));
 OAI21x1_ASAP7_75t_R _27053_ (.A1(net4550),
    .A2(_04635_),
    .B(_04638_),
    .Y(_04639_));
 OAI21x1_ASAP7_75t_R _27054_ (.A1(net5382),
    .A2(net5664),
    .B(_01309_),
    .Y(_04640_));
 INVx1_ASAP7_75t_R _27055_ (.A(_04640_),
    .Y(_04641_));
 NAND2x1_ASAP7_75t_R _27056_ (.A(net6095),
    .B(net4635),
    .Y(_04642_));
 AOI21x1_ASAP7_75t_R _27057_ (.A1(net5032),
    .A2(net5103),
    .B(net6099),
    .Y(_04643_));
 AOI21x1_ASAP7_75t_R _27058_ (.A1(net4858),
    .A2(_04643_),
    .B(net5660),
    .Y(_04644_));
 NAND2x1_ASAP7_75t_R _27059_ (.A(_04642_),
    .B(_04644_),
    .Y(_04645_));
 AOI21x1_ASAP7_75t_R _27060_ (.A1(_04639_),
    .A2(_04645_),
    .B(net6100),
    .Y(_04646_));
 NOR2x1_ASAP7_75t_R _27061_ (.A(_04591_),
    .B(net4551),
    .Y(_04647_));
 OAI21x1_ASAP7_75t_R _27062_ (.A1(net5101),
    .A2(net5379),
    .B(net6099),
    .Y(_04648_));
 OAI21x1_ASAP7_75t_R _27063_ (.A1(_04482_),
    .A2(_04648_),
    .B(net5655),
    .Y(_04649_));
 OAI21x1_ASAP7_75t_R _27064_ (.A1(_04647_),
    .A2(_04649_),
    .B(net6100),
    .Y(_04650_));
 NOR2x1_ASAP7_75t_R _27065_ (.A(net5663),
    .B(net5379),
    .Y(_04651_));
 OAI21x1_ASAP7_75t_R _27066_ (.A1(_04651_),
    .A2(_04541_),
    .B(net6105),
    .Y(_04652_));
 NAND2x1_ASAP7_75t_R _27067_ (.A(net5101),
    .B(net5383),
    .Y(_04653_));
 AO21x1_ASAP7_75t_R _27068_ (.A1(_04653_),
    .A2(_04447_),
    .B(net6103),
    .Y(_04654_));
 AOI21x1_ASAP7_75t_R _27069_ (.A1(_04652_),
    .A2(_04654_),
    .B(net5649),
    .Y(_04655_));
 NOR2x1_ASAP7_75t_R _27070_ (.A(_04650_),
    .B(_04655_),
    .Y(_04656_));
 OAI21x1_ASAP7_75t_R _27071_ (.A1(_04646_),
    .A2(_04656_),
    .B(net5644),
    .Y(_04657_));
 AO21x1_ASAP7_75t_R _27072_ (.A1(_04553_),
    .A2(_04554_),
    .B(_01310_),
    .Y(_04658_));
 AO21x1_ASAP7_75t_R _27073_ (.A1(_04658_),
    .A2(net4549),
    .B(net6098),
    .Y(_04659_));
 NAND2x1_ASAP7_75t_R _27074_ (.A(_04608_),
    .B(_04659_),
    .Y(_04660_));
 OAI21x1_ASAP7_75t_R _27075_ (.A1(net6105),
    .A2(net4636),
    .B(net5646),
    .Y(_04661_));
 INVx1_ASAP7_75t_R _27076_ (.A(_04661_),
    .Y(_04662_));
 NOR2x1_ASAP7_75t_R _27077_ (.A(net5666),
    .B(net5104),
    .Y(_04663_));
 INVx1_ASAP7_75t_R _27078_ (.A(_01319_),
    .Y(_04664_));
 NOR2x1_ASAP7_75t_R _27079_ (.A(_04664_),
    .B(net6094),
    .Y(_04665_));
 AOI21x1_ASAP7_75t_R _27080_ (.A1(net6094),
    .A2(_04663_),
    .B(_04665_),
    .Y(_04666_));
 AOI21x1_ASAP7_75t_R _27081_ (.A1(_04662_),
    .A2(_04666_),
    .B(net5658),
    .Y(_04667_));
 AOI21x1_ASAP7_75t_R _27082_ (.A1(_04660_),
    .A2(_04667_),
    .B(net5644),
    .Y(_04668_));
 OAI21x1_ASAP7_75t_R _27083_ (.A1(net5381),
    .A2(net5662),
    .B(net5036),
    .Y(_04669_));
 INVx1_ASAP7_75t_R _27084_ (.A(_04669_),
    .Y(_04670_));
 NAND2x1_ASAP7_75t_R _27085_ (.A(net6105),
    .B(_04670_),
    .Y(_04671_));
 AOI21x1_ASAP7_75t_R _27086_ (.A1(net5666),
    .A2(net5101),
    .B(net6107),
    .Y(_04672_));
 NAND2x1_ASAP7_75t_R _27087_ (.A(_04501_),
    .B(_04672_),
    .Y(_04673_));
 AOI21x1_ASAP7_75t_R _27089_ (.A1(_04671_),
    .A2(_04673_),
    .B(net5649),
    .Y(_04675_));
 AOI22x1_ASAP7_75t_R _27090_ (.A1(net5380),
    .A2(net5656),
    .B1(net6090),
    .B2(net5645),
    .Y(_04676_));
 OAI21x1_ASAP7_75t_R _27092_ (.A1(_04637_),
    .A2(_04676_),
    .B(net6096),
    .Y(_04678_));
 NAND2x1_ASAP7_75t_R _27093_ (.A(net4731),
    .B(_04552_),
    .Y(_04679_));
 AOI21x1_ASAP7_75t_R _27094_ (.A1(_04678_),
    .A2(_04679_),
    .B(net5660),
    .Y(_04680_));
 OAI21x1_ASAP7_75t_R _27095_ (.A1(_04675_),
    .A2(_04680_),
    .B(net5657),
    .Y(_04681_));
 AOI21x1_ASAP7_75t_R _27096_ (.A1(_04668_),
    .A2(_04681_),
    .B(net6088),
    .Y(_04682_));
 NAND2x1_ASAP7_75t_R _27097_ (.A(_04657_),
    .B(_04682_),
    .Y(_04683_));
 AOI21x1_ASAP7_75t_R _27098_ (.A1(_04542_),
    .A2(net5104),
    .B(net6094),
    .Y(_04684_));
 AND2x2_ASAP7_75t_R _27099_ (.A(net4634),
    .B(_04560_),
    .Y(_04685_));
 OA21x2_ASAP7_75t_R _27100_ (.A1(net5383),
    .A2(net5103),
    .B(net6098),
    .Y(_04686_));
 NAND2x1_ASAP7_75t_R _27101_ (.A(net5649),
    .B(net5657),
    .Y(_04687_));
 AO21x1_ASAP7_75t_R _27102_ (.A1(_04686_),
    .A2(_04477_),
    .B(_04687_),
    .Y(_04688_));
 OAI21x1_ASAP7_75t_R _27103_ (.A1(_04685_),
    .A2(_04688_),
    .B(net6089),
    .Y(_04689_));
 NOR2x1_ASAP7_75t_R _27104_ (.A(net5661),
    .B(net5658),
    .Y(_04690_));
 NAND2x1_ASAP7_75t_R _27105_ (.A(_04459_),
    .B(_04546_),
    .Y(_04691_));
 NAND2x1_ASAP7_75t_R _27106_ (.A(_04690_),
    .B(_04691_),
    .Y(_04692_));
 NOR2x1_ASAP7_75t_R _27107_ (.A(net5663),
    .B(net5102),
    .Y(_04693_));
 INVx1_ASAP7_75t_R _27108_ (.A(_04693_),
    .Y(_04694_));
 NAND2x1_ASAP7_75t_R _27109_ (.A(_04694_),
    .B(_04497_),
    .Y(_04695_));
 INVx1_ASAP7_75t_R _27110_ (.A(_04695_),
    .Y(_04696_));
 INVx1_ASAP7_75t_R _27111_ (.A(_01315_),
    .Y(_04697_));
 NAND2x1_ASAP7_75t_R _27112_ (.A(net6107),
    .B(net6101),
    .Y(_04698_));
 OAI21x1_ASAP7_75t_R _27113_ (.A1(_04641_),
    .A2(_04483_),
    .B(net6099),
    .Y(_04699_));
 OAI21x1_ASAP7_75t_R _27114_ (.A1(_04697_),
    .A2(_04698_),
    .B(_04699_),
    .Y(_04700_));
 OAI22x1_ASAP7_75t_R _27115_ (.A1(_04692_),
    .A2(_04696_),
    .B1(_04700_),
    .B2(net5655),
    .Y(_04701_));
 NOR2x1_ASAP7_75t_R _27116_ (.A(_04689_),
    .B(_04701_),
    .Y(_04702_));
 AO21x1_ASAP7_75t_R _27117_ (.A1(net5380),
    .A2(net5656),
    .B(net4857),
    .Y(_04703_));
 AND3x1_ASAP7_75t_R _27118_ (.A(_04555_),
    .B(_04703_),
    .C(net6096),
    .Y(_04704_));
 AO21x1_ASAP7_75t_R _27119_ (.A1(_04634_),
    .A2(net4460),
    .B(net5660),
    .Y(_04705_));
 AOI21x1_ASAP7_75t_R _27120_ (.A1(net6105),
    .A2(net4731),
    .B(net5647),
    .Y(_04706_));
 NAND2x1_ASAP7_75t_R _27121_ (.A(_04560_),
    .B(_04548_),
    .Y(_04707_));
 AOI21x1_ASAP7_75t_R _27122_ (.A1(_04706_),
    .A2(_04707_),
    .B(net5657),
    .Y(_04708_));
 OAI21x1_ASAP7_75t_R _27123_ (.A1(_04704_),
    .A2(_04705_),
    .B(_04708_),
    .Y(_04709_));
 OAI21x1_ASAP7_75t_R _27124_ (.A1(net6097),
    .A2(net4864),
    .B(net5649),
    .Y(_04710_));
 INVx1_ASAP7_75t_R _27125_ (.A(_04710_),
    .Y(_04711_));
 OAI21x1_ASAP7_75t_R _27126_ (.A1(net5379),
    .A2(net5100),
    .B(net4640),
    .Y(_04712_));
 NOR2x1p5_ASAP7_75t_R _27127_ (.A(net4549),
    .B(net6097),
    .Y(_04713_));
 AOI21x1_ASAP7_75t_R _27128_ (.A1(net6097),
    .A2(_04712_),
    .B(_04713_),
    .Y(_04714_));
 NAND2x1_ASAP7_75t_R _27129_ (.A(_04711_),
    .B(_04714_),
    .Y(_04715_));
 AOI21x1_ASAP7_75t_R _27130_ (.A1(_04477_),
    .A2(_04497_),
    .B(net5649),
    .Y(_04716_));
 AOI21x1_ASAP7_75t_R _27131_ (.A1(_04691_),
    .A2(_04716_),
    .B(net6100),
    .Y(_04717_));
 NAND2x1_ASAP7_75t_R _27132_ (.A(_04715_),
    .B(_04717_),
    .Y(_04718_));
 AOI21x1_ASAP7_75t_R _27134_ (.A1(_04709_),
    .A2(_04718_),
    .B(net6089),
    .Y(_04720_));
 OAI21x1_ASAP7_75t_R _27135_ (.A1(_04702_),
    .A2(_04720_),
    .B(net6088),
    .Y(_04721_));
 NAND2x1_ASAP7_75t_R _27136_ (.A(_04683_),
    .B(_04721_),
    .Y(_00121_));
 AOI21x1_ASAP7_75t_R _27137_ (.A1(net4636),
    .A2(_04653_),
    .B(net6096),
    .Y(_04722_));
 OA21x2_ASAP7_75t_R _27138_ (.A1(net5662),
    .A2(net5381),
    .B(_04539_),
    .Y(_04723_));
 OA21x2_ASAP7_75t_R _27140_ (.A1(_04723_),
    .A2(net4856),
    .B(net6096),
    .Y(_04725_));
 OAI21x1_ASAP7_75t_R _27141_ (.A1(_04722_),
    .A2(_04725_),
    .B(net5648),
    .Y(_04726_));
 AOI21x1_ASAP7_75t_R _27142_ (.A1(net4637),
    .A2(_04585_),
    .B(net6103),
    .Y(_04727_));
 NOR2x1_ASAP7_75t_R _27143_ (.A(net5663),
    .B(net5103),
    .Y(_04728_));
 OA21x2_ASAP7_75t_R _27144_ (.A1(_04728_),
    .A2(_04591_),
    .B(net6103),
    .Y(_04729_));
 OAI21x1_ASAP7_75t_R _27145_ (.A1(net4499),
    .A2(_04729_),
    .B(net5661),
    .Y(_04730_));
 AOI21x1_ASAP7_75t_R _27146_ (.A1(_04726_),
    .A2(_04730_),
    .B(net5657),
    .Y(_04731_));
 INVx1_ASAP7_75t_R _27147_ (.A(net4549),
    .Y(_04732_));
 NOR2x1_ASAP7_75t_R _27148_ (.A(_04732_),
    .B(net4551),
    .Y(_04733_));
 INVx1_ASAP7_75t_R _27149_ (.A(_04627_),
    .Y(_04734_));
 AOI21x1_ASAP7_75t_R _27150_ (.A1(net4633),
    .A2(_04653_),
    .B(net6103),
    .Y(_04735_));
 OAI21x1_ASAP7_75t_R _27151_ (.A1(_04733_),
    .A2(_04735_),
    .B(net5661),
    .Y(_04736_));
 AO21x1_ASAP7_75t_R _27152_ (.A1(net5104),
    .A2(net5663),
    .B(net6092),
    .Y(_04737_));
 AO21x1_ASAP7_75t_R _27153_ (.A1(net5380),
    .A2(net5656),
    .B(net5032),
    .Y(_04738_));
 AOI21x1_ASAP7_75t_R _27154_ (.A1(_04738_),
    .A2(_04497_),
    .B(net5660),
    .Y(_04739_));
 OAI21x1_ASAP7_75t_R _27155_ (.A1(net4856),
    .A2(_04737_),
    .B(_04739_),
    .Y(_04740_));
 AOI21x1_ASAP7_75t_R _27156_ (.A1(_04736_),
    .A2(_04740_),
    .B(net6101),
    .Y(_04741_));
 NOR3x1_ASAP7_75t_R _27157_ (.A(_04731_),
    .B(_04741_),
    .C(net6089),
    .Y(_04742_));
 AOI21x1_ASAP7_75t_R _27158_ (.A1(net5663),
    .A2(net5103),
    .B(net6105),
    .Y(_04743_));
 AOI21x1_ASAP7_75t_R _27159_ (.A1(net5383),
    .A2(net5100),
    .B(net6096),
    .Y(_04744_));
 AOI22x1_ASAP7_75t_R _27160_ (.A1(_04743_),
    .A2(net4460),
    .B1(_04744_),
    .B2(net4854),
    .Y(_04745_));
 AOI21x1_ASAP7_75t_R _27161_ (.A1(net6096),
    .A2(_04547_),
    .B(net5648),
    .Y(_04746_));
 NAND2x1_ASAP7_75t_R _27162_ (.A(_04555_),
    .B(_04634_),
    .Y(_04747_));
 AOI21x1_ASAP7_75t_R _27163_ (.A1(_04746_),
    .A2(_04747_),
    .B(net6100),
    .Y(_04748_));
 OAI21x1_ASAP7_75t_R _27164_ (.A1(net5660),
    .A2(_04745_),
    .B(_04748_),
    .Y(_04749_));
 OAI21x1_ASAP7_75t_R _27165_ (.A1(net6098),
    .A2(_04607_),
    .B(net5661),
    .Y(_04750_));
 NOR2x1_ASAP7_75t_R _27166_ (.A(_04598_),
    .B(_04750_),
    .Y(_04751_));
 OAI21x1_ASAP7_75t_R _27167_ (.A1(_04723_),
    .A2(_04637_),
    .B(net6099),
    .Y(_04752_));
 NAND2x1_ASAP7_75t_R _27168_ (.A(net5666),
    .B(net5102),
    .Y(_04753_));
 NAND2x1_ASAP7_75t_R _27169_ (.A(_04753_),
    .B(_04684_),
    .Y(_04754_));
 AOI21x1_ASAP7_75t_R _27171_ (.A1(_04752_),
    .A2(_04754_),
    .B(net5661),
    .Y(_04756_));
 OAI21x1_ASAP7_75t_R _27172_ (.A1(_04751_),
    .A2(_04756_),
    .B(net6101),
    .Y(_04757_));
 NAND2x1_ASAP7_75t_R _27173_ (.A(_04749_),
    .B(_04757_),
    .Y(_04758_));
 OAI21x1_ASAP7_75t_R _27174_ (.A1(net5644),
    .A2(_04758_),
    .B(net6088),
    .Y(_04759_));
 OA21x2_ASAP7_75t_R _27175_ (.A1(_01320_),
    .A2(net6102),
    .B(net5646),
    .Y(_04760_));
 NAND2x1_ASAP7_75t_R _27176_ (.A(_04760_),
    .B(_04754_),
    .Y(_04761_));
 NOR2x1_ASAP7_75t_R _27177_ (.A(net5035),
    .B(_04434_),
    .Y(_04762_));
 NAND2x1_ASAP7_75t_R _27178_ (.A(_01317_),
    .B(net6102),
    .Y(_04763_));
 OA21x2_ASAP7_75t_R _27179_ (.A1(_04762_),
    .A2(net6102),
    .B(_04763_),
    .Y(_04764_));
 AOI21x1_ASAP7_75t_R _27180_ (.A1(net5659),
    .A2(_04764_),
    .B(net5658),
    .Y(_04765_));
 NAND2x1_ASAP7_75t_R _27181_ (.A(_04761_),
    .B(_04765_),
    .Y(_04766_));
 OAI21x1_ASAP7_75t_R _27182_ (.A1(net4501),
    .A2(net4550),
    .B(net6103),
    .Y(_04767_));
 OA21x2_ASAP7_75t_R _27183_ (.A1(net6104),
    .A2(net4864),
    .B(net5661),
    .Y(_04768_));
 AOI21x1_ASAP7_75t_R _27184_ (.A1(_04767_),
    .A2(_04768_),
    .B(net6101),
    .Y(_04769_));
 NOR2x1_ASAP7_75t_R _27185_ (.A(_04512_),
    .B(net5101),
    .Y(_04770_));
 AND2x2_ASAP7_75t_R _27186_ (.A(_01302_),
    .B(_01308_),
    .Y(_04771_));
 NOR2x1_ASAP7_75t_R _27187_ (.A(_04771_),
    .B(net5103),
    .Y(_04772_));
 OAI21x1_ASAP7_75t_R _27188_ (.A1(_04770_),
    .A2(net4632),
    .B(net6107),
    .Y(_04773_));
 NAND3x1_ASAP7_75t_R _27189_ (.A(_04773_),
    .B(_04699_),
    .C(net5650),
    .Y(_04774_));
 AOI21x1_ASAP7_75t_R _27190_ (.A1(_04769_),
    .A2(_04774_),
    .B(net5644),
    .Y(_04775_));
 NAND2x1_ASAP7_75t_R _27191_ (.A(_04766_),
    .B(_04775_),
    .Y(_04776_));
 AO21x1_ASAP7_75t_R _27192_ (.A1(net4548),
    .A2(net4855),
    .B(net6093),
    .Y(_04777_));
 OA21x2_ASAP7_75t_R _27193_ (.A1(_01318_),
    .A2(net6107),
    .B(net5661),
    .Y(_04778_));
 AOI21x1_ASAP7_75t_R _27194_ (.A1(_04777_),
    .A2(_04778_),
    .B(net6101),
    .Y(_04779_));
 NAND2x1_ASAP7_75t_R _27195_ (.A(_04459_),
    .B(_04601_),
    .Y(_04780_));
 AOI21x1_ASAP7_75t_R _27196_ (.A1(net4548),
    .A2(_04672_),
    .B(net5661),
    .Y(_04781_));
 NAND2x1_ASAP7_75t_R _27197_ (.A(_04780_),
    .B(_04781_),
    .Y(_04782_));
 AOI21x1_ASAP7_75t_R _27198_ (.A1(_04779_),
    .A2(_04782_),
    .B(net6089),
    .Y(_04783_));
 NAND2x1_ASAP7_75t_R _27199_ (.A(_01315_),
    .B(net6091),
    .Y(_04784_));
 AOI21x1_ASAP7_75t_R _27200_ (.A1(net5666),
    .A2(net5102),
    .B(net6091),
    .Y(_04785_));
 AOI21x1_ASAP7_75t_R _27201_ (.A1(_04501_),
    .A2(_04785_),
    .B(net5654),
    .Y(_04786_));
 AOI21x1_ASAP7_75t_R _27202_ (.A1(_04784_),
    .A2(_04786_),
    .B(net5658),
    .Y(_04787_));
 NAND2x1p5_ASAP7_75t_R _27203_ (.A(net6106),
    .B(net4549),
    .Y(_04788_));
 NOR2x1_ASAP7_75t_R _27204_ (.A(_04522_),
    .B(_04788_),
    .Y(_04789_));
 AND2x2_ASAP7_75t_R _27205_ (.A(_04672_),
    .B(_04521_),
    .Y(_04790_));
 OAI21x1_ASAP7_75t_R _27206_ (.A1(_04789_),
    .A2(_04790_),
    .B(net5652),
    .Y(_04791_));
 NAND2x1_ASAP7_75t_R _27207_ (.A(_04787_),
    .B(_04791_),
    .Y(_04792_));
 AOI21x1_ASAP7_75t_R _27208_ (.A1(_04783_),
    .A2(_04792_),
    .B(net6088),
    .Y(_04793_));
 NAND2x1_ASAP7_75t_R _27209_ (.A(_04776_),
    .B(_04793_),
    .Y(_04794_));
 OAI21x1_ASAP7_75t_R _27210_ (.A1(_04742_),
    .A2(_04759_),
    .B(_04794_),
    .Y(_00122_));
 AO21x1_ASAP7_75t_R _27211_ (.A1(net5103),
    .A2(net5037),
    .B(net6102),
    .Y(_04795_));
 AOI21x1_ASAP7_75t_R _27212_ (.A1(net6102),
    .A2(net4856),
    .B(net6101),
    .Y(_04796_));
 OAI21x1_ASAP7_75t_R _27213_ (.A1(_04541_),
    .A2(_04795_),
    .B(_04796_),
    .Y(_04797_));
 OAI21x1_ASAP7_75t_R _27214_ (.A1(_04723_),
    .A2(_04772_),
    .B(net6105),
    .Y(_04798_));
 AOI21x1_ASAP7_75t_R _27215_ (.A1(net4731),
    .A2(_04548_),
    .B(net5658),
    .Y(_04799_));
 NAND2x1_ASAP7_75t_R _27216_ (.A(_04798_),
    .B(_04799_),
    .Y(_04800_));
 AOI21x1_ASAP7_75t_R _27217_ (.A1(_04797_),
    .A2(_04800_),
    .B(net5655),
    .Y(_04801_));
 OAI21x1_ASAP7_75t_R _27218_ (.A1(_04447_),
    .A2(_04698_),
    .B(_04623_),
    .Y(_04802_));
 NAND2x1_ASAP7_75t_R _27219_ (.A(net6101),
    .B(_04753_),
    .Y(_04803_));
 INVx1_ASAP7_75t_R _27220_ (.A(net5038),
    .Y(_04804_));
 AO21x1_ASAP7_75t_R _27221_ (.A1(net5104),
    .A2(_04804_),
    .B(net6102),
    .Y(_04805_));
 INVx1_ASAP7_75t_R _27222_ (.A(_04460_),
    .Y(_04806_));
 NAND2x1_ASAP7_75t_R _27223_ (.A(net6091),
    .B(_04806_),
    .Y(_04807_));
 OAI22x1_ASAP7_75t_R _27224_ (.A1(_04803_),
    .A2(_04805_),
    .B1(_04807_),
    .B2(net6101),
    .Y(_04808_));
 OAI21x1_ASAP7_75t_R _27225_ (.A1(_04802_),
    .A2(_04808_),
    .B(net6089),
    .Y(_04809_));
 NOR2x1_ASAP7_75t_R _27226_ (.A(_04801_),
    .B(_04809_),
    .Y(_04810_));
 OAI21x1_ASAP7_75t_R _27227_ (.A1(net4852),
    .A2(_04772_),
    .B(net6107),
    .Y(_04811_));
 AOI21x1_ASAP7_75t_R _27228_ (.A1(_04699_),
    .A2(_04811_),
    .B(net5650),
    .Y(_04812_));
 OAI21x1_ASAP7_75t_R _27229_ (.A1(_04739_),
    .A2(_04812_),
    .B(net6101),
    .Y(_04813_));
 OAI21x1_ASAP7_75t_R _27230_ (.A1(net4550),
    .A2(_04723_),
    .B(net6095),
    .Y(_04814_));
 OAI21x1_ASAP7_75t_R _27231_ (.A1(net4856),
    .A2(_04676_),
    .B(net6105),
    .Y(_04815_));
 AOI21x1_ASAP7_75t_R _27232_ (.A1(_04814_),
    .A2(_04815_),
    .B(net5660),
    .Y(_04816_));
 AOI21x1_ASAP7_75t_R _27233_ (.A1(_04613_),
    .A2(_04673_),
    .B(net5655),
    .Y(_04817_));
 OAI21x1_ASAP7_75t_R _27234_ (.A1(_04816_),
    .A2(_04817_),
    .B(net5658),
    .Y(_04818_));
 AOI21x1_ASAP7_75t_R _27235_ (.A1(_04813_),
    .A2(_04818_),
    .B(net6089),
    .Y(_04819_));
 OAI21x1_ASAP7_75t_R _27236_ (.A1(_04810_),
    .A2(_04819_),
    .B(net6088),
    .Y(_04820_));
 OAI21x1_ASAP7_75t_R _27237_ (.A1(_04611_),
    .A2(_04505_),
    .B(net6091),
    .Y(_04821_));
 OAI21x1_ASAP7_75t_R _27238_ (.A1(net4547),
    .A2(_04737_),
    .B(_04821_),
    .Y(_04822_));
 OAI21x1_ASAP7_75t_R _27239_ (.A1(_04693_),
    .A2(_04504_),
    .B(net6091),
    .Y(_04823_));
 AOI21x1_ASAP7_75t_R _27240_ (.A1(_04458_),
    .A2(_04823_),
    .B(net5658),
    .Y(_04824_));
 OAI21x1_ASAP7_75t_R _27241_ (.A1(net5655),
    .A2(_04822_),
    .B(_04824_),
    .Y(_04825_));
 NOR2x1_ASAP7_75t_R _27242_ (.A(_04522_),
    .B(_04648_),
    .Y(_04826_));
 AND3x1_ASAP7_75t_R _27243_ (.A(net4864),
    .B(_04447_),
    .C(net6104),
    .Y(_04827_));
 OAI21x1_ASAP7_75t_R _27244_ (.A1(_04826_),
    .A2(_04827_),
    .B(net5650),
    .Y(_04828_));
 AO21x1_ASAP7_75t_R _27245_ (.A1(_04658_),
    .A2(net4636),
    .B(net6095),
    .Y(_04829_));
 AOI21x1_ASAP7_75t_R _27246_ (.A1(_04516_),
    .A2(_04743_),
    .B(net5649),
    .Y(_04830_));
 AOI21x1_ASAP7_75t_R _27247_ (.A1(_04829_),
    .A2(_04830_),
    .B(net6100),
    .Y(_04831_));
 NAND2x1_ASAP7_75t_R _27248_ (.A(_04828_),
    .B(_04831_),
    .Y(_04832_));
 AOI21x1_ASAP7_75t_R _27249_ (.A1(_04825_),
    .A2(_04832_),
    .B(_04536_),
    .Y(_04833_));
 AO21x1_ASAP7_75t_R _27250_ (.A1(net4850),
    .A2(net4549),
    .B(net6105),
    .Y(_04834_));
 OAI21x1_ASAP7_75t_R _27251_ (.A1(_04670_),
    .A2(_04522_),
    .B(net6105),
    .Y(_04835_));
 AOI21x1_ASAP7_75t_R _27252_ (.A1(_04834_),
    .A2(_04835_),
    .B(net5646),
    .Y(_04836_));
 OAI21x1_ASAP7_75t_R _27253_ (.A1(_04806_),
    .A2(net4862),
    .B(net6094),
    .Y(_04837_));
 NOR2x1_ASAP7_75t_R _27254_ (.A(net5663),
    .B(net5383),
    .Y(_04838_));
 OAI21x1_ASAP7_75t_R _27255_ (.A1(_04611_),
    .A2(_04838_),
    .B(net6102),
    .Y(_04839_));
 AOI21x1_ASAP7_75t_R _27256_ (.A1(_04837_),
    .A2(_04839_),
    .B(net5659),
    .Y(_04840_));
 OAI21x1_ASAP7_75t_R _27257_ (.A1(_04836_),
    .A2(_04840_),
    .B(net5658),
    .Y(_04841_));
 INVx1_ASAP7_75t_R _27258_ (.A(net4634),
    .Y(_04842_));
 AOI21x1_ASAP7_75t_R _27259_ (.A1(_04842_),
    .A2(_04821_),
    .B(net5655),
    .Y(_04843_));
 OAI21x1_ASAP7_75t_R _27260_ (.A1(net4851),
    .A2(_04806_),
    .B(net6094),
    .Y(_04844_));
 NAND2x1_ASAP7_75t_R _27261_ (.A(_04556_),
    .B(_04643_),
    .Y(_04845_));
 AOI21x1_ASAP7_75t_R _27262_ (.A1(_04844_),
    .A2(_04845_),
    .B(net5660),
    .Y(_04846_));
 OAI21x1_ASAP7_75t_R _27263_ (.A1(_04843_),
    .A2(_04846_),
    .B(net6101),
    .Y(_04847_));
 AOI21x1_ASAP7_75t_R _27264_ (.A1(_04841_),
    .A2(_04847_),
    .B(net6089),
    .Y(_04848_));
 INVx1_ASAP7_75t_R _27265_ (.A(_04578_),
    .Y(_04849_));
 OAI21x1_ASAP7_75t_R _27266_ (.A1(_04833_),
    .A2(_04848_),
    .B(net5643),
    .Y(_04850_));
 NAND2x1_ASAP7_75t_R _27267_ (.A(_04820_),
    .B(_04850_),
    .Y(_00123_));
 NAND2x1_ASAP7_75t_R _27268_ (.A(net5103),
    .B(net6107),
    .Y(_04851_));
 AND2x2_ASAP7_75t_R _27269_ (.A(_04851_),
    .B(net5661),
    .Y(_04852_));
 NAND2x1_ASAP7_75t_R _27270_ (.A(_04540_),
    .B(_04497_),
    .Y(_04853_));
 AO21x1_ASAP7_75t_R _27271_ (.A1(_04852_),
    .A2(_04853_),
    .B(net6089),
    .Y(_04854_));
 AO21x1_ASAP7_75t_R _27272_ (.A1(_04482_),
    .A2(net6092),
    .B(net5661),
    .Y(_04855_));
 NAND2x1_ASAP7_75t_R _27273_ (.A(_04564_),
    .B(_04691_),
    .Y(_04856_));
 NOR2x1_ASAP7_75t_R _27274_ (.A(_04855_),
    .B(_04856_),
    .Y(_04857_));
 OAI21x1_ASAP7_75t_R _27275_ (.A1(_04854_),
    .A2(_04857_),
    .B(net6088),
    .Y(_04858_));
 NOR2x1_ASAP7_75t_R _27276_ (.A(net5653),
    .B(_04506_),
    .Y(_04859_));
 AO21x1_ASAP7_75t_R _27277_ (.A1(net5103),
    .A2(net5037),
    .B(net6094),
    .Y(_04860_));
 NOR2x1_ASAP7_75t_R _27278_ (.A(_04504_),
    .B(_04860_),
    .Y(_04861_));
 NAND2x1_ASAP7_75t_R _27279_ (.A(net5666),
    .B(net5378),
    .Y(_04862_));
 NAND2x1_ASAP7_75t_R _27280_ (.A(_04459_),
    .B(_04862_),
    .Y(_04863_));
 OAI21x1_ASAP7_75t_R _27281_ (.A1(net6106),
    .A2(_04863_),
    .B(net5653),
    .Y(_04864_));
 OAI21x1_ASAP7_75t_R _27282_ (.A1(_04861_),
    .A2(_04864_),
    .B(net6089),
    .Y(_04865_));
 AOI21x1_ASAP7_75t_R _27283_ (.A1(net4500),
    .A2(_04859_),
    .B(_04865_),
    .Y(_04866_));
 OAI21x1_ASAP7_75t_R _27284_ (.A1(_04858_),
    .A2(_04866_),
    .B(net6101),
    .Y(_04867_));
 AO21x1_ASAP7_75t_R _27285_ (.A1(net5102),
    .A2(net4861),
    .B(net6091),
    .Y(_04868_));
 OA21x2_ASAP7_75t_R _27286_ (.A1(_04563_),
    .A2(_04868_),
    .B(_04752_),
    .Y(_04869_));
 AO21x1_ASAP7_75t_R _27287_ (.A1(_04694_),
    .A2(net4864),
    .B(net6093),
    .Y(_04870_));
 AO21x1_ASAP7_75t_R _27288_ (.A1(_04870_),
    .A2(_04608_),
    .B(net5644),
    .Y(_04871_));
 AOI21x1_ASAP7_75t_R _27289_ (.A1(net5655),
    .A2(_04869_),
    .B(_04871_),
    .Y(_04872_));
 NAND2x1_ASAP7_75t_R _27290_ (.A(_04501_),
    .B(_04785_),
    .Y(_04873_));
 AOI21x1_ASAP7_75t_R _27291_ (.A1(_04873_),
    .A2(_04695_),
    .B(net5653),
    .Y(_04874_));
 INVx1_ASAP7_75t_R _27292_ (.A(_04521_),
    .Y(_04875_));
 OAI21x1_ASAP7_75t_R _27293_ (.A1(_04728_),
    .A2(_04875_),
    .B(net6106),
    .Y(_04876_));
 AO21x1_ASAP7_75t_R _27294_ (.A1(_04862_),
    .A2(_04459_),
    .B(net6106),
    .Y(_04877_));
 AOI21x1_ASAP7_75t_R _27295_ (.A1(_04876_),
    .A2(_04877_),
    .B(net5661),
    .Y(_04878_));
 OAI21x1_ASAP7_75t_R _27296_ (.A1(_04874_),
    .A2(_04878_),
    .B(net5644),
    .Y(_04879_));
 NAND2x1_ASAP7_75t_R _27297_ (.A(net5643),
    .B(_04879_),
    .Y(_04880_));
 NOR2x1_ASAP7_75t_R _27298_ (.A(_04872_),
    .B(_04880_),
    .Y(_04881_));
 AO21x1_ASAP7_75t_R _27299_ (.A1(net5100),
    .A2(net5034),
    .B(net6105),
    .Y(_04882_));
 NOR2x1_ASAP7_75t_R _27300_ (.A(_04732_),
    .B(_04882_),
    .Y(_04883_));
 AOI21x1_ASAP7_75t_R _27301_ (.A1(net6096),
    .A2(_04703_),
    .B(net5660),
    .Y(_04884_));
 AOI21x1_ASAP7_75t_R _27302_ (.A1(_04635_),
    .A2(_04884_),
    .B(net6089),
    .Y(_04885_));
 OAI21x1_ASAP7_75t_R _27303_ (.A1(_04583_),
    .A2(_04883_),
    .B(_04885_),
    .Y(_04886_));
 OA21x2_ASAP7_75t_R _27304_ (.A1(_04512_),
    .A2(net6107),
    .B(net5661),
    .Y(_04887_));
 AOI21x1_ASAP7_75t_R _27305_ (.A1(_04788_),
    .A2(_04887_),
    .B(net5644),
    .Y(_04888_));
 OA21x2_ASAP7_75t_R _27306_ (.A1(net6107),
    .A2(net4855),
    .B(net5649),
    .Y(_04889_));
 AO21x1_ASAP7_75t_R _27307_ (.A1(_04753_),
    .A2(_04734_),
    .B(net6098),
    .Y(_04890_));
 NAND2x1_ASAP7_75t_R _27308_ (.A(_04889_),
    .B(_04890_),
    .Y(_04891_));
 AOI21x1_ASAP7_75t_R _27309_ (.A1(_04888_),
    .A2(_04891_),
    .B(_04849_),
    .Y(_04892_));
 AOI21x1_ASAP7_75t_R _27310_ (.A1(_04886_),
    .A2(_04892_),
    .B(net6100),
    .Y(_04893_));
 OA21x2_ASAP7_75t_R _27311_ (.A1(_04585_),
    .A2(net6097),
    .B(net5649),
    .Y(_04894_));
 NOR2x1_ASAP7_75t_R _27312_ (.A(_04727_),
    .B(_04713_),
    .Y(_04895_));
 NAND2x1_ASAP7_75t_R _27313_ (.A(_04895_),
    .B(_04894_),
    .Y(_04896_));
 AO21x1_ASAP7_75t_R _27314_ (.A1(_04658_),
    .A2(net4549),
    .B(net6107),
    .Y(_04897_));
 AND2x2_ASAP7_75t_R _27315_ (.A(_04628_),
    .B(net5659),
    .Y(_04898_));
 AOI21x1_ASAP7_75t_R _27316_ (.A1(_04897_),
    .A2(_04898_),
    .B(net5644),
    .Y(_04899_));
 NAND2x1_ASAP7_75t_R _27317_ (.A(_04899_),
    .B(_04896_),
    .Y(_04900_));
 AND2x2_ASAP7_75t_R _27318_ (.A(net5655),
    .B(_04566_),
    .Y(_04901_));
 AOI21x1_ASAP7_75t_R _27319_ (.A1(_04860_),
    .A2(_04901_),
    .B(net6089),
    .Y(_04902_));
 NAND2x1_ASAP7_75t_R _27320_ (.A(_04694_),
    .B(_04601_),
    .Y(_04903_));
 AOI21x1_ASAP7_75t_R _27321_ (.A1(_04477_),
    .A2(_04686_),
    .B(net5649),
    .Y(_04904_));
 NAND2x1_ASAP7_75t_R _27322_ (.A(_04903_),
    .B(_04904_),
    .Y(_04905_));
 AOI21x1_ASAP7_75t_R _27323_ (.A1(_04902_),
    .A2(_04905_),
    .B(net6088),
    .Y(_04906_));
 NAND2x1_ASAP7_75t_R _27324_ (.A(_04906_),
    .B(_04900_),
    .Y(_04907_));
 NAND2x1_ASAP7_75t_R _27325_ (.A(_04907_),
    .B(_04893_),
    .Y(_04908_));
 OAI21x1_ASAP7_75t_R _27326_ (.A1(_04867_),
    .A2(_04881_),
    .B(_04908_),
    .Y(_00124_));
 OA21x2_ASAP7_75t_R _27327_ (.A1(_04637_),
    .A2(_04723_),
    .B(net6105),
    .Y(_04909_));
 OAI21x1_ASAP7_75t_R _27328_ (.A1(_04909_),
    .A2(_04568_),
    .B(net5657),
    .Y(_04910_));
 NAND2x1_ASAP7_75t_R _27329_ (.A(net4855),
    .B(_04734_),
    .Y(_04911_));
 INVx1_ASAP7_75t_R _27330_ (.A(_04771_),
    .Y(_04912_));
 OA21x2_ASAP7_75t_R _27331_ (.A1(net5101),
    .A2(_04589_),
    .B(net6104),
    .Y(_04913_));
 AOI221x1_ASAP7_75t_R _27332_ (.A1(net6095),
    .A2(_04911_),
    .B1(net4631),
    .B2(_04913_),
    .C(net5660),
    .Y(_04914_));
 NOR2x1_ASAP7_75t_R _27333_ (.A(_04670_),
    .B(net5660),
    .Y(_04915_));
 AOI21x1_ASAP7_75t_R _27334_ (.A1(_04915_),
    .A2(_04882_),
    .B(net5657),
    .Y(_04916_));
 OA21x2_ASAP7_75t_R _27335_ (.A1(_04806_),
    .A2(net6102),
    .B(net5661),
    .Y(_04917_));
 NAND2x1_ASAP7_75t_R _27336_ (.A(_04815_),
    .B(_04917_),
    .Y(_04918_));
 AOI21x1_ASAP7_75t_R _27337_ (.A1(_04916_),
    .A2(_04918_),
    .B(net6088),
    .Y(_04919_));
 OAI21x1_ASAP7_75t_R _27338_ (.A1(_04910_),
    .A2(_04914_),
    .B(_04919_),
    .Y(_04920_));
 NAND2x1_ASAP7_75t_R _27339_ (.A(net4731),
    .B(net4634),
    .Y(_04921_));
 OAI21x1_ASAP7_75t_R _27340_ (.A1(net4851),
    .A2(_04728_),
    .B(net6093),
    .Y(_04922_));
 AND3x1_ASAP7_75t_R _27341_ (.A(_04921_),
    .B(net5655),
    .C(_04922_),
    .Y(_04923_));
 NOR2x1_ASAP7_75t_R _27342_ (.A(net5378),
    .B(net6093),
    .Y(_04924_));
 AOI21x1_ASAP7_75t_R _27343_ (.A1(_04501_),
    .A2(_04497_),
    .B(_04924_),
    .Y(_04925_));
 AO21x1_ASAP7_75t_R _27344_ (.A1(_04925_),
    .A2(net5661),
    .B(net6101),
    .Y(_04926_));
 AOI21x1_ASAP7_75t_R _27345_ (.A1(net6104),
    .A2(net4863),
    .B(net5661),
    .Y(_04927_));
 OAI21x1_ASAP7_75t_R _27346_ (.A1(net4635),
    .A2(_04723_),
    .B(net6095),
    .Y(_04928_));
 AOI21x1_ASAP7_75t_R _27347_ (.A1(_04927_),
    .A2(_04928_),
    .B(net5657),
    .Y(_04929_));
 AO21x1_ASAP7_75t_R _27348_ (.A1(_04653_),
    .A2(net4636),
    .B(net6103),
    .Y(_04930_));
 NAND2x1_ASAP7_75t_R _27349_ (.A(_04582_),
    .B(_04930_),
    .Y(_04931_));
 AOI21x1_ASAP7_75t_R _27350_ (.A1(_04929_),
    .A2(_04931_),
    .B(_04849_),
    .Y(_04932_));
 OAI21x1_ASAP7_75t_R _27351_ (.A1(_04923_),
    .A2(_04926_),
    .B(_04932_),
    .Y(_04933_));
 AOI21x1_ASAP7_75t_R _27352_ (.A1(_04920_),
    .A2(_04933_),
    .B(net6089),
    .Y(_04934_));
 NOR2x1_ASAP7_75t_R _27353_ (.A(_04804_),
    .B(net6095),
    .Y(_04935_));
 AOI21x1_ASAP7_75t_R _27354_ (.A1(net6095),
    .A2(_04560_),
    .B(_04935_),
    .Y(_04936_));
 OAI21x1_ASAP7_75t_R _27355_ (.A1(net5649),
    .A2(_04936_),
    .B(net6100),
    .Y(_04937_));
 NAND2x1_ASAP7_75t_R _27356_ (.A(_04600_),
    .B(_04479_),
    .Y(_04938_));
 AO21x1_ASAP7_75t_R _27357_ (.A1(_04738_),
    .A2(net4731),
    .B(net6105),
    .Y(_04939_));
 AOI21x1_ASAP7_75t_R _27358_ (.A1(_04938_),
    .A2(_04939_),
    .B(net5660),
    .Y(_04940_));
 NOR2x1_ASAP7_75t_R _27359_ (.A(_04937_),
    .B(_04940_),
    .Y(_04941_));
 NOR2x1_ASAP7_75t_R _27360_ (.A(_04643_),
    .B(_04661_),
    .Y(_04942_));
 AOI21x1_ASAP7_75t_R _27361_ (.A1(_04669_),
    .A2(net4850),
    .B(net6105),
    .Y(_04943_));
 AOI21x1_ASAP7_75t_R _27362_ (.A1(_04554_),
    .A2(_04553_),
    .B(_04912_),
    .Y(_04944_));
 OAI21x1_ASAP7_75t_R _27363_ (.A1(net6099),
    .A2(_04944_),
    .B(net5659),
    .Y(_04945_));
 NOR2x1_ASAP7_75t_R _27364_ (.A(_04943_),
    .B(_04945_),
    .Y(_04946_));
 OAI21x1_ASAP7_75t_R _27365_ (.A1(_04942_),
    .A2(_04946_),
    .B(net5657),
    .Y(_04947_));
 NAND2x1_ASAP7_75t_R _27366_ (.A(net6088),
    .B(_04947_),
    .Y(_04948_));
 OAI21x1_ASAP7_75t_R _27367_ (.A1(_04941_),
    .A2(_04948_),
    .B(net6089),
    .Y(_04949_));
 INVx2_ASAP7_75t_R _27368_ (.A(_04713_),
    .Y(_04950_));
 AO21x1_ASAP7_75t_R _27369_ (.A1(net4858),
    .A2(_04610_),
    .B(net6105),
    .Y(_04951_));
 AOI21x1_ASAP7_75t_R _27370_ (.A1(_04950_),
    .A2(_04951_),
    .B(net5660),
    .Y(_04952_));
 OA21x2_ASAP7_75t_R _27371_ (.A1(_04723_),
    .A2(net6105),
    .B(net5660),
    .Y(_04953_));
 NAND2x1_ASAP7_75t_R _27372_ (.A(_04521_),
    .B(_04479_),
    .Y(_04954_));
 AO21x1_ASAP7_75t_R _27373_ (.A1(_04953_),
    .A2(_04954_),
    .B(net5657),
    .Y(_04955_));
 NOR2x1_ASAP7_75t_R _27374_ (.A(_04955_),
    .B(_04952_),
    .Y(_04956_));
 AO21x1_ASAP7_75t_R _27375_ (.A1(net5101),
    .A2(net5033),
    .B(net6094),
    .Y(_04957_));
 OAI21x1_ASAP7_75t_R _27376_ (.A1(net4863),
    .A2(_04957_),
    .B(net5650),
    .Y(_04958_));
 OA21x2_ASAP7_75t_R _27377_ (.A1(net5663),
    .A2(net5379),
    .B(_04548_),
    .Y(_04959_));
 NOR2x1_ASAP7_75t_R _27378_ (.A(_04958_),
    .B(_04959_),
    .Y(_04960_));
 AO21x1_ASAP7_75t_R _27379_ (.A1(net5663),
    .A2(net6104),
    .B(net5650),
    .Y(_04961_));
 OA21x2_ASAP7_75t_R _27380_ (.A1(_04651_),
    .A2(_04663_),
    .B(net6099),
    .Y(_04962_));
 OAI21x1_ASAP7_75t_R _27381_ (.A1(_04961_),
    .A2(_04962_),
    .B(net5658),
    .Y(_04963_));
 OAI21x1_ASAP7_75t_R _27382_ (.A1(_04960_),
    .A2(_04963_),
    .B(_04849_),
    .Y(_04964_));
 NOR2x1_ASAP7_75t_R _27383_ (.A(_04964_),
    .B(_04956_),
    .Y(_04965_));
 NOR2x1_ASAP7_75t_R _27384_ (.A(_04949_),
    .B(_04965_),
    .Y(_04966_));
 NOR2x1_ASAP7_75t_R _27385_ (.A(_04934_),
    .B(_04966_),
    .Y(_00125_));
 INVx1_ASAP7_75t_R _27386_ (.A(_04805_),
    .Y(_04967_));
 NOR2x1_ASAP7_75t_R _27387_ (.A(_04663_),
    .B(_04860_),
    .Y(_04968_));
 OAI21x1_ASAP7_75t_R _27388_ (.A1(_04967_),
    .A2(_04968_),
    .B(net5651),
    .Y(_04969_));
 AOI21x1_ASAP7_75t_R _27389_ (.A1(net4440),
    .A2(_04969_),
    .B(net5658),
    .Y(_04970_));
 NAND2x1_ASAP7_75t_R _27390_ (.A(net5103),
    .B(net5383),
    .Y(_04971_));
 NOR2x1_ASAP7_75t_R _27391_ (.A(net6104),
    .B(_04971_),
    .Y(_04972_));
 AOI211x1_ASAP7_75t_R _27392_ (.A1(net4459),
    .A2(_04643_),
    .B(_04972_),
    .C(net5661),
    .Y(_04973_));
 AOI21x1_ASAP7_75t_R _27393_ (.A1(_01313_),
    .A2(net6107),
    .B(net5654),
    .Y(_04974_));
 AO21x1_ASAP7_75t_R _27394_ (.A1(_04922_),
    .A2(_04974_),
    .B(net6101),
    .Y(_04975_));
 OAI21x1_ASAP7_75t_R _27395_ (.A1(_04973_),
    .A2(_04975_),
    .B(net6089),
    .Y(_04976_));
 OAI21x1_ASAP7_75t_R _27396_ (.A1(_04970_),
    .A2(_04976_),
    .B(net6088),
    .Y(_04977_));
 INVx1_ASAP7_75t_R _27397_ (.A(_04815_),
    .Y(_04978_));
 AO21x1_ASAP7_75t_R _27398_ (.A1(net4550),
    .A2(net6095),
    .B(net5657),
    .Y(_04979_));
 OAI21x1_ASAP7_75t_R _27399_ (.A1(_04978_),
    .A2(_04979_),
    .B(net5660),
    .Y(_04980_));
 NAND3x1_ASAP7_75t_R _27400_ (.A(net4858),
    .B(net6095),
    .C(net4849),
    .Y(_04981_));
 AO21x1_ASAP7_75t_R _27401_ (.A1(_04653_),
    .A2(_04862_),
    .B(net6099),
    .Y(_04982_));
 AOI21x1_ASAP7_75t_R _27402_ (.A1(_04981_),
    .A2(_04982_),
    .B(net6100),
    .Y(_04983_));
 OAI21x1_ASAP7_75t_R _27403_ (.A1(_04980_),
    .A2(_04983_),
    .B(net5644),
    .Y(_04984_));
 NOR2x1_ASAP7_75t_R _27404_ (.A(_04541_),
    .B(_04543_),
    .Y(_04985_));
 OAI21x1_ASAP7_75t_R _27405_ (.A1(_04665_),
    .A2(_04985_),
    .B(net6101),
    .Y(_04986_));
 INVx1_ASAP7_75t_R _27406_ (.A(_04676_),
    .Y(_04987_));
 AOI21x1_ASAP7_75t_R _27407_ (.A1(_04658_),
    .A2(_04987_),
    .B(net6105),
    .Y(_04988_));
 OA21x2_ASAP7_75t_R _27408_ (.A1(_04504_),
    .A2(_04838_),
    .B(net6102),
    .Y(_04989_));
 OAI21x1_ASAP7_75t_R _27409_ (.A1(_04988_),
    .A2(_04989_),
    .B(net5658),
    .Y(_04990_));
 AOI21x1_ASAP7_75t_R _27410_ (.A1(_04986_),
    .A2(_04990_),
    .B(net5659),
    .Y(_04991_));
 NOR2x1_ASAP7_75t_R _27411_ (.A(_04984_),
    .B(_04991_),
    .Y(_04992_));
 NAND2x1_ASAP7_75t_R _27412_ (.A(net4731),
    .B(net4853),
    .Y(_04993_));
 AOI22x1_ASAP7_75t_R _27413_ (.A1(_04993_),
    .A2(net6092),
    .B1(_04556_),
    .B2(net4634),
    .Y(_04994_));
 OA21x2_ASAP7_75t_R _27414_ (.A1(net6102),
    .A2(net4730),
    .B(net5646),
    .Y(_04995_));
 NAND2x1_ASAP7_75t_R _27415_ (.A(_04763_),
    .B(_04543_),
    .Y(_04996_));
 AOI21x1_ASAP7_75t_R _27416_ (.A1(_04995_),
    .A2(_04996_),
    .B(net6101),
    .Y(_04997_));
 OAI21x1_ASAP7_75t_R _27417_ (.A1(net5651),
    .A2(_04994_),
    .B(_04997_),
    .Y(_04998_));
 NOR2x1_ASAP7_75t_R _27418_ (.A(net4498),
    .B(_04617_),
    .Y(_04999_));
 NOR2x1_ASAP7_75t_R _27419_ (.A(_04611_),
    .B(_04868_),
    .Y(_05000_));
 OAI21x1_ASAP7_75t_R _27420_ (.A1(_05000_),
    .A2(_04999_),
    .B(net5659),
    .Y(_05001_));
 NAND2x1_ASAP7_75t_R _27421_ (.A(net6091),
    .B(net4862),
    .Y(_05002_));
 OAI21x1_ASAP7_75t_R _27422_ (.A1(_04693_),
    .A2(_04868_),
    .B(_05002_),
    .Y(_05003_));
 AOI21x1_ASAP7_75t_R _27423_ (.A1(net5651),
    .A2(_05003_),
    .B(net5658),
    .Y(_05004_));
 NAND2x1_ASAP7_75t_R _27424_ (.A(_05004_),
    .B(_05001_),
    .Y(_05005_));
 AOI21x1_ASAP7_75t_R _27425_ (.A1(_04998_),
    .A2(_05005_),
    .B(_04536_),
    .Y(_05006_));
 AOI21x1_ASAP7_75t_R _27426_ (.A1(net4639),
    .A2(_04513_),
    .B(net6093),
    .Y(_05007_));
 AOI21x1_ASAP7_75t_R _27427_ (.A1(_04734_),
    .A2(_04658_),
    .B(net6107),
    .Y(_05008_));
 OAI21x1_ASAP7_75t_R _27428_ (.A1(_05007_),
    .A2(net4497),
    .B(net5661),
    .Y(_05009_));
 AO21x1_ASAP7_75t_R _27429_ (.A1(net5380),
    .A2(net5656),
    .B(_04771_),
    .Y(_05010_));
 AOI21x1_ASAP7_75t_R _27430_ (.A1(net4638),
    .A2(_05010_),
    .B(net6092),
    .Y(_05011_));
 NOR2x1_ASAP7_75t_R _27431_ (.A(_04504_),
    .B(_04617_),
    .Y(_05012_));
 OAI21x1_ASAP7_75t_R _27432_ (.A1(_05011_),
    .A2(_05012_),
    .B(net5655),
    .Y(_05013_));
 AOI21x1_ASAP7_75t_R _27433_ (.A1(_05009_),
    .A2(_05013_),
    .B(net5658),
    .Y(_05014_));
 AOI21x1_ASAP7_75t_R _27434_ (.A1(net4638),
    .A2(net4853),
    .B(net6092),
    .Y(_05015_));
 OAI21x1_ASAP7_75t_R _27435_ (.A1(_05015_),
    .A2(_04855_),
    .B(net5658),
    .Y(_05016_));
 NAND2x1_ASAP7_75t_R _27436_ (.A(_01312_),
    .B(_01316_),
    .Y(_05017_));
 AOI21x1_ASAP7_75t_R _27437_ (.A1(net6091),
    .A2(_05017_),
    .B(net5654),
    .Y(_05018_));
 OA21x2_ASAP7_75t_R _27438_ (.A1(_04863_),
    .A2(net6091),
    .B(_05018_),
    .Y(_05019_));
 OAI21x1_ASAP7_75t_R _27439_ (.A1(_05016_),
    .A2(_05019_),
    .B(net5644),
    .Y(_05020_));
 OAI21x1_ASAP7_75t_R _27440_ (.A1(_05020_),
    .A2(_05014_),
    .B(net5643),
    .Y(_05021_));
 OAI22x1_ASAP7_75t_R _27441_ (.A1(_04977_),
    .A2(_04992_),
    .B1(_05006_),
    .B2(_05021_),
    .Y(_00126_));
 NAND2x1_ASAP7_75t_R _27442_ (.A(net4858),
    .B(_04548_),
    .Y(_05022_));
 AO21x1_ASAP7_75t_R _27443_ (.A1(net4731),
    .A2(net4549),
    .B(net6098),
    .Y(_05023_));
 AO21x1_ASAP7_75t_R _27444_ (.A1(_05022_),
    .A2(_05023_),
    .B(net5661),
    .Y(_05024_));
 AO21x1_ASAP7_75t_R _27445_ (.A1(_04585_),
    .A2(_04447_),
    .B(net6106),
    .Y(_05025_));
 OR2x2_ASAP7_75t_R _27446_ (.A(_01316_),
    .B(net6091),
    .Y(_05026_));
 AO21x1_ASAP7_75t_R _27447_ (.A1(_05025_),
    .A2(_05026_),
    .B(net5653),
    .Y(_05027_));
 AOI21x1_ASAP7_75t_R _27448_ (.A1(_05024_),
    .A2(_05027_),
    .B(net5658),
    .Y(_05028_));
 NOR2x1_ASAP7_75t_R _27449_ (.A(net5039),
    .B(net5102),
    .Y(_05029_));
 AOI21x1_ASAP7_75t_R _27450_ (.A1(net6091),
    .A2(_05029_),
    .B(net5655),
    .Y(_05030_));
 NAND2x1_ASAP7_75t_R _27451_ (.A(net5033),
    .B(net6107),
    .Y(_05031_));
 AO21x1_ASAP7_75t_R _27452_ (.A1(_05030_),
    .A2(_05031_),
    .B(net6101),
    .Y(_05032_));
 AND3x1_ASAP7_75t_R _27453_ (.A(_04691_),
    .B(_04889_),
    .C(_04564_),
    .Y(_05033_));
 OAI21x1_ASAP7_75t_R _27454_ (.A1(_05032_),
    .A2(_05033_),
    .B(net5643),
    .Y(_05034_));
 OAI21x1_ASAP7_75t_R _27455_ (.A1(_05028_),
    .A2(_05034_),
    .B(net6089),
    .Y(_05035_));
 AO21x1_ASAP7_75t_R _27456_ (.A1(_04753_),
    .A2(_04513_),
    .B(net6106),
    .Y(_05036_));
 AOI21x1_ASAP7_75t_R _27457_ (.A1(_04786_),
    .A2(_05036_),
    .B(net6101),
    .Y(_05037_));
 NAND2x1_ASAP7_75t_R _27458_ (.A(net5378),
    .B(net6092),
    .Y(_05038_));
 AO21x1_ASAP7_75t_R _27459_ (.A1(_04903_),
    .A2(_05038_),
    .B(net5661),
    .Y(_05039_));
 NAND2x1_ASAP7_75t_R _27460_ (.A(_04957_),
    .B(_04917_),
    .Y(_05040_));
 INVx1_ASAP7_75t_R _27461_ (.A(_04868_),
    .Y(_05041_));
 AOI21x1_ASAP7_75t_R _27462_ (.A1(net4730),
    .A2(_04513_),
    .B(net6107),
    .Y(_05042_));
 OAI21x1_ASAP7_75t_R _27463_ (.A1(_05041_),
    .A2(_05042_),
    .B(net5654),
    .Y(_05043_));
 AOI21x1_ASAP7_75t_R _27464_ (.A1(_05040_),
    .A2(_05043_),
    .B(net5658),
    .Y(_05044_));
 AOI211x1_ASAP7_75t_R _27465_ (.A1(_05037_),
    .A2(_05039_),
    .B(_05044_),
    .C(net5643),
    .Y(_05045_));
 OA21x2_ASAP7_75t_R _27466_ (.A1(net5034),
    .A2(net6107),
    .B(net5655),
    .Y(_05046_));
 OAI21x1_ASAP7_75t_R _27467_ (.A1(net6091),
    .A2(_04863_),
    .B(_05046_),
    .Y(_05047_));
 AOI21x1_ASAP7_75t_R _27468_ (.A1(net6107),
    .A2(_04563_),
    .B(_04482_),
    .Y(_05048_));
 AOI21x1_ASAP7_75t_R _27469_ (.A1(_05030_),
    .A2(_05048_),
    .B(net5658),
    .Y(_05049_));
 AOI21x1_ASAP7_75t_R _27470_ (.A1(_05047_),
    .A2(_05049_),
    .B(net6088),
    .Y(_05050_));
 OAI21x1_ASAP7_75t_R _27471_ (.A1(_04806_),
    .A2(net4862),
    .B(net6102),
    .Y(_05051_));
 OAI21x1_ASAP7_75t_R _27472_ (.A1(_04482_),
    .A2(_04770_),
    .B(net6094),
    .Y(_05052_));
 AOI21x1_ASAP7_75t_R _27473_ (.A1(_05051_),
    .A2(_05052_),
    .B(net5651),
    .Y(_05053_));
 OAI21x1_ASAP7_75t_R _27474_ (.A1(_04770_),
    .A2(_04663_),
    .B(net6094),
    .Y(_05054_));
 AOI21x1_ASAP7_75t_R _27475_ (.A1(_04811_),
    .A2(_05054_),
    .B(net5659),
    .Y(_05055_));
 OAI21x1_ASAP7_75t_R _27476_ (.A1(_05053_),
    .A2(_05055_),
    .B(net5658),
    .Y(_05056_));
 AOI21x1_ASAP7_75t_R _27477_ (.A1(_05050_),
    .A2(_05056_),
    .B(net6089),
    .Y(_05057_));
 INVx1_ASAP7_75t_R _27478_ (.A(_05008_),
    .Y(_05058_));
 AOI21x1_ASAP7_75t_R _27479_ (.A1(_04780_),
    .A2(_05058_),
    .B(net5652),
    .Y(_05059_));
 NAND2x1_ASAP7_75t_R _27480_ (.A(net4731),
    .B(_04548_),
    .Y(_05060_));
 AOI21x1_ASAP7_75t_R _27481_ (.A1(_05060_),
    .A2(_04659_),
    .B(net5661),
    .Y(_05061_));
 OAI21x1_ASAP7_75t_R _27482_ (.A1(_05059_),
    .A2(_05061_),
    .B(net6101),
    .Y(_05062_));
 AO21x1_ASAP7_75t_R _27483_ (.A1(_04971_),
    .A2(net4855),
    .B(net6107),
    .Y(_05063_));
 NOR2x1_ASAP7_75t_R _27484_ (.A(_04512_),
    .B(_04851_),
    .Y(_05064_));
 NOR2x1_ASAP7_75t_R _27485_ (.A(_04710_),
    .B(_05064_),
    .Y(_05065_));
 NAND2x1_ASAP7_75t_R _27486_ (.A(_05063_),
    .B(_05065_),
    .Y(_05066_));
 AOI21x1_ASAP7_75t_R _27487_ (.A1(net6097),
    .A2(_04555_),
    .B(net5649),
    .Y(_05067_));
 AOI21x1_ASAP7_75t_R _27488_ (.A1(_05067_),
    .A2(_04890_),
    .B(net6100),
    .Y(_05068_));
 AOI21x1_ASAP7_75t_R _27489_ (.A1(_05066_),
    .A2(_05068_),
    .B(_04849_),
    .Y(_05069_));
 NAND2x1_ASAP7_75t_R _27490_ (.A(_05062_),
    .B(_05069_),
    .Y(_05070_));
 NAND2x1_ASAP7_75t_R _27491_ (.A(_05057_),
    .B(_05070_),
    .Y(_05071_));
 OAI21x1_ASAP7_75t_R _27492_ (.A1(_05035_),
    .A2(_05045_),
    .B(_05071_),
    .Y(_00127_));
 NOR2x1_ASAP7_75t_R _27493_ (.A(net6672),
    .B(_00480_),
    .Y(_05072_));
 XOR2x2_ASAP7_75t_R _27494_ (.A(net6453),
    .B(net6597),
    .Y(_05073_));
 XOR2x2_ASAP7_75t_R _27495_ (.A(_10717_),
    .B(_02281_),
    .Y(_05074_));
 NAND2x1_ASAP7_75t_R _27496_ (.A(_05073_),
    .B(_05074_),
    .Y(_05075_));
 XNOR2x2_ASAP7_75t_R _27497_ (.A(net6597),
    .B(net6453),
    .Y(_05076_));
 XOR2x2_ASAP7_75t_R _27498_ (.A(_02281_),
    .B(_10719_),
    .Y(_05077_));
 NAND2x1p5_ASAP7_75t_R _27499_ (.A(_05076_),
    .B(_05077_),
    .Y(_05078_));
 AOI21x1_ASAP7_75t_R _27500_ (.A1(_05075_),
    .A2(_05078_),
    .B(net6462),
    .Y(_05079_));
 OAI21x1_ASAP7_75t_R _27501_ (.A1(_05072_),
    .A2(_05079_),
    .B(net6529),
    .Y(_05080_));
 AND2x2_ASAP7_75t_R _27502_ (.A(net6462),
    .B(_00480_),
    .Y(_05081_));
 NAND2x1_ASAP7_75t_R _27503_ (.A(_05073_),
    .B(_05077_),
    .Y(_05082_));
 NAND2x1p5_ASAP7_75t_R _27504_ (.A(_05074_),
    .B(_05076_),
    .Y(_05083_));
 AOI21x1_ASAP7_75t_R _27505_ (.A1(_05082_),
    .A2(_05083_),
    .B(net6462),
    .Y(_05084_));
 INVx1_ASAP7_75t_R _27506_ (.A(net6529),
    .Y(_05085_));
 OAI21x1_ASAP7_75t_R _27507_ (.A1(_05081_),
    .A2(_05084_),
    .B(_05085_),
    .Y(_05086_));
 NAND2x1p5_ASAP7_75t_R _27508_ (.A(_05080_),
    .B(_05086_),
    .Y(_05087_));
 OR2x2_ASAP7_75t_R _27510_ (.A(net6668),
    .B(_00481_),
    .Y(_05088_));
 NOR2x1_ASAP7_75t_R _27511_ (.A(_10858_),
    .B(_10701_),
    .Y(_05089_));
 NOR2x1p5_ASAP7_75t_R _27512_ (.A(net6560),
    .B(_10702_),
    .Y(_05090_));
 OAI21x1_ASAP7_75t_R _27513_ (.A1(_05089_),
    .A2(_05090_),
    .B(net6452),
    .Y(_05091_));
 INVx1_ASAP7_75t_R _27514_ (.A(_05091_),
    .Y(_05092_));
 NOR3x1_ASAP7_75t_R _27515_ (.A(net6382),
    .B(_05089_),
    .C(net6452),
    .Y(_05093_));
 OAI21x1_ASAP7_75t_R _27516_ (.A1(_05092_),
    .A2(_05093_),
    .B(net6668),
    .Y(_05094_));
 AOI21x1_ASAP7_75t_R _27517_ (.A1(_05088_),
    .A2(_05094_),
    .B(net6539),
    .Y(_05095_));
 NAND2x1_ASAP7_75t_R _27518_ (.A(_00481_),
    .B(net6462),
    .Y(_05096_));
 INVx1_ASAP7_75t_R _27519_ (.A(net6453),
    .Y(_05097_));
 XOR2x2_ASAP7_75t_R _27520_ (.A(_10701_),
    .B(_10858_),
    .Y(_05098_));
 NAND2x1_ASAP7_75t_R _27521_ (.A(_05097_),
    .B(_05098_),
    .Y(_05099_));
 NAND3x1_ASAP7_75t_R _27522_ (.A(_05091_),
    .B(net6668),
    .C(_05099_),
    .Y(_05100_));
 INVx1_ASAP7_75t_R _27523_ (.A(net6539),
    .Y(_05101_));
 AOI21x1_ASAP7_75t_R _27524_ (.A1(_05096_),
    .A2(net6087),
    .B(_05101_),
    .Y(_05102_));
 NOR2x1_ASAP7_75t_R _27525_ (.A(_05095_),
    .B(_05102_),
    .Y(_05103_));
 XOR2x2_ASAP7_75t_R _27527_ (.A(net6647),
    .B(net6596),
    .Y(_05104_));
 NAND2x1_ASAP7_75t_R _27528_ (.A(net6402),
    .B(_05104_),
    .Y(_05105_));
 XNOR2x2_ASAP7_75t_R _27529_ (.A(net6647),
    .B(net6596),
    .Y(_05106_));
 NAND2x1_ASAP7_75t_R _27530_ (.A(net6565),
    .B(_05106_),
    .Y(_05107_));
 AOI21x1_ASAP7_75t_R _27531_ (.A1(_05105_),
    .A2(_05107_),
    .B(_02331_),
    .Y(_05108_));
 XOR2x2_ASAP7_75t_R _27532_ (.A(net6596),
    .B(net6565),
    .Y(_05109_));
 NAND2x1_ASAP7_75t_R _27533_ (.A(net6647),
    .B(_05109_),
    .Y(_05110_));
 XNOR2x2_ASAP7_75t_R _27534_ (.A(net6596),
    .B(net6565),
    .Y(_05111_));
 NAND2x1_ASAP7_75t_R _27535_ (.A(net6419),
    .B(_05111_),
    .Y(_05112_));
 AOI21x1_ASAP7_75t_R _27536_ (.A1(_05110_),
    .A2(_05112_),
    .B(_02319_),
    .Y(_05113_));
 OAI21x1_ASAP7_75t_R _27537_ (.A1(_05108_),
    .A2(_05113_),
    .B(net6672),
    .Y(_05114_));
 NOR2x1_ASAP7_75t_R _27538_ (.A(net6672),
    .B(_00482_),
    .Y(_05115_));
 INVx1_ASAP7_75t_R _27539_ (.A(_05115_),
    .Y(_05116_));
 NAND3x1_ASAP7_75t_R _27540_ (.A(_05114_),
    .B(net6522),
    .C(_05116_),
    .Y(_05117_));
 AO21x1_ASAP7_75t_R _27541_ (.A1(_05114_),
    .A2(_05116_),
    .B(net6522),
    .Y(_05118_));
 NAND2x1_ASAP7_75t_R _27542_ (.A(_05117_),
    .B(_05118_),
    .Y(_05119_));
 AOI21x1_ASAP7_75t_R _27545_ (.A1(_05088_),
    .A2(_05094_),
    .B(_05101_),
    .Y(_05121_));
 AOI21x1_ASAP7_75t_R _27546_ (.A1(_05096_),
    .A2(_05100_),
    .B(net6539),
    .Y(_05122_));
 NOR2x1p5_ASAP7_75t_R _27547_ (.A(_05122_),
    .B(_05121_),
    .Y(_05123_));
 INVx1_ASAP7_75t_R _27549_ (.A(net6522),
    .Y(_05124_));
 NAND3x1_ASAP7_75t_R _27550_ (.A(_05114_),
    .B(_05124_),
    .C(_05116_),
    .Y(_05125_));
 AO21x1_ASAP7_75t_R _27551_ (.A1(_05114_),
    .A2(_05116_),
    .B(_05124_),
    .Y(_05126_));
 NAND2x1_ASAP7_75t_R _27552_ (.A(_05125_),
    .B(_05126_),
    .Y(_05127_));
 AO21x1_ASAP7_75t_R _27556_ (.A1(net6083),
    .A2(net6084),
    .B(_01323_),
    .Y(_05130_));
 INVx1_ASAP7_75t_R _27558_ (.A(_01327_),
    .Y(_05132_));
 XNOR2x2_ASAP7_75t_R _27559_ (.A(net6595),
    .B(_10757_),
    .Y(_05133_));
 NOR2x1_ASAP7_75t_R _27560_ (.A(_05133_),
    .B(_02364_),
    .Y(_05134_));
 XOR2x2_ASAP7_75t_R _27561_ (.A(_10757_),
    .B(net6595),
    .Y(_05135_));
 XNOR2x2_ASAP7_75t_R _27562_ (.A(_02363_),
    .B(_02362_),
    .Y(_05136_));
 OAI21x1_ASAP7_75t_R _27563_ (.A1(_05135_),
    .A2(_05136_),
    .B(net6672),
    .Y(_05137_));
 NAND2x1_ASAP7_75t_R _27564_ (.A(_00489_),
    .B(net6462),
    .Y(_05138_));
 OAI21x1_ASAP7_75t_R _27565_ (.A1(_05134_),
    .A2(_05137_),
    .B(_05138_),
    .Y(_05139_));
 XOR2x2_ASAP7_75t_R _27566_ (.A(_05139_),
    .B(net6519),
    .Y(_05140_));
 AOI21x1_ASAP7_75t_R _27568_ (.A1(_05132_),
    .A2(net5639),
    .B(net6077),
    .Y(_05142_));
 NAND2x1_ASAP7_75t_R _27569_ (.A(_05130_),
    .B(_05142_),
    .Y(_05143_));
 AO21x1_ASAP7_75t_R _27572_ (.A1(net6085),
    .A2(net6086),
    .B(_01323_),
    .Y(_05146_));
 XNOR2x2_ASAP7_75t_R _27573_ (.A(net6519),
    .B(_05139_),
    .Y(_05147_));
 INVx1_ASAP7_75t_R _27575_ (.A(_01324_),
    .Y(_05149_));
 AOI21x1_ASAP7_75t_R _27576_ (.A1(net6084),
    .A2(net6083),
    .B(_05149_),
    .Y(_05150_));
 NOR2x1p5_ASAP7_75t_R _27577_ (.A(_05150_),
    .B(_05147_),
    .Y(_05151_));
 NAND2x1_ASAP7_75t_R _27578_ (.A(_05146_),
    .B(_05151_),
    .Y(_05152_));
 XNOR2x2_ASAP7_75t_R _27579_ (.A(_00643_),
    .B(_10773_),
    .Y(_05153_));
 XOR2x2_ASAP7_75t_R _27580_ (.A(_05153_),
    .B(_02351_),
    .Y(_05154_));
 NOR2x1_ASAP7_75t_R _27581_ (.A(net6668),
    .B(_00568_),
    .Y(_05155_));
 AOI21x1_ASAP7_75t_R _27582_ (.A1(net6668),
    .A2(_05154_),
    .B(_05155_),
    .Y(_05156_));
 XOR2x2_ASAP7_75t_R _27583_ (.A(_05156_),
    .B(net6518),
    .Y(_05157_));
 AO21x1_ASAP7_75t_R _27585_ (.A1(_05143_),
    .A2(_05152_),
    .B(net6068),
    .Y(_05159_));
 NAND2x1_ASAP7_75t_R _27587_ (.A(net5638),
    .B(net5641),
    .Y(_05161_));
 AO21x2_ASAP7_75t_R _27588_ (.A1(net6083),
    .A2(net6084),
    .B(net4721),
    .Y(_05162_));
 AO21x1_ASAP7_75t_R _27591_ (.A1(net5377),
    .A2(_05162_),
    .B(net6078),
    .Y(_05165_));
 NOR2x1_ASAP7_75t_R _27594_ (.A(net4546),
    .B(net5636),
    .Y(_05168_));
 NAND2x1_ASAP7_75t_R _27595_ (.A(net6078),
    .B(_05168_),
    .Y(_05169_));
 XNOR2x2_ASAP7_75t_R _27596_ (.A(net6518),
    .B(_05156_),
    .Y(_05170_));
 AO21x1_ASAP7_75t_R _27599_ (.A1(_05165_),
    .A2(_05169_),
    .B(net6065),
    .Y(_05173_));
 XOR2x2_ASAP7_75t_R _27600_ (.A(_00579_),
    .B(_00580_),
    .Y(_05174_));
 XOR2x2_ASAP7_75t_R _27601_ (.A(_10802_),
    .B(net6562),
    .Y(_05175_));
 NAND2x1_ASAP7_75t_R _27602_ (.A(_05174_),
    .B(_05175_),
    .Y(_05176_));
 INVx1_ASAP7_75t_R _27603_ (.A(_05174_),
    .Y(_05177_));
 XNOR2x2_ASAP7_75t_R _27604_ (.A(net6562),
    .B(_10802_),
    .Y(_05178_));
 NAND2x1_ASAP7_75t_R _27605_ (.A(_05177_),
    .B(_05178_),
    .Y(_05179_));
 AOI21x1_ASAP7_75t_R _27606_ (.A1(_05176_),
    .A2(_05179_),
    .B(net6462),
    .Y(_05180_));
 NOR2x1_ASAP7_75t_R _27607_ (.A(net6668),
    .B(_00567_),
    .Y(_05181_));
 INVx1_ASAP7_75t_R _27608_ (.A(net6517),
    .Y(_05182_));
 OA21x2_ASAP7_75t_R _27609_ (.A1(_05180_),
    .A2(_05181_),
    .B(_05182_),
    .Y(_05183_));
 INVx1_ASAP7_75t_R _27610_ (.A(_00567_),
    .Y(_05184_));
 AOI211x1_ASAP7_75t_R _27611_ (.A1(net6462),
    .A2(_05184_),
    .B(_05180_),
    .C(_05182_),
    .Y(_05185_));
 NOR2x1_ASAP7_75t_R _27612_ (.A(_05183_),
    .B(_05185_),
    .Y(_05186_));
 AOI21x1_ASAP7_75t_R _27615_ (.A1(_05159_),
    .A2(_05173_),
    .B(net5633),
    .Y(_05189_));
 AO21x1_ASAP7_75t_R _27616_ (.A1(net5097),
    .A2(net5641),
    .B(net5637),
    .Y(_05190_));
 AOI21x1_ASAP7_75t_R _27619_ (.A1(net4544),
    .A2(_05190_),
    .B(net6077),
    .Y(_05193_));
 INVx1_ASAP7_75t_R _27621_ (.A(_01323_),
    .Y(_05195_));
 AO21x1_ASAP7_75t_R _27622_ (.A1(net6085),
    .A2(net6086),
    .B(_05195_),
    .Y(_05196_));
 AO21x1_ASAP7_75t_R _27623_ (.A1(net6083),
    .A2(net6084),
    .B(_05132_),
    .Y(_05197_));
 AO21x1_ASAP7_75t_R _27625_ (.A1(_05196_),
    .A2(_05197_),
    .B(net6073),
    .Y(_05199_));
 NAND2x1_ASAP7_75t_R _27626_ (.A(net6064),
    .B(_05199_),
    .Y(_05200_));
 OAI21x1_ASAP7_75t_R _27628_ (.A1(_05193_),
    .A2(_05200_),
    .B(net5633),
    .Y(_05202_));
 INVx3_ASAP7_75t_R _27629_ (.A(_05087_),
    .Y(_01321_));
 NAND2x1_ASAP7_75t_R _27630_ (.A(net5096),
    .B(net5373),
    .Y(_05203_));
 AOI21x1_ASAP7_75t_R _27631_ (.A1(net5637),
    .A2(net5097),
    .B(net6077),
    .Y(_05204_));
 NAND2x1_ASAP7_75t_R _27632_ (.A(_05203_),
    .B(_05204_),
    .Y(_05205_));
 NAND2x1_ASAP7_75t_R _27633_ (.A(net5638),
    .B(net5097),
    .Y(_05206_));
 AOI21x1_ASAP7_75t_R _27636_ (.A1(net5641),
    .A2(net5095),
    .B(net6073),
    .Y(_05209_));
 NAND2x1_ASAP7_75t_R _27637_ (.A(_05206_),
    .B(_05209_),
    .Y(_05210_));
 AND3x1_ASAP7_75t_R _27639_ (.A(_05205_),
    .B(_05210_),
    .C(net6068),
    .Y(_05212_));
 XOR2x2_ASAP7_75t_R _27640_ (.A(_00580_),
    .B(_00581_),
    .Y(_05213_));
 XOR2x2_ASAP7_75t_R _27641_ (.A(_05213_),
    .B(_10803_),
    .Y(_05214_));
 XOR2x2_ASAP7_75t_R _27642_ (.A(_05214_),
    .B(_10744_),
    .Y(_05215_));
 NOR2x1_ASAP7_75t_R _27643_ (.A(net6668),
    .B(_00566_),
    .Y(_05216_));
 AO21x1_ASAP7_75t_R _27644_ (.A1(_05215_),
    .A2(net6668),
    .B(_05216_),
    .Y(_05217_));
 XOR2x2_ASAP7_75t_R _27645_ (.A(_05217_),
    .B(net6516),
    .Y(_05218_));
 OAI21x1_ASAP7_75t_R _27647_ (.A1(_05202_),
    .A2(_05212_),
    .B(net6060),
    .Y(_05220_));
 NOR2x1_ASAP7_75t_R _27648_ (.A(_05189_),
    .B(_05220_),
    .Y(_05221_));
 INVx1_ASAP7_75t_R _27649_ (.A(_01332_),
    .Y(_05222_));
 AO21x1_ASAP7_75t_R _27650_ (.A1(net6085),
    .A2(net6086),
    .B(_05222_),
    .Y(_05223_));
 NAND2x1_ASAP7_75t_R _27651_ (.A(net6082),
    .B(_05223_),
    .Y(_05224_));
 NAND2x1_ASAP7_75t_R _27652_ (.A(net5640),
    .B(net5095),
    .Y(_05225_));
 AOI21x1_ASAP7_75t_R _27653_ (.A1(net5636),
    .A2(net5095),
    .B(net6079),
    .Y(_05226_));
 AOI21x1_ASAP7_75t_R _27655_ (.A1(net4845),
    .A2(_05226_),
    .B(net6063),
    .Y(_05228_));
 OA21x2_ASAP7_75t_R _27656_ (.A1(net4458),
    .A2(net4439),
    .B(_05228_),
    .Y(_05229_));
 AOI21x1_ASAP7_75t_R _27657_ (.A1(net5638),
    .A2(net5095),
    .B(net6082),
    .Y(_05230_));
 INVx1_ASAP7_75t_R _27658_ (.A(_05230_),
    .Y(_05231_));
 NAND2x1_ASAP7_75t_R _27659_ (.A(net6065),
    .B(_05231_),
    .Y(_05232_));
 INVx1_ASAP7_75t_R _27660_ (.A(net4800),
    .Y(_05233_));
 OA21x2_ASAP7_75t_R _27661_ (.A1(net5638),
    .A2(_05233_),
    .B(net6079),
    .Y(_05234_));
 OA21x2_ASAP7_75t_R _27662_ (.A1(net5637),
    .A2(net4845),
    .B(_05234_),
    .Y(_05235_));
 OAI21x1_ASAP7_75t_R _27663_ (.A1(_05232_),
    .A2(_05235_),
    .B(net5634),
    .Y(_05236_));
 INVx1_ASAP7_75t_R _27664_ (.A(_05218_),
    .Y(_05237_));
 OAI21x1_ASAP7_75t_R _27665_ (.A1(_05229_),
    .A2(_05236_),
    .B(_05237_),
    .Y(_05238_));
 OAI21x1_ASAP7_75t_R _27668_ (.A1(net5097),
    .A2(net5376),
    .B(net6073),
    .Y(_05241_));
 NOR2x1_ASAP7_75t_R _27669_ (.A(net5638),
    .B(net5640),
    .Y(_05242_));
 AO21x1_ASAP7_75t_R _27670_ (.A1(net6083),
    .A2(net6084),
    .B(net4630),
    .Y(_05243_));
 AOI21x1_ASAP7_75t_R _27671_ (.A1(net5638),
    .A2(net5095),
    .B(net6074),
    .Y(_05244_));
 NAND2x1_ASAP7_75t_R _27672_ (.A(net4496),
    .B(_05244_),
    .Y(_05245_));
 OA21x2_ASAP7_75t_R _27673_ (.A1(_05241_),
    .A2(net5372),
    .B(_05245_),
    .Y(_05246_));
 INVx1_ASAP7_75t_R _27674_ (.A(_05244_),
    .Y(_05247_));
 NAND2x1_ASAP7_75t_R _27675_ (.A(_05127_),
    .B(net5640),
    .Y(_05248_));
 NOR2x1_ASAP7_75t_R _27676_ (.A(net5095),
    .B(net5371),
    .Y(_05249_));
 NOR2x1_ASAP7_75t_R _27677_ (.A(net6402),
    .B(_05104_),
    .Y(_05250_));
 NOR2x1_ASAP7_75t_R _27678_ (.A(net6565),
    .B(_05106_),
    .Y(_05251_));
 OAI21x1_ASAP7_75t_R _27679_ (.A1(_05250_),
    .A2(_05251_),
    .B(_02319_),
    .Y(_05252_));
 NOR2x1_ASAP7_75t_R _27680_ (.A(net6647),
    .B(_05109_),
    .Y(_05253_));
 NOR2x1_ASAP7_75t_R _27681_ (.A(net6419),
    .B(_05111_),
    .Y(_05254_));
 OAI21x1_ASAP7_75t_R _27682_ (.A1(_05253_),
    .A2(_05254_),
    .B(_02331_),
    .Y(_05255_));
 AOI21x1_ASAP7_75t_R _27683_ (.A1(_05252_),
    .A2(_05255_),
    .B(net6462),
    .Y(_05256_));
 NOR3x1_ASAP7_75t_R _27684_ (.A(_05256_),
    .B(net6522),
    .C(net6394),
    .Y(_05257_));
 OA21x2_ASAP7_75t_R _27685_ (.A1(_05256_),
    .A2(net6394),
    .B(net6522),
    .Y(_05258_));
 INVx1_ASAP7_75t_R _27686_ (.A(_01325_),
    .Y(_05259_));
 OAI21x1_ASAP7_75t_R _27687_ (.A1(_05257_),
    .A2(_05258_),
    .B(_05259_),
    .Y(_05260_));
 INVx1_ASAP7_75t_R _27688_ (.A(_05260_),
    .Y(_05261_));
 NOR2x1_ASAP7_75t_R _27689_ (.A(net5637),
    .B(net5641),
    .Y(_05262_));
 OAI21x1_ASAP7_75t_R _27691_ (.A1(_05261_),
    .A2(net5368),
    .B(net6075),
    .Y(_05264_));
 OAI21x1_ASAP7_75t_R _27692_ (.A1(_05247_),
    .A2(_05249_),
    .B(_05264_),
    .Y(_05265_));
 INVx1_ASAP7_75t_R _27693_ (.A(_05186_),
    .Y(_05266_));
 OAI21x1_ASAP7_75t_R _27696_ (.A1(net6069),
    .A2(_05265_),
    .B(net5366),
    .Y(_05269_));
 AOI21x1_ASAP7_75t_R _27697_ (.A1(net6069),
    .A2(_05246_),
    .B(_05269_),
    .Y(_05270_));
 XOR2x2_ASAP7_75t_R _27698_ (.A(_00581_),
    .B(net6644),
    .Y(_05271_));
 XOR2x2_ASAP7_75t_R _27699_ (.A(_05271_),
    .B(_00677_),
    .Y(_05272_));
 XOR2x2_ASAP7_75t_R _27700_ (.A(_05272_),
    .B(_10860_),
    .Y(_05273_));
 NOR2x1_ASAP7_75t_R _27701_ (.A(net6671),
    .B(_00565_),
    .Y(_05274_));
 AO21x1_ASAP7_75t_R _27702_ (.A1(_05273_),
    .A2(net6671),
    .B(_05274_),
    .Y(_05275_));
 XOR2x2_ASAP7_75t_R _27703_ (.A(_05275_),
    .B(net6515),
    .Y(_05276_));
 OAI21x1_ASAP7_75t_R _27705_ (.A1(_05238_),
    .A2(_05270_),
    .B(net6059),
    .Y(_05278_));
 INVx1_ASAP7_75t_R _27706_ (.A(_01340_),
    .Y(_05279_));
 AO21x1_ASAP7_75t_R _27708_ (.A1(net6085),
    .A2(net6086),
    .B(net4721),
    .Y(_05281_));
 NAND2x1_ASAP7_75t_R _27710_ (.A(net6073),
    .B(_05281_),
    .Y(_05283_));
 OAI21x1_ASAP7_75t_R _27711_ (.A1(_05279_),
    .A2(net6072),
    .B(_05283_),
    .Y(_05284_));
 AOI21x1_ASAP7_75t_R _27713_ (.A1(_05130_),
    .A2(_05244_),
    .B(net6069),
    .Y(_05286_));
 AND2x2_ASAP7_75t_R _27714_ (.A(_01325_),
    .B(_01330_),
    .Y(_05287_));
 NOR2x1_ASAP7_75t_R _27715_ (.A(net4629),
    .B(net5636),
    .Y(_05288_));
 AOI21x1_ASAP7_75t_R _27716_ (.A1(net5640),
    .A2(net5095),
    .B(net5639),
    .Y(_05289_));
 OAI21x1_ASAP7_75t_R _27717_ (.A1(_05288_),
    .A2(_05289_),
    .B(net6072),
    .Y(_05290_));
 AOI221x1_ASAP7_75t_R _27718_ (.A1(net6068),
    .A2(_05284_),
    .B1(_05286_),
    .B2(_05290_),
    .C(net5635),
    .Y(_05291_));
 NOR2x1_ASAP7_75t_R _27719_ (.A(net6075),
    .B(_05260_),
    .Y(_05292_));
 NOR2x1_ASAP7_75t_R _27720_ (.A(net6065),
    .B(_05292_),
    .Y(_05293_));
 INVx1_ASAP7_75t_R _27721_ (.A(_05293_),
    .Y(_05294_));
 INVx1_ASAP7_75t_R _27722_ (.A(_05142_),
    .Y(_05295_));
 NOR2x1_ASAP7_75t_R _27723_ (.A(net5099),
    .B(net5371),
    .Y(_05296_));
 NOR2x1_ASAP7_75t_R _27724_ (.A(_05295_),
    .B(_05296_),
    .Y(_05297_));
 OAI21x1_ASAP7_75t_R _27725_ (.A1(_05294_),
    .A2(_05297_),
    .B(net5632),
    .Y(_05298_));
 AOI21x1_ASAP7_75t_R _27727_ (.A1(net4801),
    .A2(net5639),
    .B(net6073),
    .Y(_05300_));
 INVx1_ASAP7_75t_R _27728_ (.A(_05300_),
    .Y(_05301_));
 NAND2x1_ASAP7_75t_R _27729_ (.A(net6075),
    .B(_05261_),
    .Y(_05302_));
 OA211x2_ASAP7_75t_R _27730_ (.A1(_05296_),
    .A2(_05301_),
    .B(_05302_),
    .C(net6061),
    .Y(_05303_));
 OAI21x1_ASAP7_75t_R _27731_ (.A1(_05298_),
    .A2(_05303_),
    .B(net6060),
    .Y(_05304_));
 AOI21x1_ASAP7_75t_R _27732_ (.A1(net5636),
    .A2(net5640),
    .B(_05140_),
    .Y(_05305_));
 NAND2x1_ASAP7_75t_R _27733_ (.A(net4543),
    .B(net5365),
    .Y(_05306_));
 INVx1_ASAP7_75t_R _27734_ (.A(_05306_),
    .Y(_05307_));
 AO21x1_ASAP7_75t_R _27735_ (.A1(net6085),
    .A2(net6086),
    .B(net4802),
    .Y(_05308_));
 AND2x2_ASAP7_75t_R _27736_ (.A(_05308_),
    .B(net6077),
    .Y(_05309_));
 NAND2x1_ASAP7_75t_R _27737_ (.A(net5636),
    .B(net5095),
    .Y(_05310_));
 AO21x1_ASAP7_75t_R _27738_ (.A1(_05309_),
    .A2(_05310_),
    .B(net6069),
    .Y(_05311_));
 AO21x1_ASAP7_75t_R _27739_ (.A1(net6083),
    .A2(net6084),
    .B(_05233_),
    .Y(_05312_));
 AOI21x1_ASAP7_75t_R _27740_ (.A1(net6081),
    .A2(_05312_),
    .B(net6062),
    .Y(_05313_));
 AO21x1_ASAP7_75t_R _27741_ (.A1(_05196_),
    .A2(_05260_),
    .B(net6081),
    .Y(_05314_));
 AOI21x1_ASAP7_75t_R _27743_ (.A1(_05313_),
    .A2(_05314_),
    .B(net5366),
    .Y(_05316_));
 OAI21x1_ASAP7_75t_R _27744_ (.A1(_05307_),
    .A2(_05311_),
    .B(_05316_),
    .Y(_05317_));
 NOR2x1_ASAP7_75t_R _27745_ (.A(net6061),
    .B(_05151_),
    .Y(_05318_));
 NOR2x1_ASAP7_75t_R _27746_ (.A(net4800),
    .B(net5636),
    .Y(_05319_));
 AO21x1_ASAP7_75t_R _27747_ (.A1(net6083),
    .A2(net6084),
    .B(_01328_),
    .Y(_05320_));
 INVx1_ASAP7_75t_R _27748_ (.A(_05320_),
    .Y(_05321_));
 OAI21x1_ASAP7_75t_R _27749_ (.A1(net4628),
    .A2(_05321_),
    .B(net6072),
    .Y(_05322_));
 AOI21x1_ASAP7_75t_R _27750_ (.A1(_05318_),
    .A2(_05322_),
    .B(net5632),
    .Y(_05323_));
 AO21x1_ASAP7_75t_R _27751_ (.A1(net6085),
    .A2(net6086),
    .B(_01330_),
    .Y(_05324_));
 NOR2x1_ASAP7_75t_R _27752_ (.A(net6081),
    .B(_05324_),
    .Y(_05325_));
 NOR2x1_ASAP7_75t_R _27753_ (.A(net6069),
    .B(_05325_),
    .Y(_05326_));
 OAI21x1_ASAP7_75t_R _27754_ (.A1(_05247_),
    .A2(_05249_),
    .B(_05326_),
    .Y(_05327_));
 AOI21x1_ASAP7_75t_R _27756_ (.A1(_05327_),
    .A2(_05323_),
    .B(net6060),
    .Y(_05329_));
 AOI21x1_ASAP7_75t_R _27757_ (.A1(_05329_),
    .A2(_05317_),
    .B(net6059),
    .Y(_05330_));
 OAI21x1_ASAP7_75t_R _27758_ (.A1(_05291_),
    .A2(_05304_),
    .B(_05330_),
    .Y(_05331_));
 OAI21x1_ASAP7_75t_R _27759_ (.A1(_05221_),
    .A2(_05278_),
    .B(_05331_),
    .Y(_00128_));
 NAND2x1_ASAP7_75t_R _27760_ (.A(_05305_),
    .B(_05203_),
    .Y(_05332_));
 NOR2x1_ASAP7_75t_R _27761_ (.A(net5636),
    .B(_05147_),
    .Y(_05333_));
 NAND2x1_ASAP7_75t_R _27762_ (.A(_05333_),
    .B(net4846),
    .Y(_05334_));
 AND3x1_ASAP7_75t_R _27763_ (.A(_05332_),
    .B(net6065),
    .C(_05334_),
    .Y(_05335_));
 AO21x1_ASAP7_75t_R _27764_ (.A1(net6083),
    .A2(net6084),
    .B(net4800),
    .Y(_05336_));
 NAND2x1_ASAP7_75t_R _27765_ (.A(net5638),
    .B(net5095),
    .Y(_05337_));
 AOI21x1_ASAP7_75t_R _27766_ (.A1(net4624),
    .A2(_05337_),
    .B(net6078),
    .Y(_05338_));
 INVx3_ASAP7_75t_R _27767_ (.A(_05150_),
    .Y(_05339_));
 AO21x1_ASAP7_75t_R _27768_ (.A1(_05244_),
    .A2(_05339_),
    .B(net6062),
    .Y(_05340_));
 OAI21x1_ASAP7_75t_R _27769_ (.A1(_05338_),
    .A2(_05340_),
    .B(net5634),
    .Y(_05341_));
 NOR2x1_ASAP7_75t_R _27770_ (.A(_05335_),
    .B(_05341_),
    .Y(_05342_));
 AO21x1_ASAP7_75t_R _27771_ (.A1(_05319_),
    .A2(net6075),
    .B(net6065),
    .Y(_05343_));
 INVx1_ASAP7_75t_R _27772_ (.A(_05242_),
    .Y(_05344_));
 AOI21x1_ASAP7_75t_R _27773_ (.A1(net5638),
    .A2(net5641),
    .B(net6074),
    .Y(_05345_));
 INVx1_ASAP7_75t_R _27774_ (.A(_05345_),
    .Y(_05346_));
 NAND2x1_ASAP7_75t_R _27775_ (.A(net5094),
    .B(_05346_),
    .Y(_05347_));
 OAI21x1_ASAP7_75t_R _27776_ (.A1(net4495),
    .A2(_05347_),
    .B(net5367),
    .Y(_05348_));
 AOI21x1_ASAP7_75t_R _27777_ (.A1(net4721),
    .A2(net5639),
    .B(net6073),
    .Y(_05349_));
 AO21x1_ASAP7_75t_R _27778_ (.A1(_05349_),
    .A2(net4496),
    .B(net6069),
    .Y(_05350_));
 AO21x1_ASAP7_75t_R _27780_ (.A1(net6075),
    .A2(_05289_),
    .B(_05325_),
    .Y(_05352_));
 NOR2x1_ASAP7_75t_R _27781_ (.A(_05350_),
    .B(_05352_),
    .Y(_05353_));
 OAI21x1_ASAP7_75t_R _27782_ (.A1(_05348_),
    .A2(_05353_),
    .B(net6060),
    .Y(_05354_));
 INVx1_ASAP7_75t_R _27783_ (.A(_05276_),
    .Y(_05355_));
 OAI21x1_ASAP7_75t_R _27784_ (.A1(_05342_),
    .A2(_05354_),
    .B(_05355_),
    .Y(_05356_));
 OAI21x1_ASAP7_75t_R _27786_ (.A1(net5095),
    .A2(net5375),
    .B(net6080),
    .Y(_05358_));
 INVx2_ASAP7_75t_R _27787_ (.A(_05162_),
    .Y(_05359_));
 OA21x2_ASAP7_75t_R _27788_ (.A1(_05336_),
    .A2(net6080),
    .B(net6065),
    .Y(_05360_));
 OA21x2_ASAP7_75t_R _27789_ (.A1(_05358_),
    .A2(net4457),
    .B(_05360_),
    .Y(_05361_));
 OAI21x1_ASAP7_75t_R _27790_ (.A1(net5372),
    .A2(_05224_),
    .B(net6070),
    .Y(_05362_));
 AOI21x1_ASAP7_75t_R _27791_ (.A1(net5640),
    .A2(net5097),
    .B(net5638),
    .Y(_05363_));
 INVx1_ASAP7_75t_R _27792_ (.A(_05363_),
    .Y(_05364_));
 NOR2x1_ASAP7_75t_R _27793_ (.A(net6080),
    .B(_05364_),
    .Y(_05365_));
 OAI21x1_ASAP7_75t_R _27794_ (.A1(net4425),
    .A2(_05365_),
    .B(net5634),
    .Y(_05366_));
 OAI21x1_ASAP7_75t_R _27795_ (.A1(_05361_),
    .A2(_05366_),
    .B(net5631),
    .Y(_05367_));
 OA21x2_ASAP7_75t_R _27796_ (.A1(net5641),
    .A2(net5095),
    .B(_05244_),
    .Y(_05368_));
 AO21x1_ASAP7_75t_R _27797_ (.A1(_05226_),
    .A2(net4543),
    .B(net6070),
    .Y(_05369_));
 OAI21x1_ASAP7_75t_R _27798_ (.A1(_05368_),
    .A2(_05369_),
    .B(net5367),
    .Y(_05370_));
 NOR2x1_ASAP7_75t_R _27799_ (.A(_05195_),
    .B(net5639),
    .Y(_05371_));
 INVx1_ASAP7_75t_R _27800_ (.A(_05371_),
    .Y(_05372_));
 NAND2x1_ASAP7_75t_R _27801_ (.A(_05372_),
    .B(net4847),
    .Y(_05373_));
 OA21x2_ASAP7_75t_R _27802_ (.A1(_05319_),
    .A2(net4458),
    .B(net6079),
    .Y(_05374_));
 AOI211x1_ASAP7_75t_R _27804_ (.A1(_05373_),
    .A2(net6074),
    .B(_05374_),
    .C(net6067),
    .Y(_05376_));
 NOR2x1_ASAP7_75t_R _27805_ (.A(_05370_),
    .B(_05376_),
    .Y(_05377_));
 NOR2x1_ASAP7_75t_R _27806_ (.A(_05367_),
    .B(_05377_),
    .Y(_05378_));
 NOR2x1_ASAP7_75t_R _27807_ (.A(_05119_),
    .B(net5096),
    .Y(_05379_));
 NAND2x1_ASAP7_75t_R _27808_ (.A(net5641),
    .B(_05379_),
    .Y(_05380_));
 NOR2x1_ASAP7_75t_R _27809_ (.A(net6072),
    .B(net5635),
    .Y(_05381_));
 AOI22x1_ASAP7_75t_R _27810_ (.A1(net4623),
    .A2(_05142_),
    .B1(_01337_),
    .B2(_05381_),
    .Y(_05382_));
 OAI21x1_ASAP7_75t_R _27811_ (.A1(net6070),
    .A2(_05382_),
    .B(net6060),
    .Y(_05383_));
 AOI21x1_ASAP7_75t_R _27812_ (.A1(_05146_),
    .A2(_05226_),
    .B(net5367),
    .Y(_05384_));
 AOI21x1_ASAP7_75t_R _27813_ (.A1(net5640),
    .A2(net5095),
    .B(net5636),
    .Y(_05385_));
 OAI21x1_ASAP7_75t_R _27814_ (.A1(net4844),
    .A2(_05385_),
    .B(net6079),
    .Y(_05386_));
 AO21x1_ASAP7_75t_R _27815_ (.A1(net5641),
    .A2(net5638),
    .B(net6077),
    .Y(_05387_));
 NOR2x1_ASAP7_75t_R _27816_ (.A(net4842),
    .B(_05387_),
    .Y(_05388_));
 NAND2x1_ASAP7_75t_R _27817_ (.A(net6078),
    .B(_05312_),
    .Y(_05389_));
 OAI21x1_ASAP7_75t_R _27818_ (.A1(net5368),
    .A2(_05389_),
    .B(net5367),
    .Y(_05390_));
 OAI21x1_ASAP7_75t_R _27819_ (.A1(_05388_),
    .A2(_05390_),
    .B(net6071),
    .Y(_05391_));
 AOI21x1_ASAP7_75t_R _27820_ (.A1(_05384_),
    .A2(_05386_),
    .B(_05391_),
    .Y(_05392_));
 OAI21x1_ASAP7_75t_R _27821_ (.A1(_05383_),
    .A2(_05392_),
    .B(net6059),
    .Y(_05393_));
 AO21x1_ASAP7_75t_R _27822_ (.A1(net6080),
    .A2(net4431),
    .B(net6070),
    .Y(_05394_));
 NOR2x1_ASAP7_75t_R _27823_ (.A(_05231_),
    .B(_05249_),
    .Y(_05395_));
 OAI21x1_ASAP7_75t_R _27824_ (.A1(_05395_),
    .A2(_05394_),
    .B(net5367),
    .Y(_05396_));
 NOR2x1_ASAP7_75t_R _27825_ (.A(net4457),
    .B(_05358_),
    .Y(_05397_));
 OA21x2_ASAP7_75t_R _27826_ (.A1(net5638),
    .A2(net4630),
    .B(net6073),
    .Y(_05398_));
 AO21x1_ASAP7_75t_R _27827_ (.A1(net6085),
    .A2(net6086),
    .B(_05259_),
    .Y(_05399_));
 AO21x1_ASAP7_75t_R _27828_ (.A1(_05398_),
    .A2(_05399_),
    .B(net6065),
    .Y(_05400_));
 NOR2x1_ASAP7_75t_R _27829_ (.A(_05397_),
    .B(_05400_),
    .Y(_05401_));
 OAI21x1_ASAP7_75t_R _27830_ (.A1(_05401_),
    .A2(_05396_),
    .B(net5631),
    .Y(_05402_));
 NOR2x1_ASAP7_75t_R _27831_ (.A(net5637),
    .B(net5095),
    .Y(_05403_));
 AOI21x1_ASAP7_75t_R _27832_ (.A1(net6074),
    .A2(_05403_),
    .B(net6067),
    .Y(_05404_));
 NAND2x1_ASAP7_75t_R _27833_ (.A(_05130_),
    .B(_05349_),
    .Y(_05405_));
 AND3x1_ASAP7_75t_R _27834_ (.A(_05404_),
    .B(_05302_),
    .C(_05405_),
    .Y(_05406_));
 AND2x2_ASAP7_75t_R _27835_ (.A(_05204_),
    .B(_05146_),
    .Y(_05407_));
 INVx1_ASAP7_75t_R _27836_ (.A(_05262_),
    .Y(_05408_));
 AO21x1_ASAP7_75t_R _27837_ (.A1(_05234_),
    .A2(_05408_),
    .B(net6071),
    .Y(_05409_));
 OAI21x1_ASAP7_75t_R _27838_ (.A1(_05407_),
    .A2(_05409_),
    .B(net5634),
    .Y(_05410_));
 NOR2x1_ASAP7_75t_R _27839_ (.A(_05406_),
    .B(_05410_),
    .Y(_05411_));
 NOR2x1_ASAP7_75t_R _27840_ (.A(_05411_),
    .B(_05402_),
    .Y(_05412_));
 OAI22x1_ASAP7_75t_R _27841_ (.A1(_05356_),
    .A2(_05378_),
    .B1(_05412_),
    .B2(_05393_),
    .Y(_00129_));
 NAND2x1_ASAP7_75t_R _27842_ (.A(net6061),
    .B(_05322_),
    .Y(_05413_));
 INVx1_ASAP7_75t_R _27843_ (.A(net5371),
    .Y(_05414_));
 OA21x2_ASAP7_75t_R _27844_ (.A1(_05414_),
    .A2(net4628),
    .B(net6081),
    .Y(_05415_));
 OA21x2_ASAP7_75t_R _27845_ (.A1(_05413_),
    .A2(_05415_),
    .B(net5366),
    .Y(_05416_));
 NAND2x1_ASAP7_75t_R _27846_ (.A(_05140_),
    .B(_05324_),
    .Y(_05417_));
 NOR2x1_ASAP7_75t_R _27847_ (.A(net4843),
    .B(_05417_),
    .Y(_05418_));
 AO21x1_ASAP7_75t_R _27848_ (.A1(net6085),
    .A2(net6086),
    .B(net4799),
    .Y(_05419_));
 AND3x1_ASAP7_75t_R _27850_ (.A(net4626),
    .B(net4621),
    .C(net6072),
    .Y(_05421_));
 OAI21x1_ASAP7_75t_R _27851_ (.A1(_05418_),
    .A2(_05421_),
    .B(net6068),
    .Y(_05422_));
 OA21x2_ASAP7_75t_R _27852_ (.A1(net5640),
    .A2(net5636),
    .B(net6082),
    .Y(_05423_));
 INVx1_ASAP7_75t_R _27853_ (.A(_05423_),
    .Y(_05424_));
 AOI21x1_ASAP7_75t_R _27854_ (.A1(net4622),
    .A2(_05204_),
    .B(net6065),
    .Y(_05425_));
 OAI21x1_ASAP7_75t_R _27855_ (.A1(_05321_),
    .A2(_05424_),
    .B(_05425_),
    .Y(_05426_));
 AO21x1_ASAP7_75t_R _27856_ (.A1(net6085),
    .A2(net6086),
    .B(net4546),
    .Y(_05427_));
 AO21x1_ASAP7_75t_R _27857_ (.A1(_05427_),
    .A2(_05162_),
    .B(net6075),
    .Y(_05428_));
 AOI21x1_ASAP7_75t_R _27858_ (.A1(net4801),
    .A2(net5639),
    .B(_05140_),
    .Y(_05429_));
 NAND2x1_ASAP7_75t_R _27859_ (.A(_05310_),
    .B(net4619),
    .Y(_05430_));
 AO21x1_ASAP7_75t_R _27860_ (.A1(_05428_),
    .A2(_05430_),
    .B(net6069),
    .Y(_05431_));
 AOI21x1_ASAP7_75t_R _27861_ (.A1(_05426_),
    .A2(_05431_),
    .B(net5366),
    .Y(_05432_));
 AOI211x1_ASAP7_75t_R _27862_ (.A1(_05416_),
    .A2(_05422_),
    .B(_05432_),
    .C(net6060),
    .Y(_05433_));
 OAI21x1_ASAP7_75t_R _27863_ (.A1(net5637),
    .A2(net5095),
    .B(net5641),
    .Y(_05434_));
 NAND2x1_ASAP7_75t_R _27864_ (.A(net6077),
    .B(_05434_),
    .Y(_05435_));
 AO21x1_ASAP7_75t_R _27865_ (.A1(net4621),
    .A2(_05336_),
    .B(net6081),
    .Y(_05436_));
 AO21x1_ASAP7_75t_R _27866_ (.A1(_05435_),
    .A2(_05436_),
    .B(net6061),
    .Y(_05437_));
 OA21x2_ASAP7_75t_R _27867_ (.A1(_05417_),
    .A2(_05289_),
    .B(net6061),
    .Y(_05438_));
 NAND2x1_ASAP7_75t_R _27868_ (.A(_05306_),
    .B(_05438_),
    .Y(_05439_));
 AOI21x1_ASAP7_75t_R _27869_ (.A1(_05437_),
    .A2(_05439_),
    .B(net5632),
    .Y(_05440_));
 NAND2x1_ASAP7_75t_R _27870_ (.A(net6066),
    .B(_05241_),
    .Y(_05441_));
 AO21x1_ASAP7_75t_R _27871_ (.A1(net6083),
    .A2(net6084),
    .B(net4799),
    .Y(_05442_));
 AOI21x1_ASAP7_75t_R _27872_ (.A1(_05442_),
    .A2(_05190_),
    .B(net6073),
    .Y(_05443_));
 OAI21x1_ASAP7_75t_R _27873_ (.A1(_05441_),
    .A2(_05443_),
    .B(net5635),
    .Y(_05444_));
 AO21x1_ASAP7_75t_R _27874_ (.A1(net5377),
    .A2(_05339_),
    .B(net6076),
    .Y(_05445_));
 NOR2x1_ASAP7_75t_R _27875_ (.A(net4803),
    .B(net5637),
    .Y(_05446_));
 OR3x1_ASAP7_75t_R _27876_ (.A(net4841),
    .B(net6073),
    .C(_05446_),
    .Y(_05447_));
 AOI21x1_ASAP7_75t_R _27877_ (.A1(_05447_),
    .A2(_05445_),
    .B(net6066),
    .Y(_05448_));
 OAI21x1_ASAP7_75t_R _27878_ (.A1(_05444_),
    .A2(_05448_),
    .B(net6060),
    .Y(_05449_));
 OAI21x1_ASAP7_75t_R _27879_ (.A1(_05440_),
    .A2(_05449_),
    .B(net6059),
    .Y(_05450_));
 AO21x1_ASAP7_75t_R _27880_ (.A1(net6083),
    .A2(net6084),
    .B(_05287_),
    .Y(_05451_));
 AOI21x1_ASAP7_75t_R _27881_ (.A1(net4494),
    .A2(_05190_),
    .B(net6073),
    .Y(_05452_));
 OAI21x1_ASAP7_75t_R _27882_ (.A1(net5095),
    .A2(net5370),
    .B(_05142_),
    .Y(_05453_));
 NAND2x1_ASAP7_75t_R _27883_ (.A(net6068),
    .B(_05453_),
    .Y(_05454_));
 AOI21x1_ASAP7_75t_R _27884_ (.A1(net6073),
    .A2(_05371_),
    .B(net6068),
    .Y(_05455_));
 AO21x1_ASAP7_75t_R _27885_ (.A1(net4625),
    .A2(net4544),
    .B(net6073),
    .Y(_05456_));
 AOI21x1_ASAP7_75t_R _27886_ (.A1(_05455_),
    .A2(_05456_),
    .B(net5367),
    .Y(_05457_));
 OAI21x1_ASAP7_75t_R _27887_ (.A1(_05452_),
    .A2(_05454_),
    .B(_05457_),
    .Y(_05458_));
 NAND2x1_ASAP7_75t_R _27888_ (.A(_01339_),
    .B(net6076),
    .Y(_05459_));
 NAND2x1_ASAP7_75t_R _27889_ (.A(_05459_),
    .B(_05241_),
    .Y(_05460_));
 OA21x2_ASAP7_75t_R _27890_ (.A1(_01341_),
    .A2(net6077),
    .B(net6068),
    .Y(_05461_));
 AOI21x1_ASAP7_75t_R _27892_ (.A1(_05461_),
    .A2(_05435_),
    .B(net5635),
    .Y(_05463_));
 OAI21x1_ASAP7_75t_R _27893_ (.A1(net6068),
    .A2(_05460_),
    .B(_05463_),
    .Y(_05464_));
 AOI21x1_ASAP7_75t_R _27894_ (.A1(_05458_),
    .A2(_05464_),
    .B(_05237_),
    .Y(_05465_));
 OA21x2_ASAP7_75t_R _27895_ (.A1(_01340_),
    .A2(_05140_),
    .B(net6065),
    .Y(_05466_));
 OAI21x1_ASAP7_75t_R _27896_ (.A1(net5099),
    .A2(net5369),
    .B(_05349_),
    .Y(_05467_));
 AOI21x1_ASAP7_75t_R _27897_ (.A1(_05466_),
    .A2(_05467_),
    .B(net5366),
    .Y(_05468_));
 AOI21x1_ASAP7_75t_R _27898_ (.A1(net4543),
    .A2(net5365),
    .B(net6061),
    .Y(_05469_));
 NAND2x1_ASAP7_75t_R _27899_ (.A(_05310_),
    .B(_05423_),
    .Y(_05470_));
 NAND2x1_ASAP7_75t_R _27900_ (.A(_05469_),
    .B(_05470_),
    .Y(_05471_));
 NAND2x1_ASAP7_75t_R _27901_ (.A(_05468_),
    .B(_05471_),
    .Y(_05472_));
 AOI21x1_ASAP7_75t_R _27902_ (.A1(net5636),
    .A2(net5640),
    .B(net6072),
    .Y(_05473_));
 AND2x2_ASAP7_75t_R _27903_ (.A(net6072),
    .B(_01337_),
    .Y(_05474_));
 AOI21x1_ASAP7_75t_R _27904_ (.A1(_05473_),
    .A2(net4848),
    .B(_05474_),
    .Y(_05475_));
 AOI21x1_ASAP7_75t_R _27905_ (.A1(net6064),
    .A2(_05475_),
    .B(net5635),
    .Y(_05476_));
 INVx1_ASAP7_75t_R _27906_ (.A(net4543),
    .Y(_05477_));
 NAND2x1_ASAP7_75t_R _27907_ (.A(net6077),
    .B(_05197_),
    .Y(_05478_));
 NOR2x1_ASAP7_75t_R _27908_ (.A(_05477_),
    .B(_05478_),
    .Y(_05479_));
 AND2x2_ASAP7_75t_R _27909_ (.A(_05305_),
    .B(_05196_),
    .Y(_05480_));
 OAI21x1_ASAP7_75t_R _27910_ (.A1(_05479_),
    .A2(_05480_),
    .B(net6068),
    .Y(_05481_));
 NAND2x1_ASAP7_75t_R _27911_ (.A(_05476_),
    .B(_05481_),
    .Y(_05482_));
 AOI21x1_ASAP7_75t_R _27912_ (.A1(_05472_),
    .A2(_05482_),
    .B(net6060),
    .Y(_05483_));
 OAI21x1_ASAP7_75t_R _27913_ (.A1(_05465_),
    .A2(_05483_),
    .B(_05355_),
    .Y(_05484_));
 OAI21x1_ASAP7_75t_R _27914_ (.A1(_05433_),
    .A2(_05450_),
    .B(_05484_),
    .Y(_00130_));
 AOI21x1_ASAP7_75t_R _27915_ (.A1(net4625),
    .A2(_05442_),
    .B(net6073),
    .Y(_05485_));
 NAND2x1_ASAP7_75t_R _27916_ (.A(net5635),
    .B(_05445_),
    .Y(_05486_));
 NAND2x1_ASAP7_75t_R _27917_ (.A(_05151_),
    .B(_05408_),
    .Y(_05487_));
 AOI21x1_ASAP7_75t_R _27918_ (.A1(net4845),
    .A2(_05204_),
    .B(net5635),
    .Y(_05488_));
 AOI21x1_ASAP7_75t_R _27919_ (.A1(_05487_),
    .A2(_05488_),
    .B(net6068),
    .Y(_05489_));
 OAI21x1_ASAP7_75t_R _27920_ (.A1(_05485_),
    .A2(_05486_),
    .B(_05489_),
    .Y(_05490_));
 AO21x1_ASAP7_75t_R _27921_ (.A1(_05349_),
    .A2(_05372_),
    .B(net5367),
    .Y(_05491_));
 AOI211x1_ASAP7_75t_R _27922_ (.A1(net4802),
    .A2(net5637),
    .B(net4840),
    .C(net6076),
    .Y(_05492_));
 AOI21x1_ASAP7_75t_R _27923_ (.A1(net6076),
    .A2(_05168_),
    .B(net5635),
    .Y(_05493_));
 OAI21x1_ASAP7_75t_R _27924_ (.A1(net4841),
    .A2(_05387_),
    .B(_05493_),
    .Y(_05494_));
 OAI21x1_ASAP7_75t_R _27925_ (.A1(_05491_),
    .A2(_05492_),
    .B(_05494_),
    .Y(_05495_));
 AOI21x1_ASAP7_75t_R _27926_ (.A1(net6068),
    .A2(_05495_),
    .B(_05237_),
    .Y(_05496_));
 NAND2x1_ASAP7_75t_R _27927_ (.A(_05490_),
    .B(_05496_),
    .Y(_05497_));
 NOR2x1_ASAP7_75t_R _27928_ (.A(_05385_),
    .B(_05478_),
    .Y(_05498_));
 OAI21x1_ASAP7_75t_R _27929_ (.A1(net4844),
    .A2(_05283_),
    .B(net6065),
    .Y(_05499_));
 NOR2x1_ASAP7_75t_R _27930_ (.A(_05498_),
    .B(_05499_),
    .Y(_05500_));
 AO21x1_ASAP7_75t_R _27931_ (.A1(net6085),
    .A2(net6086),
    .B(_05132_),
    .Y(_05501_));
 AO21x1_ASAP7_75t_R _27932_ (.A1(_05501_),
    .A2(_05339_),
    .B(net6076),
    .Y(_05502_));
 NOR2x1_ASAP7_75t_R _27933_ (.A(net5097),
    .B(net5373),
    .Y(_05503_));
 OAI21x1_ASAP7_75t_R _27934_ (.A1(net4840),
    .A2(_05503_),
    .B(net6076),
    .Y(_05504_));
 AOI21x1_ASAP7_75t_R _27935_ (.A1(_05502_),
    .A2(_05504_),
    .B(net6066),
    .Y(_05505_));
 OAI21x1_ASAP7_75t_R _27936_ (.A1(_05500_),
    .A2(_05505_),
    .B(net5633),
    .Y(_05506_));
 NAND2x1_ASAP7_75t_R _27937_ (.A(net4847),
    .B(_05203_),
    .Y(_05507_));
 AO21x1_ASAP7_75t_R _27938_ (.A1(net5637),
    .A2(net6076),
    .B(net6068),
    .Y(_05508_));
 OA21x2_ASAP7_75t_R _27939_ (.A1(_05507_),
    .A2(_05508_),
    .B(net5367),
    .Y(_05509_));
 NAND2x1_ASAP7_75t_R _27940_ (.A(net4545),
    .B(net4620),
    .Y(_05510_));
 INVx1_ASAP7_75t_R _27941_ (.A(_05362_),
    .Y(_05511_));
 NAND2x1_ASAP7_75t_R _27942_ (.A(_05510_),
    .B(_05511_),
    .Y(_05512_));
 AOI21x1_ASAP7_75t_R _27943_ (.A1(_05509_),
    .A2(_05512_),
    .B(net6060),
    .Y(_05513_));
 AOI21x1_ASAP7_75t_R _27944_ (.A1(_05506_),
    .A2(_05513_),
    .B(net6059),
    .Y(_05514_));
 NAND2x1_ASAP7_75t_R _27945_ (.A(_05497_),
    .B(_05514_),
    .Y(_05515_));
 NOR2x1_ASAP7_75t_R _27946_ (.A(net6072),
    .B(_05320_),
    .Y(_05516_));
 NOR2x1_ASAP7_75t_R _27947_ (.A(net5366),
    .B(_05516_),
    .Y(_05517_));
 NAND2x1_ASAP7_75t_R _27948_ (.A(_05430_),
    .B(_05517_),
    .Y(_05518_));
 AND3x1_ASAP7_75t_R _27949_ (.A(net6085),
    .B(net6086),
    .C(_05287_),
    .Y(_05519_));
 AOI21x1_ASAP7_75t_R _27950_ (.A1(_05339_),
    .A2(_05230_),
    .B(net5634),
    .Y(_05520_));
 OAI21x1_ASAP7_75t_R _27951_ (.A1(net4439),
    .A2(net4493),
    .B(_05520_),
    .Y(_05521_));
 NAND2x1_ASAP7_75t_R _27952_ (.A(_05518_),
    .B(_05521_),
    .Y(_05522_));
 NAND2x1p5_ASAP7_75t_R _27953_ (.A(net6074),
    .B(net4458),
    .Y(_05523_));
 OAI21x1_ASAP7_75t_R _27954_ (.A1(net5367),
    .A2(_05523_),
    .B(_05293_),
    .Y(_05524_));
 NAND2x1_ASAP7_75t_R _27955_ (.A(net5370),
    .B(_05142_),
    .Y(_05525_));
 AOI21x1_ASAP7_75t_R _27956_ (.A1(_05169_),
    .A2(_05525_),
    .B(net5632),
    .Y(_05526_));
 OAI21x1_ASAP7_75t_R _27957_ (.A1(_05524_),
    .A2(_05526_),
    .B(net6060),
    .Y(_05527_));
 AOI21x1_ASAP7_75t_R _27958_ (.A1(net6065),
    .A2(_05522_),
    .B(_05527_),
    .Y(_05528_));
 AO21x1_ASAP7_75t_R _27959_ (.A1(net6085),
    .A2(net6086),
    .B(net4801),
    .Y(_05529_));
 AO21x1_ASAP7_75t_R _27960_ (.A1(_05529_),
    .A2(_05451_),
    .B(net6073),
    .Y(_05530_));
 AOI21x1_ASAP7_75t_R _27961_ (.A1(_05453_),
    .A2(_05530_),
    .B(net6068),
    .Y(_05531_));
 OAI21x1_ASAP7_75t_R _27962_ (.A1(_05425_),
    .A2(_05531_),
    .B(net5367),
    .Y(_05532_));
 AOI21x1_ASAP7_75t_R _27963_ (.A1(_05332_),
    .A2(_05286_),
    .B(net5367),
    .Y(_05533_));
 OA21x2_ASAP7_75t_R _27964_ (.A1(net4627),
    .A2(net6075),
    .B(net6068),
    .Y(_05534_));
 AO21x1_ASAP7_75t_R _27965_ (.A1(_05162_),
    .A2(net4622),
    .B(net6078),
    .Y(_05535_));
 NAND2x1_ASAP7_75t_R _27966_ (.A(net5095),
    .B(_05333_),
    .Y(_05536_));
 NAND3x1_ASAP7_75t_R _27967_ (.A(_05534_),
    .B(_05535_),
    .C(_05536_),
    .Y(_05537_));
 NAND2x1_ASAP7_75t_R _27968_ (.A(_05533_),
    .B(_05537_),
    .Y(_05538_));
 AOI21x1_ASAP7_75t_R _27969_ (.A1(_05532_),
    .A2(_05538_),
    .B(net6060),
    .Y(_05539_));
 OAI21x1_ASAP7_75t_R _27970_ (.A1(_05528_),
    .A2(_05539_),
    .B(net6059),
    .Y(_05540_));
 NAND2x1_ASAP7_75t_R _27971_ (.A(_05515_),
    .B(_05540_),
    .Y(_00131_));
 AO21x1_ASAP7_75t_R _27972_ (.A1(net4543),
    .A2(net4626),
    .B(net6072),
    .Y(_05541_));
 AO21x1_ASAP7_75t_R _27973_ (.A1(_05541_),
    .A2(_05322_),
    .B(net6061),
    .Y(_05542_));
 AND3x1_ASAP7_75t_R _27974_ (.A(net4456),
    .B(_05243_),
    .C(net6075),
    .Y(_05543_));
 NOR2x1_ASAP7_75t_R _27975_ (.A(_05301_),
    .B(_05296_),
    .Y(_05544_));
 OAI21x1_ASAP7_75t_R _27976_ (.A1(_05543_),
    .A2(_05544_),
    .B(net6061),
    .Y(_05545_));
 AOI21x1_ASAP7_75t_R _27977_ (.A1(_05542_),
    .A2(_05545_),
    .B(net5366),
    .Y(_05546_));
 AO21x1_ASAP7_75t_R _27978_ (.A1(_05423_),
    .A2(_05130_),
    .B(net6069),
    .Y(_05547_));
 NOR2x1_ASAP7_75t_R _27979_ (.A(_05352_),
    .B(_05547_),
    .Y(_05548_));
 OAI21x1_ASAP7_75t_R _27980_ (.A1(_05296_),
    .A2(_05424_),
    .B(_05436_),
    .Y(_05549_));
 OAI21x1_ASAP7_75t_R _27981_ (.A1(net6061),
    .A2(_05549_),
    .B(net5366),
    .Y(_05550_));
 OAI21x1_ASAP7_75t_R _27982_ (.A1(_05548_),
    .A2(_05550_),
    .B(_05355_),
    .Y(_05551_));
 OAI21x1_ASAP7_75t_R _27983_ (.A1(_05546_),
    .A2(_05551_),
    .B(net6060),
    .Y(_05552_));
 NAND2x1_ASAP7_75t_R _27984_ (.A(net6075),
    .B(_05289_),
    .Y(_05553_));
 NAND2x1_ASAP7_75t_R _27985_ (.A(_05300_),
    .B(net5094),
    .Y(_05554_));
 AO21x1_ASAP7_75t_R _27986_ (.A1(_05553_),
    .A2(_05554_),
    .B(net6062),
    .Y(_05555_));
 INVx1_ASAP7_75t_R _27987_ (.A(_01331_),
    .Y(_05556_));
 AO221x1_ASAP7_75t_R _27988_ (.A1(_05556_),
    .A2(net6074),
    .B1(net4546),
    .B2(_05333_),
    .C(net6071),
    .Y(_05557_));
 AOI21x1_ASAP7_75t_R _27989_ (.A1(_05555_),
    .A2(_05557_),
    .B(net5366),
    .Y(_05558_));
 NOR2x1_ASAP7_75t_R _27990_ (.A(net4843),
    .B(_05301_),
    .Y(_05559_));
 NAND2x1_ASAP7_75t_R _27991_ (.A(net5640),
    .B(net5099),
    .Y(_05560_));
 AOI21x1_ASAP7_75t_R _27992_ (.A1(_05560_),
    .A2(net5094),
    .B(net6081),
    .Y(_05561_));
 OAI21x1_ASAP7_75t_R _27993_ (.A1(_05559_),
    .A2(_05561_),
    .B(net6069),
    .Y(_05562_));
 AO21x1_ASAP7_75t_R _27994_ (.A1(_05210_),
    .A2(_05314_),
    .B(net6069),
    .Y(_05563_));
 AOI21x1_ASAP7_75t_R _27995_ (.A1(_05562_),
    .A2(_05563_),
    .B(net5632),
    .Y(_05564_));
 NOR3x1_ASAP7_75t_R _27996_ (.A(_05558_),
    .B(_05564_),
    .C(_05355_),
    .Y(_05565_));
 AO21x1_ASAP7_75t_R _27997_ (.A1(_05203_),
    .A2(_05473_),
    .B(net6069),
    .Y(_05566_));
 OAI21x1_ASAP7_75t_R _27998_ (.A1(_05388_),
    .A2(_05566_),
    .B(net5367),
    .Y(_05567_));
 AND2x2_ASAP7_75t_R _27999_ (.A(_05473_),
    .B(_05196_),
    .Y(_05568_));
 OA21x2_ASAP7_75t_R _28000_ (.A1(_05568_),
    .A2(_05561_),
    .B(net6070),
    .Y(_05569_));
 NAND2x1_ASAP7_75t_R _28001_ (.A(_05260_),
    .B(net6069),
    .Y(_05570_));
 OA21x2_ASAP7_75t_R _28002_ (.A1(_05570_),
    .A2(_05300_),
    .B(net5632),
    .Y(_05571_));
 NAND2x1_ASAP7_75t_R _28003_ (.A(_05310_),
    .B(_05345_),
    .Y(_05572_));
 AOI21x1_ASAP7_75t_R _28004_ (.A1(_05146_),
    .A2(_05226_),
    .B(net6070),
    .Y(_05573_));
 NAND2x1_ASAP7_75t_R _28005_ (.A(_05572_),
    .B(_05573_),
    .Y(_05574_));
 AOI21x1_ASAP7_75t_R _28006_ (.A1(_05571_),
    .A2(_05574_),
    .B(net6059),
    .Y(_05575_));
 OAI21x1_ASAP7_75t_R _28007_ (.A1(_05567_),
    .A2(_05569_),
    .B(_05575_),
    .Y(_05576_));
 NOR2x1_ASAP7_75t_R _28008_ (.A(net6071),
    .B(_05333_),
    .Y(_05577_));
 NAND2x1_ASAP7_75t_R _28009_ (.A(_05223_),
    .B(_05204_),
    .Y(_05578_));
 AOI21x1_ASAP7_75t_R _28010_ (.A1(_05577_),
    .A2(_05578_),
    .B(net5633),
    .Y(_05579_));
 OAI21x1_ASAP7_75t_R _28011_ (.A1(_05371_),
    .A2(net5368),
    .B(net6073),
    .Y(_05580_));
 AOI21x1_ASAP7_75t_R _28012_ (.A1(_05408_),
    .A2(_05234_),
    .B(_05170_),
    .Y(_05581_));
 NAND2x1_ASAP7_75t_R _28013_ (.A(_05580_),
    .B(_05581_),
    .Y(_05582_));
 AOI21x1_ASAP7_75t_R _28014_ (.A1(_05579_),
    .A2(_05582_),
    .B(_05355_),
    .Y(_05583_));
 NAND2x1_ASAP7_75t_R _28015_ (.A(net6074),
    .B(_05399_),
    .Y(_05584_));
 AND2x2_ASAP7_75t_R _28016_ (.A(_05584_),
    .B(net6071),
    .Y(_05585_));
 AOI21x1_ASAP7_75t_R _28017_ (.A1(_05358_),
    .A2(_05585_),
    .B(net5367),
    .Y(_05586_));
 AO21x1_ASAP7_75t_R _28018_ (.A1(_05427_),
    .A2(_05336_),
    .B(net6079),
    .Y(_05587_));
 AOI21x1_ASAP7_75t_R _28019_ (.A1(_05244_),
    .A2(_05380_),
    .B(net6071),
    .Y(_05588_));
 NAND2x1_ASAP7_75t_R _28020_ (.A(_05587_),
    .B(_05588_),
    .Y(_05589_));
 NAND2x1_ASAP7_75t_R _28021_ (.A(_05586_),
    .B(_05589_),
    .Y(_05590_));
 AOI21x1_ASAP7_75t_R _28022_ (.A1(_05583_),
    .A2(_05590_),
    .B(net6060),
    .Y(_05591_));
 NAND2x1_ASAP7_75t_R _28023_ (.A(_05576_),
    .B(_05591_),
    .Y(_05592_));
 OAI21x1_ASAP7_75t_R _28024_ (.A1(_05552_),
    .A2(_05565_),
    .B(_05592_),
    .Y(_00132_));
 NAND2x1_ASAP7_75t_R _28025_ (.A(_05339_),
    .B(net4622),
    .Y(_05593_));
 AO22x1_ASAP7_75t_R _28026_ (.A1(_05308_),
    .A2(_05151_),
    .B1(_05593_),
    .B2(net6074),
    .Y(_05594_));
 OA21x2_ASAP7_75t_R _28027_ (.A1(_05132_),
    .A2(net6073),
    .B(net6065),
    .Y(_05595_));
 AO21x1_ASAP7_75t_R _28028_ (.A1(net4842),
    .A2(net5641),
    .B(net6077),
    .Y(_05596_));
 AOI21x1_ASAP7_75t_R _28029_ (.A1(_05595_),
    .A2(_05596_),
    .B(net5633),
    .Y(_05597_));
 OAI21x1_ASAP7_75t_R _28030_ (.A1(net6066),
    .A2(_05594_),
    .B(_05597_),
    .Y(_05598_));
 OA21x2_ASAP7_75t_R _28031_ (.A1(_05519_),
    .A2(net6075),
    .B(net6065),
    .Y(_05599_));
 OAI21x1_ASAP7_75t_R _28032_ (.A1(_05249_),
    .A2(_05241_),
    .B(_05599_),
    .Y(_05600_));
 INVx1_ASAP7_75t_R _28033_ (.A(_05224_),
    .Y(_05601_));
 OA21x2_ASAP7_75t_R _28034_ (.A1(_05343_),
    .A2(_05601_),
    .B(net5634),
    .Y(_05602_));
 AOI21x1_ASAP7_75t_R _28035_ (.A1(_05600_),
    .A2(_05602_),
    .B(_05237_),
    .Y(_05603_));
 NAND2x1_ASAP7_75t_R _28036_ (.A(_05598_),
    .B(_05603_),
    .Y(_05604_));
 OAI21x1_ASAP7_75t_R _28037_ (.A1(net5097),
    .A2(net5377),
    .B(_05151_),
    .Y(_05605_));
 AOI21x1_ASAP7_75t_R _28038_ (.A1(net4620),
    .A2(net5094),
    .B(_05170_),
    .Y(_05606_));
 NAND2x1_ASAP7_75t_R _28039_ (.A(_05605_),
    .B(_05606_),
    .Y(_05607_));
 OA21x2_ASAP7_75t_R _28040_ (.A1(net5095),
    .A2(net6074),
    .B(net6065),
    .Y(_05608_));
 AOI21x1_ASAP7_75t_R _28041_ (.A1(_05608_),
    .A2(_05205_),
    .B(net5367),
    .Y(_05609_));
 AOI21x1_ASAP7_75t_R _28042_ (.A1(_05607_),
    .A2(_05609_),
    .B(net6060),
    .Y(_05610_));
 OA21x2_ASAP7_75t_R _28043_ (.A1(_05501_),
    .A2(net6074),
    .B(net6071),
    .Y(_05611_));
 INVx1_ASAP7_75t_R _28044_ (.A(net4622),
    .Y(_05612_));
 OAI21x1_ASAP7_75t_R _28045_ (.A1(_05612_),
    .A2(net4844),
    .B(net6074),
    .Y(_05613_));
 AOI21x1_ASAP7_75t_R _28046_ (.A1(_05611_),
    .A2(_05613_),
    .B(net5635),
    .Y(_05614_));
 NAND2x1_ASAP7_75t_R _28047_ (.A(net5637),
    .B(net5097),
    .Y(_05615_));
 AO21x1_ASAP7_75t_R _28048_ (.A1(_05615_),
    .A2(net4625),
    .B(net6076),
    .Y(_05616_));
 NAND2x1_ASAP7_75t_R _28049_ (.A(_05616_),
    .B(_05588_),
    .Y(_05617_));
 NAND2x1_ASAP7_75t_R _28050_ (.A(_05614_),
    .B(_05617_),
    .Y(_05618_));
 AOI21x1_ASAP7_75t_R _28051_ (.A1(_05610_),
    .A2(_05618_),
    .B(_05355_),
    .Y(_05619_));
 NAND2x1_ASAP7_75t_R _28052_ (.A(_05604_),
    .B(_05619_),
    .Y(_05620_));
 AO21x1_ASAP7_75t_R _28053_ (.A1(net6075),
    .A2(_05339_),
    .B(net6069),
    .Y(_05621_));
 AO21x1_ASAP7_75t_R _28054_ (.A1(_05337_),
    .A2(net4627),
    .B(net6075),
    .Y(_05622_));
 INVx1_ASAP7_75t_R _28055_ (.A(_05622_),
    .Y(_05623_));
 AOI21x1_ASAP7_75t_R _28056_ (.A1(net6075),
    .A2(_05312_),
    .B(net6063),
    .Y(_05624_));
 AOI21x1_ASAP7_75t_R _28057_ (.A1(_05624_),
    .A2(_05334_),
    .B(net5634),
    .Y(_05625_));
 OAI21x1_ASAP7_75t_R _28058_ (.A1(_05621_),
    .A2(_05623_),
    .B(_05625_),
    .Y(_05626_));
 AO21x1_ASAP7_75t_R _28059_ (.A1(_05260_),
    .A2(net4800),
    .B(net6075),
    .Y(_05627_));
 OAI21x1_ASAP7_75t_R _28060_ (.A1(net5099),
    .A2(net5371),
    .B(net4619),
    .Y(_05628_));
 AOI21x1_ASAP7_75t_R _28061_ (.A1(_05627_),
    .A2(_05628_),
    .B(net6062),
    .Y(_05629_));
 AO21x1_ASAP7_75t_R _28062_ (.A1(net4621),
    .A2(_05336_),
    .B(net6075),
    .Y(_05630_));
 AOI21x1_ASAP7_75t_R _28063_ (.A1(_05264_),
    .A2(_05630_),
    .B(net6069),
    .Y(_05631_));
 OAI21x1_ASAP7_75t_R _28064_ (.A1(_05629_),
    .A2(_05631_),
    .B(net5632),
    .Y(_05632_));
 AOI21x1_ASAP7_75t_R _28065_ (.A1(_05626_),
    .A2(_05632_),
    .B(net6060),
    .Y(_05633_));
 AND2x2_ASAP7_75t_R _28066_ (.A(_05501_),
    .B(net6078),
    .Y(_05634_));
 AOI22x1_ASAP7_75t_R _28067_ (.A1(_05634_),
    .A2(_05364_),
    .B1(_05560_),
    .B2(_05230_),
    .Y(_05635_));
 OA21x2_ASAP7_75t_R _28068_ (.A1(net6075),
    .A2(net4543),
    .B(net5367),
    .Y(_05636_));
 OAI21x1_ASAP7_75t_R _28069_ (.A1(_05414_),
    .A2(net4438),
    .B(_05636_),
    .Y(_05637_));
 OAI21x1_ASAP7_75t_R _28070_ (.A1(net5367),
    .A2(_05635_),
    .B(_05637_),
    .Y(_05638_));
 AO21x1_ASAP7_75t_R _28071_ (.A1(net5374),
    .A2(net6081),
    .B(net5367),
    .Y(_05639_));
 NOR2x1_ASAP7_75t_R _28072_ (.A(_05639_),
    .B(_05561_),
    .Y(_05640_));
 AO21x1_ASAP7_75t_R _28073_ (.A1(net4621),
    .A2(net6075),
    .B(net5632),
    .Y(_05641_));
 AND2x2_ASAP7_75t_R _28074_ (.A(_05196_),
    .B(_05151_),
    .Y(_05642_));
 OAI21x1_ASAP7_75t_R _28075_ (.A1(_05641_),
    .A2(_05642_),
    .B(net6061),
    .Y(_05643_));
 OAI21x1_ASAP7_75t_R _28076_ (.A1(_05640_),
    .A2(_05643_),
    .B(net6060),
    .Y(_05644_));
 AOI21x1_ASAP7_75t_R _28077_ (.A1(net6069),
    .A2(_05638_),
    .B(_05644_),
    .Y(_05645_));
 OAI21x1_ASAP7_75t_R _28078_ (.A1(_05633_),
    .A2(_05645_),
    .B(_05355_),
    .Y(_05646_));
 NAND2x1_ASAP7_75t_R _28079_ (.A(_05620_),
    .B(_05646_),
    .Y(_00133_));
 NAND2x1_ASAP7_75t_R _28080_ (.A(net4846),
    .B(_05423_),
    .Y(_05647_));
 AO21x1_ASAP7_75t_R _28081_ (.A1(_01334_),
    .A2(_01338_),
    .B(net6079),
    .Y(_05648_));
 AND2x2_ASAP7_75t_R _28082_ (.A(_05648_),
    .B(net5635),
    .Y(_05649_));
 AOI21x1_ASAP7_75t_R _28083_ (.A1(_05647_),
    .A2(_05649_),
    .B(net6070),
    .Y(_05650_));
 AOI21x1_ASAP7_75t_R _28084_ (.A1(_05333_),
    .A2(_05560_),
    .B(_05292_),
    .Y(_05651_));
 NAND2x1_ASAP7_75t_R _28085_ (.A(_05243_),
    .B(_05429_),
    .Y(_05652_));
 NAND3x1_ASAP7_75t_R _28086_ (.A(_05651_),
    .B(_05652_),
    .C(net5367),
    .Y(_05653_));
 AOI21x1_ASAP7_75t_R _28087_ (.A1(_05650_),
    .A2(_05653_),
    .B(net6060),
    .Y(_05654_));
 AND3x1_ASAP7_75t_R _28088_ (.A(net6072),
    .B(net5636),
    .C(_01323_),
    .Y(_05655_));
 OA21x2_ASAP7_75t_R _28089_ (.A1(_05655_),
    .A2(_05516_),
    .B(net5635),
    .Y(_05656_));
 OAI21x1_ASAP7_75t_R _28090_ (.A1(net4628),
    .A2(_05321_),
    .B(_05381_),
    .Y(_05657_));
 INVx1_ASAP7_75t_R _28091_ (.A(_05283_),
    .Y(_05658_));
 NOR2x1_ASAP7_75t_R _28092_ (.A(net5635),
    .B(net4843),
    .Y(_05659_));
 AND3x1_ASAP7_75t_R _28093_ (.A(_05140_),
    .B(net5639),
    .C(_05259_),
    .Y(_05660_));
 AOI21x1_ASAP7_75t_R _28094_ (.A1(_05658_),
    .A2(_05659_),
    .B(_05660_),
    .Y(_05661_));
 NAND2x1_ASAP7_75t_R _28095_ (.A(_05657_),
    .B(_05661_),
    .Y(_05662_));
 OAI21x1_ASAP7_75t_R _28096_ (.A1(_05656_),
    .A2(_05662_),
    .B(net6068),
    .Y(_05663_));
 NAND2x1_ASAP7_75t_R _28097_ (.A(_05654_),
    .B(_05663_),
    .Y(_05664_));
 NAND2x1_ASAP7_75t_R _28098_ (.A(net6071),
    .B(_05523_),
    .Y(_05665_));
 AOI21x1_ASAP7_75t_R _28099_ (.A1(_05459_),
    .A2(_05241_),
    .B(_05665_),
    .Y(_05666_));
 OAI21x1_ASAP7_75t_R _28100_ (.A1(_05414_),
    .A2(_05385_),
    .B(net6079),
    .Y(_05667_));
 AO21x1_ASAP7_75t_R _28101_ (.A1(_05359_),
    .A2(net6075),
    .B(net6070),
    .Y(_05668_));
 AOI21x1_ASAP7_75t_R _28102_ (.A1(net4438),
    .A2(_05667_),
    .B(_05668_),
    .Y(_05669_));
 OAI21x1_ASAP7_75t_R _28103_ (.A1(_05666_),
    .A2(_05669_),
    .B(net5634),
    .Y(_05670_));
 NAND2x1_ASAP7_75t_R _28104_ (.A(net4845),
    .B(_05345_),
    .Y(_05671_));
 OA21x2_ASAP7_75t_R _28105_ (.A1(_05501_),
    .A2(net6079),
    .B(net6071),
    .Y(_05672_));
 AOI21x1_ASAP7_75t_R _28106_ (.A1(_05671_),
    .A2(_05672_),
    .B(net5635),
    .Y(_05673_));
 INVx1_ASAP7_75t_R _28107_ (.A(_05451_),
    .Y(_05674_));
 OAI21x1_ASAP7_75t_R _28108_ (.A1(_05168_),
    .A2(_05674_),
    .B(net6073),
    .Y(_05675_));
 AOI21x1_ASAP7_75t_R _28109_ (.A1(net5095),
    .A2(_05333_),
    .B(net6068),
    .Y(_05676_));
 NAND3x1_ASAP7_75t_R _28110_ (.A(_05210_),
    .B(_05675_),
    .C(_05676_),
    .Y(_05677_));
 AOI21x1_ASAP7_75t_R _28111_ (.A1(_05673_),
    .A2(_05677_),
    .B(_05237_),
    .Y(_05678_));
 AOI21x1_ASAP7_75t_R _28112_ (.A1(_05670_),
    .A2(_05678_),
    .B(net6059),
    .Y(_05679_));
 NAND2x1_ASAP7_75t_R _28113_ (.A(_05664_),
    .B(_05679_),
    .Y(_05680_));
 AOI21x1_ASAP7_75t_R _28114_ (.A1(_01335_),
    .A2(net6080),
    .B(net6071),
    .Y(_05681_));
 NAND2x1_ASAP7_75t_R _28115_ (.A(net4620),
    .B(net5094),
    .Y(_05682_));
 AOI21x1_ASAP7_75t_R _28116_ (.A1(_05681_),
    .A2(_05682_),
    .B(net5367),
    .Y(_05683_));
 OAI21x1_ASAP7_75t_R _28117_ (.A1(net4457),
    .A2(_05224_),
    .B(_05404_),
    .Y(_05684_));
 NAND2x1_ASAP7_75t_R _28118_ (.A(_05683_),
    .B(_05684_),
    .Y(_05685_));
 AOI21x1_ASAP7_75t_R _28119_ (.A1(_05295_),
    .A2(_05554_),
    .B(net6062),
    .Y(_05686_));
 OAI21x1_ASAP7_75t_R _28120_ (.A1(_05438_),
    .A2(_05686_),
    .B(net5366),
    .Y(_05687_));
 AOI21x1_ASAP7_75t_R _28121_ (.A1(_05685_),
    .A2(_05687_),
    .B(_05237_),
    .Y(_05688_));
 INVx1_ASAP7_75t_R _28122_ (.A(_05668_),
    .Y(_05689_));
 NAND2x1_ASAP7_75t_R _28123_ (.A(_05622_),
    .B(_05689_),
    .Y(_05690_));
 AOI21x1_ASAP7_75t_R _28124_ (.A1(_05346_),
    .A2(_05228_),
    .B(net5634),
    .Y(_05691_));
 NAND2x1_ASAP7_75t_R _28125_ (.A(_05690_),
    .B(_05691_),
    .Y(_05692_));
 NAND2x1_ASAP7_75t_R _28126_ (.A(net6073),
    .B(_05434_),
    .Y(_05693_));
 NOR2x1_ASAP7_75t_R _28127_ (.A(net5641),
    .B(net5097),
    .Y(_05694_));
 OAI21x1_ASAP7_75t_R _28128_ (.A1(net4840),
    .A2(_05694_),
    .B(net6076),
    .Y(_05695_));
 AOI21x1_ASAP7_75t_R _28129_ (.A1(_05693_),
    .A2(_05695_),
    .B(net6071),
    .Y(_05696_));
 NAND2x1_ASAP7_75t_R _28130_ (.A(net4847),
    .B(_05398_),
    .Y(_05697_));
 OAI21x1_ASAP7_75t_R _28131_ (.A1(net4841),
    .A2(_05503_),
    .B(net6076),
    .Y(_05698_));
 AOI21x1_ASAP7_75t_R _28132_ (.A1(_05697_),
    .A2(_05698_),
    .B(net6066),
    .Y(_05699_));
 OAI21x1_ASAP7_75t_R _28133_ (.A1(_05696_),
    .A2(_05699_),
    .B(net5635),
    .Y(_05700_));
 AOI21x1_ASAP7_75t_R _28134_ (.A1(_05692_),
    .A2(_05700_),
    .B(net6060),
    .Y(_05701_));
 OAI21x1_ASAP7_75t_R _28135_ (.A1(_05688_),
    .A2(_05701_),
    .B(net6059),
    .Y(_05702_));
 NAND2x1_ASAP7_75t_R _28136_ (.A(_05680_),
    .B(_05702_),
    .Y(_00134_));
 AO21x1_ASAP7_75t_R _28137_ (.A1(net6078),
    .A2(_05364_),
    .B(_05621_),
    .Y(_05703_));
 NOR2x1_ASAP7_75t_R _28138_ (.A(net6075),
    .B(_05296_),
    .Y(_05704_));
 AOI21x1_ASAP7_75t_R _28139_ (.A1(net4429),
    .A2(_05190_),
    .B(net6078),
    .Y(_05705_));
 OAI21x1_ASAP7_75t_R _28140_ (.A1(_05704_),
    .A2(_05705_),
    .B(net6069),
    .Y(_05706_));
 AOI21x1_ASAP7_75t_R _28141_ (.A1(_05703_),
    .A2(_05706_),
    .B(net5632),
    .Y(_05707_));
 NAND2x1_ASAP7_75t_R _28142_ (.A(net6075),
    .B(net5095),
    .Y(_05708_));
 AOI21x1_ASAP7_75t_R _28143_ (.A1(_05708_),
    .A2(_05572_),
    .B(net6062),
    .Y(_05709_));
 AOI21x1_ASAP7_75t_R _28144_ (.A1(net5370),
    .A2(_05190_),
    .B(net6081),
    .Y(_05710_));
 OAI21x1_ASAP7_75t_R _28145_ (.A1(_05566_),
    .A2(_05710_),
    .B(net5632),
    .Y(_05711_));
 OAI21x1_ASAP7_75t_R _28146_ (.A1(_05709_),
    .A2(_05711_),
    .B(net6060),
    .Y(_05712_));
 NOR2x1_ASAP7_75t_R _28147_ (.A(_05712_),
    .B(_05707_),
    .Y(_05713_));
 NOR2x1_ASAP7_75t_R _28148_ (.A(net6071),
    .B(_05398_),
    .Y(_05714_));
 AO21x1_ASAP7_75t_R _28149_ (.A1(_05714_),
    .A2(_05554_),
    .B(net5366),
    .Y(_05715_));
 OAI21x1_ASAP7_75t_R _28150_ (.A1(net5095),
    .A2(net5375),
    .B(_05130_),
    .Y(_05716_));
 NOR2x1_ASAP7_75t_R _28151_ (.A(net6075),
    .B(_05716_),
    .Y(_05717_));
 NAND2x1_ASAP7_75t_R _28152_ (.A(_05553_),
    .B(_05404_),
    .Y(_05718_));
 NOR2x1_ASAP7_75t_R _28153_ (.A(_05717_),
    .B(_05718_),
    .Y(_05719_));
 OAI21x1_ASAP7_75t_R _28154_ (.A1(_05715_),
    .A2(_05719_),
    .B(_05237_),
    .Y(_05720_));
 NAND2x1_ASAP7_75t_R _28155_ (.A(net4430),
    .B(_05230_),
    .Y(_05721_));
 NAND2x1_ASAP7_75t_R _28156_ (.A(net4496),
    .B(_05349_),
    .Y(_05722_));
 AO21x1_ASAP7_75t_R _28157_ (.A1(_05721_),
    .A2(_05722_),
    .B(net6062),
    .Y(_05723_));
 AO21x1_ASAP7_75t_R _28158_ (.A1(_05470_),
    .A2(_05652_),
    .B(net6069),
    .Y(_05724_));
 AOI21x1_ASAP7_75t_R _28159_ (.A1(_05723_),
    .A2(_05724_),
    .B(net5632),
    .Y(_05725_));
 OAI21x1_ASAP7_75t_R _28160_ (.A1(_05720_),
    .A2(_05725_),
    .B(net6059),
    .Y(_05726_));
 AND3x1_ASAP7_75t_R _28161_ (.A(_05427_),
    .B(net4545),
    .C(net6079),
    .Y(_05727_));
 AO21x1_ASAP7_75t_R _28162_ (.A1(_05230_),
    .A2(net5094),
    .B(net6063),
    .Y(_05728_));
 OA21x2_ASAP7_75t_R _28163_ (.A1(_01338_),
    .A2(net6074),
    .B(_05170_),
    .Y(_05729_));
 AO21x1_ASAP7_75t_R _28164_ (.A1(_05427_),
    .A2(net4627),
    .B(net6079),
    .Y(_05730_));
 AOI21x1_ASAP7_75t_R _28165_ (.A1(_05729_),
    .A2(_05730_),
    .B(net5634),
    .Y(_05731_));
 OAI21x1_ASAP7_75t_R _28166_ (.A1(_05727_),
    .A2(_05728_),
    .B(_05731_),
    .Y(_05732_));
 NAND2x1_ASAP7_75t_R _28167_ (.A(net6073),
    .B(_05446_),
    .Y(_05733_));
 OA21x2_ASAP7_75t_R _28168_ (.A1(_05556_),
    .A2(net6073),
    .B(net6066),
    .Y(_05734_));
 AOI21x1_ASAP7_75t_R _28169_ (.A1(_05733_),
    .A2(_05734_),
    .B(net5367),
    .Y(_05735_));
 AO21x1_ASAP7_75t_R _28170_ (.A1(_05615_),
    .A2(net5641),
    .B(net6076),
    .Y(_05736_));
 NAND2x1_ASAP7_75t_R _28171_ (.A(_05581_),
    .B(_05736_),
    .Y(_05737_));
 AOI21x1_ASAP7_75t_R _28172_ (.A1(_05735_),
    .A2(_05737_),
    .B(_05237_),
    .Y(_05738_));
 AOI21x1_ASAP7_75t_R _28173_ (.A1(_05732_),
    .A2(_05738_),
    .B(net6059),
    .Y(_05739_));
 AO21x1_ASAP7_75t_R _28174_ (.A1(_05501_),
    .A2(_05339_),
    .B(net6075),
    .Y(_05740_));
 OAI21x1_ASAP7_75t_R _28175_ (.A1(net6078),
    .A2(_05716_),
    .B(_05740_),
    .Y(_05741_));
 NAND2x1_ASAP7_75t_R _28176_ (.A(_05130_),
    .B(net5367),
    .Y(_05742_));
 AOI21x1_ASAP7_75t_R _28177_ (.A1(_05346_),
    .A2(net4438),
    .B(_05742_),
    .Y(_05743_));
 AOI21x1_ASAP7_75t_R _28178_ (.A1(net5634),
    .A2(_05741_),
    .B(_05743_),
    .Y(_05744_));
 AOI21x1_ASAP7_75t_R _28179_ (.A1(_05560_),
    .A2(net5365),
    .B(net5367),
    .Y(_05745_));
 NAND2x1_ASAP7_75t_R _28180_ (.A(_05530_),
    .B(_05745_),
    .Y(_05746_));
 OA21x2_ASAP7_75t_R _28181_ (.A1(net4800),
    .A2(net6078),
    .B(net5367),
    .Y(_05747_));
 AOI21x1_ASAP7_75t_R _28182_ (.A1(_05747_),
    .A2(_05647_),
    .B(net6063),
    .Y(_05748_));
 AOI21x1_ASAP7_75t_R _28183_ (.A1(_05746_),
    .A2(_05748_),
    .B(net6060),
    .Y(_05749_));
 OAI21x1_ASAP7_75t_R _28184_ (.A1(net6069),
    .A2(_05744_),
    .B(_05749_),
    .Y(_05750_));
 NAND2x1_ASAP7_75t_R _28185_ (.A(_05739_),
    .B(_05750_),
    .Y(_05751_));
 OAI21x1_ASAP7_75t_R _28186_ (.A1(_05726_),
    .A2(_05713_),
    .B(_05751_),
    .Y(_00135_));
 NOR2x1_ASAP7_75t_R _28187_ (.A(net6668),
    .B(_00483_),
    .Y(_05752_));
 XOR2x2_ASAP7_75t_R _28188_ (.A(_11396_),
    .B(net6590),
    .Y(_05753_));
 XOR2x2_ASAP7_75t_R _28189_ (.A(_11428_),
    .B(_02981_),
    .Y(_05754_));
 NAND2x1_ASAP7_75t_R _28190_ (.A(_05753_),
    .B(_05754_),
    .Y(_05755_));
 OR2x2_ASAP7_75t_R _28191_ (.A(_05753_),
    .B(_05754_),
    .Y(_05756_));
 AOI21x1_ASAP7_75t_R _28192_ (.A1(_05755_),
    .A2(_05756_),
    .B(net6461),
    .Y(_05757_));
 OAI21x1_ASAP7_75t_R _28193_ (.A1(net6393),
    .A2(net6345),
    .B(net6505),
    .Y(_05758_));
 INVx1_ASAP7_75t_R _28194_ (.A(_00483_),
    .Y(_05759_));
 NOR2x1_ASAP7_75t_R _28195_ (.A(net6668),
    .B(_05759_),
    .Y(_05760_));
 XOR2x2_ASAP7_75t_R _28196_ (.A(_11430_),
    .B(_02981_),
    .Y(_05761_));
 XOR2x2_ASAP7_75t_R _28197_ (.A(_05761_),
    .B(_05753_),
    .Y(_05762_));
 NOR2x1_ASAP7_75t_R _28198_ (.A(net6461),
    .B(_05762_),
    .Y(_05763_));
 INVx1_ASAP7_75t_R _28199_ (.A(net6505),
    .Y(_05764_));
 OAI21x1_ASAP7_75t_R _28200_ (.A1(_05760_),
    .A2(net6344),
    .B(_05764_),
    .Y(_05765_));
 NAND2x1_ASAP7_75t_R _28201_ (.A(_05758_),
    .B(_05765_),
    .Y(_05766_));
 NOR2x1_ASAP7_75t_R _28203_ (.A(net6668),
    .B(_00484_),
    .Y(_05767_));
 INVx1_ASAP7_75t_R _28204_ (.A(_05767_),
    .Y(_05768_));
 XOR2x2_ASAP7_75t_R _28205_ (.A(net6442),
    .B(net6554),
    .Y(_05769_));
 NOR2x1_ASAP7_75t_R _28206_ (.A(net6444),
    .B(_05769_),
    .Y(_05770_));
 INVx1_ASAP7_75t_R _28207_ (.A(net6444),
    .Y(_05771_));
 XOR2x2_ASAP7_75t_R _28208_ (.A(_11565_),
    .B(_11415_),
    .Y(_05772_));
 NOR2x1_ASAP7_75t_R _28209_ (.A(net6385),
    .B(net6384),
    .Y(_05773_));
 OAI21x1_ASAP7_75t_R _28210_ (.A1(_05770_),
    .A2(_05773_),
    .B(net6668),
    .Y(_05774_));
 NAND2x1_ASAP7_75t_R _28211_ (.A(_05768_),
    .B(_05774_),
    .Y(_05775_));
 INVx1_ASAP7_75t_R _28212_ (.A(net6512),
    .Y(_05776_));
 XOR2x2_ASAP7_75t_R _28213_ (.A(_05775_),
    .B(_05776_),
    .Y(_05777_));
 XOR2x2_ASAP7_75t_R _28215_ (.A(net6641),
    .B(net6589),
    .Y(_05778_));
 NAND2x1_ASAP7_75t_R _28216_ (.A(net6400),
    .B(_05778_),
    .Y(_05779_));
 XNOR2x2_ASAP7_75t_R _28217_ (.A(net6641),
    .B(net6589),
    .Y(_05780_));
 NAND2x1_ASAP7_75t_R _28218_ (.A(net6558),
    .B(_05780_),
    .Y(_05781_));
 AOI21x1_ASAP7_75t_R _28219_ (.A1(_05779_),
    .A2(_05781_),
    .B(_03026_),
    .Y(_05782_));
 XOR2x2_ASAP7_75t_R _28220_ (.A(net6589),
    .B(net6558),
    .Y(_05783_));
 NAND2x1_ASAP7_75t_R _28221_ (.A(net6641),
    .B(_05783_),
    .Y(_05784_));
 INVx1_ASAP7_75t_R _28222_ (.A(net6641),
    .Y(_05785_));
 XNOR2x2_ASAP7_75t_R _28223_ (.A(net6589),
    .B(net6558),
    .Y(_05786_));
 NAND2x1_ASAP7_75t_R _28224_ (.A(_05785_),
    .B(_05786_),
    .Y(_05787_));
 AOI21x1_ASAP7_75t_R _28225_ (.A1(_05784_),
    .A2(_05787_),
    .B(_03014_),
    .Y(_05788_));
 OAI21x1_ASAP7_75t_R _28226_ (.A1(_05782_),
    .A2(_05788_),
    .B(net6668),
    .Y(_05789_));
 OR2x2_ASAP7_75t_R _28227_ (.A(net6668),
    .B(_00485_),
    .Y(_05790_));
 NAND3x1_ASAP7_75t_R _28228_ (.A(_05789_),
    .B(net6499),
    .C(_05790_),
    .Y(_05791_));
 AO21x1_ASAP7_75t_R _28229_ (.A1(_05789_),
    .A2(_05790_),
    .B(net6499),
    .Y(_05792_));
 NAND2x1_ASAP7_75t_R _28230_ (.A(_05791_),
    .B(_05792_),
    .Y(_05793_));
 AOI21x1_ASAP7_75t_R _28232_ (.A1(_05768_),
    .A2(_05774_),
    .B(_05776_),
    .Y(_05794_));
 AND2x2_ASAP7_75t_R _28233_ (.A(net6464),
    .B(_00484_),
    .Y(_05795_));
 INVx1_ASAP7_75t_R _28234_ (.A(_05795_),
    .Y(_05796_));
 XOR2x2_ASAP7_75t_R _28235_ (.A(_05771_),
    .B(_05772_),
    .Y(_05797_));
 NAND2x1p5_ASAP7_75t_R _28236_ (.A(net6668),
    .B(_05797_),
    .Y(_05798_));
 AOI21x1_ASAP7_75t_R _28237_ (.A1(_05798_),
    .A2(_05796_),
    .B(net6512),
    .Y(_05799_));
 NOR2x2_ASAP7_75t_R _28238_ (.A(_05799_),
    .B(_05794_),
    .Y(_05800_));
 INVx1_ASAP7_75t_R _28241_ (.A(net6499),
    .Y(_05802_));
 NAND3x1_ASAP7_75t_R _28242_ (.A(_05789_),
    .B(_05802_),
    .C(_05790_),
    .Y(_05803_));
 AO21x1_ASAP7_75t_R _28243_ (.A1(_05789_),
    .A2(_05790_),
    .B(_05802_),
    .Y(_05804_));
 NAND2x1_ASAP7_75t_R _28244_ (.A(_05803_),
    .B(_05804_),
    .Y(_05805_));
 NAND2x1_ASAP7_75t_R _28246_ (.A(net5623),
    .B(net5628),
    .Y(_05806_));
 INVx1_ASAP7_75t_R _28249_ (.A(_01345_),
    .Y(_05809_));
 AOI21x1_ASAP7_75t_R _28250_ (.A1(net6054),
    .A2(net6053),
    .B(_05809_),
    .Y(_05810_));
 INVx1_ASAP7_75t_R _28251_ (.A(_00650_),
    .Y(_05811_));
 XOR2x2_ASAP7_75t_R _28252_ (.A(_11468_),
    .B(_05811_),
    .Y(_05812_));
 NOR2x1_ASAP7_75t_R _28253_ (.A(_05812_),
    .B(_03043_),
    .Y(_05813_));
 AO21x1_ASAP7_75t_R _28254_ (.A1(_03043_),
    .A2(_05812_),
    .B(net6461),
    .Y(_05814_));
 NAND2x1_ASAP7_75t_R _28255_ (.A(_00511_),
    .B(net6461),
    .Y(_05815_));
 OAI21x1_ASAP7_75t_R _28256_ (.A1(_05813_),
    .A2(_05814_),
    .B(_05815_),
    .Y(_05816_));
 XOR2x2_ASAP7_75t_R _28257_ (.A(_05816_),
    .B(net6498),
    .Y(_05817_));
 NOR2x1_ASAP7_75t_R _28259_ (.A(net4729),
    .B(net6046),
    .Y(_05819_));
 OA21x2_ASAP7_75t_R _28260_ (.A1(net5364),
    .A2(net5617),
    .B(_05819_),
    .Y(_05820_));
 INVx1_ASAP7_75t_R _28263_ (.A(_01344_),
    .Y(_05823_));
 AO21x1_ASAP7_75t_R _28264_ (.A1(net6057),
    .A2(net6058),
    .B(_05823_),
    .Y(_05824_));
 INVx1_ASAP7_75t_R _28265_ (.A(_05824_),
    .Y(_05825_));
 INVx1_ASAP7_75t_R _28266_ (.A(_01348_),
    .Y(_05826_));
 NOR2x1_ASAP7_75t_R _28268_ (.A(_05826_),
    .B(net5620),
    .Y(_05828_));
 OA21x2_ASAP7_75t_R _28271_ (.A1(_05825_),
    .A2(_05828_),
    .B(net6049),
    .Y(_05831_));
 XNOR2x2_ASAP7_75t_R _28272_ (.A(_00651_),
    .B(_11480_),
    .Y(_05832_));
 XOR2x2_ASAP7_75t_R _28273_ (.A(_11507_),
    .B(_03059_),
    .Y(_05833_));
 NOR2x1_ASAP7_75t_R _28274_ (.A(_05832_),
    .B(_05833_),
    .Y(_05834_));
 AO21x1_ASAP7_75t_R _28275_ (.A1(_05833_),
    .A2(_05832_),
    .B(net6461),
    .Y(_05835_));
 NAND2x1_ASAP7_75t_R _28276_ (.A(_00510_),
    .B(net6461),
    .Y(_05836_));
 OAI21x1_ASAP7_75t_R _28277_ (.A1(_05834_),
    .A2(_05835_),
    .B(_05836_),
    .Y(_05837_));
 XNOR2x2_ASAP7_75t_R _28278_ (.A(net6497),
    .B(_05837_),
    .Y(_05838_));
 INVx2_ASAP7_75t_R _28279_ (.A(_05838_),
    .Y(_05839_));
 OR3x1_ASAP7_75t_R _28282_ (.A(_05820_),
    .B(_05831_),
    .C(net5612),
    .Y(_05842_));
 OAI21x1_ASAP7_75t_R _28283_ (.A1(_05752_),
    .A2(_05757_),
    .B(_05764_),
    .Y(_05843_));
 OAI21x1_ASAP7_75t_R _28284_ (.A1(_05760_),
    .A2(_05763_),
    .B(net6505),
    .Y(_05844_));
 NAND2x1_ASAP7_75t_R _28285_ (.A(_05843_),
    .B(_05844_),
    .Y(_05845_));
 NAND2x1_ASAP7_75t_R _28286_ (.A(net5617),
    .B(net5607),
    .Y(_05846_));
 AOI21x1_ASAP7_75t_R _28289_ (.A1(net5616),
    .A2(net5626),
    .B(net6052),
    .Y(_05849_));
 NAND2x1_ASAP7_75t_R _28290_ (.A(net5363),
    .B(_05849_),
    .Y(_05850_));
 OAI21x1_ASAP7_75t_R _28291_ (.A1(net6056),
    .A2(net6055),
    .B(_05793_),
    .Y(_05851_));
 INVx1_ASAP7_75t_R _28292_ (.A(net6498),
    .Y(_05852_));
 XOR2x2_ASAP7_75t_R _28293_ (.A(_05816_),
    .B(_05852_),
    .Y(_05853_));
 AOI21x1_ASAP7_75t_R _28295_ (.A1(net5617),
    .A2(net5630),
    .B(net6041),
    .Y(_05855_));
 AOI21x1_ASAP7_75t_R _28298_ (.A1(net5362),
    .A2(_05855_),
    .B(net6045),
    .Y(_05858_));
 XOR2x2_ASAP7_75t_R _28299_ (.A(_00587_),
    .B(_00588_),
    .Y(_05859_));
 XOR2x2_ASAP7_75t_R _28300_ (.A(_11504_),
    .B(net6556),
    .Y(_05860_));
 NAND2x1_ASAP7_75t_R _28301_ (.A(_05859_),
    .B(_05860_),
    .Y(_05861_));
 INVx1_ASAP7_75t_R _28302_ (.A(_05859_),
    .Y(_05862_));
 XNOR2x2_ASAP7_75t_R _28303_ (.A(net6556),
    .B(_11504_),
    .Y(_05863_));
 NAND2x1_ASAP7_75t_R _28304_ (.A(_05862_),
    .B(_05863_),
    .Y(_05864_));
 AOI21x1_ASAP7_75t_R _28305_ (.A1(_05861_),
    .A2(_05864_),
    .B(net6463),
    .Y(_05865_));
 NOR2x1_ASAP7_75t_R _28306_ (.A(net6665),
    .B(_00509_),
    .Y(_05866_));
 OA21x2_ASAP7_75t_R _28307_ (.A1(_05865_),
    .A2(_05866_),
    .B(net6496),
    .Y(_05867_));
 INVx1_ASAP7_75t_R _28308_ (.A(_00509_),
    .Y(_05868_));
 AOI211x1_ASAP7_75t_R _28309_ (.A1(net6461),
    .A2(_05868_),
    .B(_05865_),
    .C(net6496),
    .Y(_05869_));
 NOR2x1_ASAP7_75t_R _28310_ (.A(_05867_),
    .B(_05869_),
    .Y(_05870_));
 AOI21x1_ASAP7_75t_R _28313_ (.A1(_05850_),
    .A2(_05858_),
    .B(net5605),
    .Y(_05873_));
 XOR2x2_ASAP7_75t_R _28314_ (.A(_00588_),
    .B(_00589_),
    .Y(_05874_));
 XOR2x2_ASAP7_75t_R _28315_ (.A(_05874_),
    .B(_11508_),
    .Y(_05875_));
 XOR2x2_ASAP7_75t_R _28316_ (.A(_05875_),
    .B(_11455_),
    .Y(_05876_));
 NOR2x1_ASAP7_75t_R _28317_ (.A(net6665),
    .B(_00507_),
    .Y(_05877_));
 AO21x1_ASAP7_75t_R _28318_ (.A1(_05876_),
    .A2(net6665),
    .B(_05877_),
    .Y(_05878_));
 XNOR2x2_ASAP7_75t_R _28319_ (.A(net6495),
    .B(_05878_),
    .Y(_05879_));
 INVx1_ASAP7_75t_R _28320_ (.A(_05879_),
    .Y(_05880_));
 AOI21x1_ASAP7_75t_R _28322_ (.A1(net6058),
    .A2(net6057),
    .B(net4995),
    .Y(_05882_));
 NAND2x1_ASAP7_75t_R _28324_ (.A(net4728),
    .B(net6046),
    .Y(_05884_));
 AOI21x1_ASAP7_75t_R _28326_ (.A1(net5620),
    .A2(net5607),
    .B(net6052),
    .Y(_05885_));
 INVx1_ASAP7_75t_R _28327_ (.A(net5361),
    .Y(_05886_));
 AO21x1_ASAP7_75t_R _28329_ (.A1(net4729),
    .A2(net6041),
    .B(net6045),
    .Y(_05888_));
 AOI21x1_ASAP7_75t_R _28330_ (.A1(_05884_),
    .A2(_05886_),
    .B(_05888_),
    .Y(_05889_));
 AO21x1_ASAP7_75t_R _28331_ (.A1(net6053),
    .A2(net6054),
    .B(_01344_),
    .Y(_05890_));
 AOI21x1_ASAP7_75t_R _28333_ (.A1(net6058),
    .A2(net6057),
    .B(_01348_),
    .Y(_05892_));
 NOR2x1_ASAP7_75t_R _28334_ (.A(_05892_),
    .B(_05817_),
    .Y(_05893_));
 NAND2x1_ASAP7_75t_R _28335_ (.A(_05890_),
    .B(_05893_),
    .Y(_05894_));
 AOI21x1_ASAP7_75t_R _28336_ (.A1(net6054),
    .A2(net6053),
    .B(net5253),
    .Y(_05895_));
 INVx1_ASAP7_75t_R _28337_ (.A(_05895_),
    .Y(_05896_));
 AO21x1_ASAP7_75t_R _28340_ (.A1(_05824_),
    .A2(_05896_),
    .B(net6040),
    .Y(_05899_));
 AOI21x1_ASAP7_75t_R _28343_ (.A1(_05894_),
    .A2(_05899_),
    .B(net5612),
    .Y(_05902_));
 OAI21x1_ASAP7_75t_R _28345_ (.A1(_05889_),
    .A2(_05902_),
    .B(net5605),
    .Y(_05904_));
 NAND2x1_ASAP7_75t_R _28346_ (.A(net5604),
    .B(_05904_),
    .Y(_05905_));
 AOI21x1_ASAP7_75t_R _28347_ (.A1(_05842_),
    .A2(_05873_),
    .B(_05905_),
    .Y(_05906_));
 AOI21x1_ASAP7_75t_R _28349_ (.A1(net5622),
    .A2(net5618),
    .B(net6049),
    .Y(_05908_));
 NOR2x1_ASAP7_75t_R _28350_ (.A(net5609),
    .B(_05908_),
    .Y(_05909_));
 INVx1_ASAP7_75t_R _28351_ (.A(_01351_),
    .Y(_05910_));
 AOI21x1_ASAP7_75t_R _28352_ (.A1(net6054),
    .A2(net6053),
    .B(_05910_),
    .Y(_05911_));
 NOR2x1p5_ASAP7_75t_R _28353_ (.A(_05911_),
    .B(net6042),
    .Y(_05912_));
 OAI21x1_ASAP7_75t_R _28354_ (.A1(net5625),
    .A2(net5364),
    .B(_05912_),
    .Y(_05913_));
 AO21x1_ASAP7_75t_R _28355_ (.A1(_05909_),
    .A2(_05913_),
    .B(net5606),
    .Y(_05914_));
 INVx3_ASAP7_75t_R _28356_ (.A(_05810_),
    .Y(_05915_));
 AOI21x1_ASAP7_75t_R _28357_ (.A1(net5272),
    .A2(net5623),
    .B(net6042),
    .Y(_05916_));
 OAI21x1_ASAP7_75t_R _28358_ (.A1(net5623),
    .A2(net5625),
    .B(net6042),
    .Y(_05917_));
 NAND2x1_ASAP7_75t_R _28359_ (.A(net5618),
    .B(net5628),
    .Y(_05918_));
 INVx1_ASAP7_75t_R _28360_ (.A(_05918_),
    .Y(_05919_));
 OAI21x1_ASAP7_75t_R _28361_ (.A1(_05917_),
    .A2(_05919_),
    .B(net5609),
    .Y(_05920_));
 AOI21x1_ASAP7_75t_R _28362_ (.A1(net4542),
    .A2(_05916_),
    .B(_05920_),
    .Y(_05921_));
 OAI21x1_ASAP7_75t_R _28365_ (.A1(_05914_),
    .A2(_05921_),
    .B(net6039),
    .Y(_05924_));
 INVx1_ASAP7_75t_R _28366_ (.A(net6054),
    .Y(_05925_));
 INVx1_ASAP7_75t_R _28367_ (.A(net6053),
    .Y(_05926_));
 INVx1_ASAP7_75t_R _28368_ (.A(_01346_),
    .Y(_05927_));
 OAI21x1_ASAP7_75t_R _28369_ (.A1(_05925_),
    .A2(_05926_),
    .B(_05927_),
    .Y(_05928_));
 OAI21x1_ASAP7_75t_R _28370_ (.A1(net5615),
    .A2(net5628),
    .B(net4837),
    .Y(_05929_));
 AND2x2_ASAP7_75t_R _28372_ (.A(_05929_),
    .B(net6043),
    .Y(_05931_));
 NAND2x1_ASAP7_75t_R _28373_ (.A(net5627),
    .B(net5624),
    .Y(_05932_));
 AOI21x1_ASAP7_75t_R _28374_ (.A1(net5623),
    .A2(net5618),
    .B(net6044),
    .Y(_05933_));
 OAI21x1_ASAP7_75t_R _28375_ (.A1(net5622),
    .A2(_05932_),
    .B(_05933_),
    .Y(_05934_));
 NAND2x1_ASAP7_75t_R _28376_ (.A(net6045),
    .B(_05934_),
    .Y(_05935_));
 NOR2x1_ASAP7_75t_R _28377_ (.A(_05931_),
    .B(_05935_),
    .Y(_05936_));
 INVx1_ASAP7_75t_R _28378_ (.A(_01353_),
    .Y(_05937_));
 AO21x1_ASAP7_75t_R _28379_ (.A1(net6053),
    .A2(net6054),
    .B(_05937_),
    .Y(_05938_));
 AO21x1_ASAP7_75t_R _28380_ (.A1(net5357),
    .A2(net4834),
    .B(net6045),
    .Y(_05939_));
 INVx1_ASAP7_75t_R _28381_ (.A(net6393),
    .Y(_05940_));
 NAND2x1_ASAP7_75t_R _28382_ (.A(net6673),
    .B(net6381),
    .Y(_05941_));
 AOI21x1_ASAP7_75t_R _28383_ (.A1(_05940_),
    .A2(_05941_),
    .B(net6505),
    .Y(_05942_));
 AOI211x1_ASAP7_75t_R _28384_ (.A1(net6381),
    .A2(net6673),
    .B(net6393),
    .C(_05764_),
    .Y(_05943_));
 OAI21x1_ASAP7_75t_R _28385_ (.A1(_05942_),
    .A2(_05943_),
    .B(_05805_),
    .Y(_05944_));
 INVx1_ASAP7_75t_R _28386_ (.A(_05944_),
    .Y(_05945_));
 OAI21x1_ASAP7_75t_R _28387_ (.A1(net5624),
    .A2(net5364),
    .B(net6041),
    .Y(_05946_));
 NOR2x1_ASAP7_75t_R _28388_ (.A(_05945_),
    .B(_05946_),
    .Y(_05947_));
 OAI21x1_ASAP7_75t_R _28389_ (.A1(_05939_),
    .A2(_05947_),
    .B(net5606),
    .Y(_05948_));
 NOR2x1_ASAP7_75t_R _28390_ (.A(_05936_),
    .B(_05948_),
    .Y(_05949_));
 XOR2x2_ASAP7_75t_R _28391_ (.A(_00589_),
    .B(net6640),
    .Y(_05950_));
 XOR2x2_ASAP7_75t_R _28392_ (.A(_05950_),
    .B(_00685_),
    .Y(_05951_));
 XOR2x2_ASAP7_75t_R _28393_ (.A(_05951_),
    .B(_11567_),
    .Y(_05952_));
 NOR2x1_ASAP7_75t_R _28394_ (.A(net6665),
    .B(_00506_),
    .Y(_05953_));
 AO21x1_ASAP7_75t_R _28395_ (.A1(_05952_),
    .A2(net6665),
    .B(_05953_),
    .Y(_05954_));
 XOR2x2_ASAP7_75t_R _28396_ (.A(_05954_),
    .B(_00899_),
    .Y(_05955_));
 OAI21x1_ASAP7_75t_R _28397_ (.A1(_05924_),
    .A2(_05949_),
    .B(net6038),
    .Y(_05956_));
 AO21x1_ASAP7_75t_R _28398_ (.A1(net6057),
    .A2(net6058),
    .B(_05910_),
    .Y(_05957_));
 OAI21x1_ASAP7_75t_R _28399_ (.A1(net5623),
    .A2(net5624),
    .B(_05957_),
    .Y(_05958_));
 AOI21x1_ASAP7_75t_R _28400_ (.A1(_05944_),
    .A2(_05958_),
    .B(net6047),
    .Y(_05959_));
 AO21x1_ASAP7_75t_R _28401_ (.A1(net6057),
    .A2(net6058),
    .B(_01346_),
    .Y(_05960_));
 INVx1_ASAP7_75t_R _28402_ (.A(_05960_),
    .Y(_05961_));
 NAND2x1_ASAP7_75t_R _28403_ (.A(net6043),
    .B(_05961_),
    .Y(_05962_));
 AOI21x1_ASAP7_75t_R _28404_ (.A1(_05890_),
    .A2(net5357),
    .B(net5611),
    .Y(_05963_));
 NAND2x1_ASAP7_75t_R _28405_ (.A(_05962_),
    .B(_05963_),
    .Y(_05964_));
 AOI21x1_ASAP7_75t_R _28407_ (.A1(net6058),
    .A2(net6057),
    .B(net5253),
    .Y(_05966_));
 NOR2x1_ASAP7_75t_R _28408_ (.A(_05966_),
    .B(net6052),
    .Y(_05967_));
 AO21x1_ASAP7_75t_R _28409_ (.A1(_01361_),
    .A2(net6048),
    .B(_05967_),
    .Y(_05968_));
 INVx1_ASAP7_75t_R _28410_ (.A(_05870_),
    .Y(_05969_));
 AOI21x1_ASAP7_75t_R _28412_ (.A1(net5611),
    .A2(_05968_),
    .B(net5355),
    .Y(_05971_));
 OA21x2_ASAP7_75t_R _28413_ (.A1(_05959_),
    .A2(_05964_),
    .B(_05971_),
    .Y(_05972_));
 OA21x2_ASAP7_75t_R _28414_ (.A1(net4835),
    .A2(_05853_),
    .B(_05839_),
    .Y(_05973_));
 INVx1_ASAP7_75t_R _28415_ (.A(_05973_),
    .Y(_05974_));
 INVx1_ASAP7_75t_R _28416_ (.A(_05758_),
    .Y(_05975_));
 INVx1_ASAP7_75t_R _28417_ (.A(_05765_),
    .Y(_05976_));
 OAI21x1_ASAP7_75t_R _28418_ (.A1(_05975_),
    .A2(_05976_),
    .B(_05805_),
    .Y(_05977_));
 OA21x2_ASAP7_75t_R _28419_ (.A1(_05977_),
    .A2(net5626),
    .B(net4839),
    .Y(_05978_));
 OAI21x1_ASAP7_75t_R _28421_ (.A1(_05974_),
    .A2(_05978_),
    .B(net5355),
    .Y(_05980_));
 INVx1_ASAP7_75t_R _28422_ (.A(_05977_),
    .Y(_05981_));
 NAND2x1_ASAP7_75t_R _28423_ (.A(net5618),
    .B(_05981_),
    .Y(_05982_));
 INVx1_ASAP7_75t_R _28424_ (.A(net5275),
    .Y(_05983_));
 OA21x2_ASAP7_75t_R _28425_ (.A1(_05983_),
    .A2(net5616),
    .B(net6052),
    .Y(_05984_));
 NOR2x1_ASAP7_75t_R _28427_ (.A(net6052),
    .B(net4836),
    .Y(_05986_));
 AOI211x1_ASAP7_75t_R _28428_ (.A1(_05982_),
    .A2(net4833),
    .B(_05986_),
    .C(net5610),
    .Y(_05987_));
 OAI21x1_ASAP7_75t_R _28429_ (.A1(_05980_),
    .A2(_05987_),
    .B(net5604),
    .Y(_05988_));
 OAI21x1_ASAP7_75t_R _28430_ (.A1(net6056),
    .A2(net6055),
    .B(_05805_),
    .Y(_05989_));
 INVx1_ASAP7_75t_R _28431_ (.A(_05989_),
    .Y(_05990_));
 NOR2x1_ASAP7_75t_R _28432_ (.A(_05826_),
    .B(net5616),
    .Y(_05991_));
 OA21x2_ASAP7_75t_R _28434_ (.A1(_05990_),
    .A2(net4832),
    .B(net6049),
    .Y(_05993_));
 AOI21x1_ASAP7_75t_R _28435_ (.A1(net5616),
    .A2(net5627),
    .B(net6049),
    .Y(_05994_));
 INVx2_ASAP7_75t_R _28436_ (.A(_05966_),
    .Y(_05995_));
 AO21x1_ASAP7_75t_R _28437_ (.A1(_05994_),
    .A2(_05995_),
    .B(net5611),
    .Y(_05996_));
 NOR2x1_ASAP7_75t_R _28439_ (.A(net6045),
    .B(_05912_),
    .Y(_05998_));
 AO21x1_ASAP7_75t_R _28440_ (.A1(_05824_),
    .A2(_05928_),
    .B(net6052),
    .Y(_05999_));
 AOI21x1_ASAP7_75t_R _28441_ (.A1(_05998_),
    .A2(_05999_),
    .B(net5606),
    .Y(_06000_));
 OAI21x1_ASAP7_75t_R _28442_ (.A1(_05993_),
    .A2(_05996_),
    .B(_06000_),
    .Y(_06001_));
 AOI21x1_ASAP7_75t_R _28443_ (.A1(net6054),
    .A2(net6053),
    .B(_01349_),
    .Y(_06002_));
 NOR2x1_ASAP7_75t_R _28444_ (.A(net5273),
    .B(net5616),
    .Y(_06003_));
 OAI21x1_ASAP7_75t_R _28446_ (.A1(net5090),
    .A2(_06003_),
    .B(net6043),
    .Y(_06005_));
 NOR2x1p5_ASAP7_75t_R _28447_ (.A(net6041),
    .B(_05810_),
    .Y(_06006_));
 NOR2x1_ASAP7_75t_R _28448_ (.A(net6045),
    .B(_06006_),
    .Y(_06007_));
 AOI21x1_ASAP7_75t_R _28449_ (.A1(_06007_),
    .A2(_06005_),
    .B(net5355),
    .Y(_06008_));
 AO21x1_ASAP7_75t_R _28450_ (.A1(net6057),
    .A2(net6058),
    .B(net5274),
    .Y(_06009_));
 OA21x2_ASAP7_75t_R _28452_ (.A1(net5089),
    .A2(net6048),
    .B(net6045),
    .Y(_06011_));
 NAND2x1_ASAP7_75t_R _28453_ (.A(_06011_),
    .B(_05934_),
    .Y(_06012_));
 AOI21x1_ASAP7_75t_R _28454_ (.A1(_06012_),
    .A2(_06008_),
    .B(net5604),
    .Y(_06013_));
 AOI21x1_ASAP7_75t_R _28455_ (.A1(_06013_),
    .A2(_06001_),
    .B(net6038),
    .Y(_06014_));
 OAI21x1_ASAP7_75t_R _28456_ (.A1(_05972_),
    .A2(_05988_),
    .B(_06014_),
    .Y(_06015_));
 OAI21x1_ASAP7_75t_R _28457_ (.A1(_05906_),
    .A2(_05956_),
    .B(_06015_),
    .Y(_00136_));
 OAI21x1_ASAP7_75t_R _28458_ (.A1(net5616),
    .A2(net5608),
    .B(net6052),
    .Y(_06016_));
 NAND2x1_ASAP7_75t_R _28459_ (.A(_05944_),
    .B(_06016_),
    .Y(_06017_));
 OA21x2_ASAP7_75t_R _28460_ (.A1(net5087),
    .A2(net6050),
    .B(net5611),
    .Y(_06018_));
 INVx1_ASAP7_75t_R _28461_ (.A(_06018_),
    .Y(_06019_));
 OAI21x1_ASAP7_75t_R _28462_ (.A1(_06017_),
    .A2(_06019_),
    .B(net5606),
    .Y(_06020_));
 NOR2x1_ASAP7_75t_R _28463_ (.A(_05882_),
    .B(_05853_),
    .Y(_06021_));
 AO21x1_ASAP7_75t_R _28464_ (.A1(_06021_),
    .A2(net4834),
    .B(net5611),
    .Y(_06022_));
 NOR2x1_ASAP7_75t_R _28465_ (.A(_06022_),
    .B(_05959_),
    .Y(_06023_));
 OAI21x1_ASAP7_75t_R _28466_ (.A1(_06020_),
    .A2(_06023_),
    .B(net5604),
    .Y(_06024_));
 OAI21x1_ASAP7_75t_R _28467_ (.A1(net5615),
    .A2(net5625),
    .B(net6052),
    .Y(_06025_));
 OAI21x1_ASAP7_75t_R _28468_ (.A1(net4729),
    .A2(_06025_),
    .B(net5610),
    .Y(_06026_));
 INVx1_ASAP7_75t_R _28469_ (.A(_05911_),
    .Y(_06027_));
 AND3x1_ASAP7_75t_R _28470_ (.A(_05851_),
    .B(net6042),
    .C(_06027_),
    .Y(_06028_));
 OAI21x1_ASAP7_75t_R _28471_ (.A1(_06026_),
    .A2(_06028_),
    .B(net5355),
    .Y(_06029_));
 NOR2x1_ASAP7_75t_R _28472_ (.A(net5616),
    .B(net6042),
    .Y(_06030_));
 NAND2x1_ASAP7_75t_R _28473_ (.A(_06030_),
    .B(_05918_),
    .Y(_06031_));
 NAND2x1_ASAP7_75t_R _28474_ (.A(net5363),
    .B(_05994_),
    .Y(_06032_));
 NAND2x1_ASAP7_75t_R _28475_ (.A(_06031_),
    .B(_06032_),
    .Y(_06033_));
 NOR2x1_ASAP7_75t_R _28476_ (.A(net5611),
    .B(_06033_),
    .Y(_06034_));
 NOR2x1_ASAP7_75t_R _28477_ (.A(_06029_),
    .B(_06034_),
    .Y(_06035_));
 INVx1_ASAP7_75t_R _28478_ (.A(_05955_),
    .Y(_06036_));
 OAI21x1_ASAP7_75t_R _28479_ (.A1(_06024_),
    .A2(_06035_),
    .B(_06036_),
    .Y(_06037_));
 INVx2_ASAP7_75t_R _28480_ (.A(_06006_),
    .Y(_06038_));
 NOR2x1_ASAP7_75t_R _28481_ (.A(_06003_),
    .B(net4455),
    .Y(_06039_));
 AO21x1_ASAP7_75t_R _28483_ (.A1(net6053),
    .A2(net6054),
    .B(_05823_),
    .Y(_06041_));
 AND3x1_ASAP7_75t_R _28484_ (.A(net5362),
    .B(net6041),
    .C(_06041_),
    .Y(_06042_));
 OAI21x1_ASAP7_75t_R _28485_ (.A1(_06039_),
    .A2(_06042_),
    .B(net5611),
    .Y(_06043_));
 NOR2x1_ASAP7_75t_R _28486_ (.A(net5623),
    .B(net5625),
    .Y(_06044_));
 INVx1_ASAP7_75t_R _28487_ (.A(_06044_),
    .Y(_06045_));
 AO21x1_ASAP7_75t_R _28488_ (.A1(_06045_),
    .A2(_05967_),
    .B(net5611),
    .Y(_06046_));
 OA21x2_ASAP7_75t_R _28489_ (.A1(net5627),
    .A2(net5618),
    .B(net5357),
    .Y(_06047_));
 OA21x2_ASAP7_75t_R _28490_ (.A1(_06046_),
    .A2(_06047_),
    .B(net5606),
    .Y(_06048_));
 NOR2x1_ASAP7_75t_R _28491_ (.A(net5273),
    .B(net6052),
    .Y(_06049_));
 AO21x1_ASAP7_75t_R _28492_ (.A1(_06049_),
    .A2(net5616),
    .B(net5610),
    .Y(_06050_));
 OAI21x1_ASAP7_75t_R _28493_ (.A1(net5618),
    .A2(net5607),
    .B(net5623),
    .Y(_06051_));
 AOI21x1_ASAP7_75t_R _28494_ (.A1(_06051_),
    .A2(net4541),
    .B(net6041),
    .Y(_06052_));
 NOR2x1_ASAP7_75t_R _28495_ (.A(_06050_),
    .B(_06052_),
    .Y(_06053_));
 OAI21x1_ASAP7_75t_R _28496_ (.A1(net5618),
    .A2(net5607),
    .B(net5616),
    .Y(_06054_));
 NOR2x1_ASAP7_75t_R _28497_ (.A(net6048),
    .B(net5353),
    .Y(_06055_));
 AO21x1_ASAP7_75t_R _28498_ (.A1(net6057),
    .A2(net6058),
    .B(_05937_),
    .Y(_06056_));
 NAND2x1_ASAP7_75t_R _28499_ (.A(net6052),
    .B(_06056_),
    .Y(_06057_));
 OAI21x1_ASAP7_75t_R _28500_ (.A1(_05945_),
    .A2(_06057_),
    .B(net5611),
    .Y(_06058_));
 OAI21x1_ASAP7_75t_R _28501_ (.A1(_06055_),
    .A2(_06058_),
    .B(net5355),
    .Y(_06059_));
 OAI21x1_ASAP7_75t_R _28502_ (.A1(_06053_),
    .A2(_06059_),
    .B(net6039),
    .Y(_06060_));
 AOI21x1_ASAP7_75t_R _28503_ (.A1(_06043_),
    .A2(_06048_),
    .B(_06060_),
    .Y(_06061_));
 OAI21x1_ASAP7_75t_R _28504_ (.A1(net6052),
    .A2(_05851_),
    .B(net5610),
    .Y(_06062_));
 AOI211x1_ASAP7_75t_R _28505_ (.A1(_05890_),
    .A2(_06021_),
    .B(_06062_),
    .C(_05986_),
    .Y(_06063_));
 NOR2x1_ASAP7_75t_R _28506_ (.A(net5276),
    .B(net5616),
    .Y(_06064_));
 OAI21x1_ASAP7_75t_R _28507_ (.A1(net5621),
    .A2(net5618),
    .B(net6042),
    .Y(_06065_));
 NOR2x1_ASAP7_75t_R _28508_ (.A(_06064_),
    .B(_06065_),
    .Y(_06066_));
 NAND2x1_ASAP7_75t_R _28509_ (.A(net5623),
    .B(net5608),
    .Y(_06067_));
 AO21x1_ASAP7_75t_R _28510_ (.A1(_06067_),
    .A2(_05912_),
    .B(net5609),
    .Y(_06068_));
 OAI21x1_ASAP7_75t_R _28511_ (.A1(_06066_),
    .A2(_06068_),
    .B(net5355),
    .Y(_06069_));
 NOR2x1_ASAP7_75t_R _28512_ (.A(_06063_),
    .B(_06069_),
    .Y(_06070_));
 AO21x1_ASAP7_75t_R _28513_ (.A1(net6053),
    .A2(net6054),
    .B(_01353_),
    .Y(_06071_));
 AO21x1_ASAP7_75t_R _28514_ (.A1(_06071_),
    .A2(_05960_),
    .B(net6049),
    .Y(_06072_));
 NAND2x1_ASAP7_75t_R _28515_ (.A(net5611),
    .B(_06072_),
    .Y(_06073_));
 NOR2x1_ASAP7_75t_R _28516_ (.A(_06073_),
    .B(_06052_),
    .Y(_06074_));
 AO21x1_ASAP7_75t_R _28517_ (.A1(net4541),
    .A2(net6048),
    .B(net5611),
    .Y(_06075_));
 AOI21x1_ASAP7_75t_R _28518_ (.A1(net5362),
    .A2(net5352),
    .B(net6048),
    .Y(_06076_));
 OAI21x1_ASAP7_75t_R _28519_ (.A1(_06075_),
    .A2(_06076_),
    .B(net5606),
    .Y(_06077_));
 OAI21x1_ASAP7_75t_R _28520_ (.A1(_06074_),
    .A2(_06077_),
    .B(net6039),
    .Y(_06078_));
 NOR2x1_ASAP7_75t_R _28521_ (.A(_06070_),
    .B(_06078_),
    .Y(_06079_));
 INVx1_ASAP7_75t_R _28522_ (.A(_01358_),
    .Y(_06080_));
 NAND2x1_ASAP7_75t_R _28523_ (.A(net6046),
    .B(net5606),
    .Y(_06081_));
 OAI21x1_ASAP7_75t_R _28524_ (.A1(net5617),
    .A2(_05977_),
    .B(_05893_),
    .Y(_06082_));
 OAI21x1_ASAP7_75t_R _28525_ (.A1(_06080_),
    .A2(_06081_),
    .B(_06082_),
    .Y(_06083_));
 AO21x1_ASAP7_75t_R _28527_ (.A1(_06083_),
    .A2(net6045),
    .B(net6039),
    .Y(_06085_));
 INVx1_ASAP7_75t_R _28528_ (.A(net5364),
    .Y(_06086_));
 NOR2x1_ASAP7_75t_R _28529_ (.A(_06065_),
    .B(_06086_),
    .Y(_06087_));
 OAI21x1_ASAP7_75t_R _28530_ (.A1(net5616),
    .A2(net5628),
    .B(net6051),
    .Y(_06088_));
 OAI21x1_ASAP7_75t_R _28532_ (.A1(net4838),
    .A2(_06088_),
    .B(net5606),
    .Y(_06090_));
 OAI21x1_ASAP7_75t_R _28533_ (.A1(_06087_),
    .A2(_06090_),
    .B(net5609),
    .Y(_06091_));
 OAI21x1_ASAP7_75t_R _28534_ (.A1(net5607),
    .A2(net5624),
    .B(net5620),
    .Y(_06092_));
 NAND2x1_ASAP7_75t_R _28535_ (.A(net5353),
    .B(_06092_),
    .Y(_06093_));
 OAI21x1_ASAP7_75t_R _28536_ (.A1(_06064_),
    .A2(_05917_),
    .B(net5355),
    .Y(_06094_));
 AOI21x1_ASAP7_75t_R _28537_ (.A1(net6051),
    .A2(_06093_),
    .B(_06094_),
    .Y(_06095_));
 NOR2x1_ASAP7_75t_R _28538_ (.A(_06091_),
    .B(_06095_),
    .Y(_06096_));
 OAI21x1_ASAP7_75t_R _28539_ (.A1(_06085_),
    .A2(_06096_),
    .B(net6038),
    .Y(_06097_));
 OAI22x1_ASAP7_75t_R _28540_ (.A1(_06037_),
    .A2(_06061_),
    .B1(_06079_),
    .B2(_06097_),
    .Y(_00137_));
 AO21x1_ASAP7_75t_R _28541_ (.A1(net6057),
    .A2(net6058),
    .B(_01349_),
    .Y(_06098_));
 AO21x1_ASAP7_75t_R _28542_ (.A1(_05989_),
    .A2(_06098_),
    .B(net6049),
    .Y(_06099_));
 INVx1_ASAP7_75t_R _28543_ (.A(_05882_),
    .Y(_06100_));
 AO21x1_ASAP7_75t_R _28544_ (.A1(_05896_),
    .A2(_06100_),
    .B(net6041),
    .Y(_06101_));
 AO21x1_ASAP7_75t_R _28545_ (.A1(_06099_),
    .A2(_06101_),
    .B(net5613),
    .Y(_06102_));
 INVx1_ASAP7_75t_R _28546_ (.A(_06002_),
    .Y(_06103_));
 AOI21x1_ASAP7_75t_R _28547_ (.A1(net5623),
    .A2(net5607),
    .B(net6041),
    .Y(_06104_));
 AOI21x1_ASAP7_75t_R _28548_ (.A1(net6058),
    .A2(net6057),
    .B(_01353_),
    .Y(_06105_));
 OAI21x1_ASAP7_75t_R _28549_ (.A1(_06105_),
    .A2(_06065_),
    .B(net5614),
    .Y(_06106_));
 AO21x1_ASAP7_75t_R _28550_ (.A1(net4831),
    .A2(_06104_),
    .B(_06106_),
    .Y(_06107_));
 AOI21x1_ASAP7_75t_R _28551_ (.A1(_06102_),
    .A2(_06107_),
    .B(net5604),
    .Y(_06108_));
 AOI21x1_ASAP7_75t_R _28552_ (.A1(net5616),
    .A2(net5624),
    .B(net6041),
    .Y(_06109_));
 AOI22x1_ASAP7_75t_R _28553_ (.A1(_06109_),
    .A2(net5091),
    .B1(net5361),
    .B2(_05896_),
    .Y(_06110_));
 OAI21x1_ASAP7_75t_R _28555_ (.A1(net6045),
    .A2(_06110_),
    .B(net5604),
    .Y(_06112_));
 NAND2x1_ASAP7_75t_R _28556_ (.A(_06071_),
    .B(_06051_),
    .Y(_06113_));
 INVx1_ASAP7_75t_R _28557_ (.A(_05946_),
    .Y(_06114_));
 AOI211x1_ASAP7_75t_R _28558_ (.A1(_06113_),
    .A2(net6046),
    .B(_06114_),
    .C(net5613),
    .Y(_06115_));
 OAI21x1_ASAP7_75t_R _28559_ (.A1(_06112_),
    .A2(_06115_),
    .B(net5355),
    .Y(_06116_));
 NOR2x1_ASAP7_75t_R _28560_ (.A(_06108_),
    .B(_06116_),
    .Y(_06117_));
 OAI21x1_ASAP7_75t_R _28561_ (.A1(net5620),
    .A2(net5607),
    .B(net6041),
    .Y(_06118_));
 NOR2x1_ASAP7_75t_R _28562_ (.A(net4993),
    .B(_06118_),
    .Y(_06119_));
 NAND2x1_ASAP7_75t_R _28563_ (.A(net6049),
    .B(_06009_),
    .Y(_06120_));
 AOI21x1_ASAP7_75t_R _28564_ (.A1(net5617),
    .A2(net5630),
    .B(net5620),
    .Y(_06121_));
 OAI21x1_ASAP7_75t_R _28565_ (.A1(_06120_),
    .A2(_06121_),
    .B(net6045),
    .Y(_06122_));
 NOR2x1_ASAP7_75t_R _28566_ (.A(_06119_),
    .B(_06122_),
    .Y(_06123_));
 OAI21x1_ASAP7_75t_R _28567_ (.A1(net5616),
    .A2(net5617),
    .B(net5630),
    .Y(_06124_));
 NAND2x1_ASAP7_75t_R _28568_ (.A(net6049),
    .B(_06124_),
    .Y(_06125_));
 NOR2x1_ASAP7_75t_R _28569_ (.A(_05911_),
    .B(net6052),
    .Y(_06126_));
 AOI21x1_ASAP7_75t_R _28570_ (.A1(net5272),
    .A2(net5621),
    .B(net6045),
    .Y(_06127_));
 AOI21x1_ASAP7_75t_R _28571_ (.A1(_06126_),
    .A2(_06127_),
    .B(_05879_),
    .Y(_06128_));
 OAI21x1_ASAP7_75t_R _28572_ (.A1(net6045),
    .A2(_06125_),
    .B(_06128_),
    .Y(_06129_));
 NOR2x1_ASAP7_75t_R _28573_ (.A(_06123_),
    .B(_06129_),
    .Y(_06130_));
 NOR3x1_ASAP7_75t_R _28574_ (.A(net6046),
    .B(_06105_),
    .C(net5090),
    .Y(_06131_));
 NOR2x1_ASAP7_75t_R _28575_ (.A(_05990_),
    .B(_06120_),
    .Y(_06132_));
 OAI21x1_ASAP7_75t_R _28576_ (.A1(_06131_),
    .A2(_06132_),
    .B(net5613),
    .Y(_06133_));
 NAND2x1_ASAP7_75t_R _28577_ (.A(_06103_),
    .B(net5089),
    .Y(_06134_));
 AOI21x1_ASAP7_75t_R _28578_ (.A1(net6041),
    .A2(_06134_),
    .B(net5614),
    .Y(_06135_));
 AO21x1_ASAP7_75t_R _28579_ (.A1(_05977_),
    .A2(net5089),
    .B(net6041),
    .Y(_06136_));
 NAND2x1_ASAP7_75t_R _28580_ (.A(_06135_),
    .B(_06136_),
    .Y(_06137_));
 AOI21x1_ASAP7_75t_R _28581_ (.A1(_06133_),
    .A2(_06137_),
    .B(net5604),
    .Y(_06138_));
 OAI21x1_ASAP7_75t_R _28582_ (.A1(_06130_),
    .A2(_06138_),
    .B(net5605),
    .Y(_06139_));
 NAND2x1_ASAP7_75t_R _28583_ (.A(net6038),
    .B(_06139_),
    .Y(_06140_));
 AND2x2_ASAP7_75t_R _28584_ (.A(_01346_),
    .B(net5274),
    .Y(_06141_));
 AO21x1_ASAP7_75t_R _28585_ (.A1(net6053),
    .A2(net6054),
    .B(_06141_),
    .Y(_06142_));
 AOI21x1_ASAP7_75t_R _28586_ (.A1(net4828),
    .A2(_06051_),
    .B(net6041),
    .Y(_06143_));
 NAND2x1_ASAP7_75t_R _28587_ (.A(net5614),
    .B(_06082_),
    .Y(_06144_));
 NAND2x1p5_ASAP7_75t_R _28588_ (.A(_06006_),
    .B(_05957_),
    .Y(_06145_));
 NOR2x1_ASAP7_75t_R _28589_ (.A(net6046),
    .B(_06041_),
    .Y(_06146_));
 NOR2x1_ASAP7_75t_R _28590_ (.A(net5614),
    .B(_06146_),
    .Y(_06147_));
 AOI21x1_ASAP7_75t_R _28591_ (.A1(_06145_),
    .A2(_06147_),
    .B(net6039),
    .Y(_06148_));
 OAI21x1_ASAP7_75t_R _28592_ (.A1(_06143_),
    .A2(_06144_),
    .B(_06148_),
    .Y(_06149_));
 OA21x2_ASAP7_75t_R _28593_ (.A1(net6049),
    .A2(_01361_),
    .B(net6045),
    .Y(_06150_));
 OAI21x1_ASAP7_75t_R _28594_ (.A1(net5624),
    .A2(_05977_),
    .B(_06021_),
    .Y(_06151_));
 AOI21x1_ASAP7_75t_R _28595_ (.A1(_06150_),
    .A2(_06151_),
    .B(net5604),
    .Y(_06152_));
 NAND2x1_ASAP7_75t_R _28596_ (.A(_06104_),
    .B(_06045_),
    .Y(_06153_));
 AOI21x1_ASAP7_75t_R _28597_ (.A1(_05995_),
    .A2(_05994_),
    .B(net6045),
    .Y(_06154_));
 NAND2x1_ASAP7_75t_R _28598_ (.A(_06153_),
    .B(_06154_),
    .Y(_06155_));
 AOI21x1_ASAP7_75t_R _28599_ (.A1(_06152_),
    .A2(_06155_),
    .B(net5606),
    .Y(_06156_));
 AOI21x1_ASAP7_75t_R _28600_ (.A1(_06149_),
    .A2(_06156_),
    .B(net6038),
    .Y(_06157_));
 NOR2x1_ASAP7_75t_R _28601_ (.A(_01362_),
    .B(net6049),
    .Y(_06158_));
 AOI21x1_ASAP7_75t_R _28602_ (.A1(net5614),
    .A2(_06158_),
    .B(_05879_),
    .Y(_06159_));
 OAI21x1_ASAP7_75t_R _28603_ (.A1(net6045),
    .A2(_06125_),
    .B(_06159_),
    .Y(_06160_));
 NAND2x1_ASAP7_75t_R _28604_ (.A(_01360_),
    .B(net6049),
    .Y(_06161_));
 AOI21x1_ASAP7_75t_R _28605_ (.A1(_06161_),
    .A2(_05946_),
    .B(net5613),
    .Y(_06162_));
 NOR2x1_ASAP7_75t_R _28606_ (.A(_06160_),
    .B(_06162_),
    .Y(_06163_));
 NAND2x1_ASAP7_75t_R _28607_ (.A(_01358_),
    .B(net6041),
    .Y(_06164_));
 AOI21x1_ASAP7_75t_R _28608_ (.A1(net5616),
    .A2(net5627),
    .B(net6042),
    .Y(_06165_));
 AOI21x1_ASAP7_75t_R _28609_ (.A1(_05846_),
    .A2(_06165_),
    .B(_05839_),
    .Y(_06166_));
 NAND2x1_ASAP7_75t_R _28610_ (.A(_06164_),
    .B(_06166_),
    .Y(_06167_));
 NOR3x1_ASAP7_75t_R _28611_ (.A(_05828_),
    .B(net6041),
    .C(net4993),
    .Y(_06168_));
 NOR2x1_ASAP7_75t_R _28612_ (.A(_05825_),
    .B(_06118_),
    .Y(_06169_));
 OAI21x1_ASAP7_75t_R _28613_ (.A1(_06168_),
    .A2(_06169_),
    .B(net5612),
    .Y(_06170_));
 AOI21x1_ASAP7_75t_R _28614_ (.A1(_06167_),
    .A2(_06170_),
    .B(net5604),
    .Y(_06171_));
 OAI21x1_ASAP7_75t_R _28615_ (.A1(_06163_),
    .A2(_06171_),
    .B(net5605),
    .Y(_06172_));
 NAND2x1_ASAP7_75t_R _28616_ (.A(_06157_),
    .B(_06172_),
    .Y(_06173_));
 OAI21x1_ASAP7_75t_R _28617_ (.A1(_06117_),
    .A2(_06140_),
    .B(_06173_),
    .Y(_00138_));
 AO21x1_ASAP7_75t_R _28618_ (.A1(net6050),
    .A2(net4728),
    .B(net6045),
    .Y(_06174_));
 AO21x1_ASAP7_75t_R _28619_ (.A1(net5364),
    .A2(_05849_),
    .B(_06174_),
    .Y(_06175_));
 NAND2x1_ASAP7_75t_R _28620_ (.A(net5360),
    .B(_05849_),
    .Y(_06176_));
 NAND2x1_ASAP7_75t_R _28621_ (.A(net4541),
    .B(_06104_),
    .Y(_06177_));
 AO21x1_ASAP7_75t_R _28622_ (.A1(_06176_),
    .A2(_06177_),
    .B(net5611),
    .Y(_06178_));
 AOI21x1_ASAP7_75t_R _28623_ (.A1(_06175_),
    .A2(_06178_),
    .B(net5355),
    .Y(_06179_));
 INVx1_ASAP7_75t_R _28624_ (.A(net5362),
    .Y(_06180_));
 OAI21x1_ASAP7_75t_R _28625_ (.A1(_05828_),
    .A2(_06180_),
    .B(net6040),
    .Y(_06181_));
 AO21x1_ASAP7_75t_R _28626_ (.A1(_06041_),
    .A2(_06100_),
    .B(net6041),
    .Y(_06182_));
 AND3x1_ASAP7_75t_R _28627_ (.A(_06181_),
    .B(_05839_),
    .C(_06182_),
    .Y(_06183_));
 AND3x1_ASAP7_75t_R _28628_ (.A(net4834),
    .B(_05957_),
    .C(net6049),
    .Y(_06184_));
 AO21x1_ASAP7_75t_R _28629_ (.A1(net5361),
    .A2(_05896_),
    .B(net5614),
    .Y(_06185_));
 OAI21x1_ASAP7_75t_R _28630_ (.A1(_06184_),
    .A2(_06185_),
    .B(net5355),
    .Y(_06186_));
 OAI21x1_ASAP7_75t_R _28631_ (.A1(_06183_),
    .A2(_06186_),
    .B(net5604),
    .Y(_06187_));
 AOI21x1_ASAP7_75t_R _28632_ (.A1(_05967_),
    .A2(net5352),
    .B(_05839_),
    .Y(_06188_));
 NOR2x1_ASAP7_75t_R _28633_ (.A(net6041),
    .B(_05828_),
    .Y(_06189_));
 NAND2x1_ASAP7_75t_R _28634_ (.A(_06189_),
    .B(_06092_),
    .Y(_06190_));
 OAI21x1_ASAP7_75t_R _28635_ (.A1(net5093),
    .A2(net5616),
    .B(_05819_),
    .Y(_06191_));
 AOI22x1_ASAP7_75t_R _28636_ (.A1(_06188_),
    .A2(_06190_),
    .B1(_05858_),
    .B2(_06191_),
    .Y(_06192_));
 OA21x2_ASAP7_75t_R _28637_ (.A1(net6040),
    .A2(net5620),
    .B(net6045),
    .Y(_06193_));
 NAND2x1_ASAP7_75t_R _28638_ (.A(_05989_),
    .B(net5360),
    .Y(_06194_));
 AOI21x1_ASAP7_75t_R _28639_ (.A1(_06193_),
    .A2(_06194_),
    .B(net5355),
    .Y(_06195_));
 AO21x1_ASAP7_75t_R _28640_ (.A1(_05915_),
    .A2(_06098_),
    .B(net6050),
    .Y(_06196_));
 AOI21x1_ASAP7_75t_R _28641_ (.A1(_05944_),
    .A2(_05916_),
    .B(net6045),
    .Y(_06197_));
 NAND2x1_ASAP7_75t_R _28642_ (.A(_06197_),
    .B(_06196_),
    .Y(_06198_));
 AOI21x1_ASAP7_75t_R _28643_ (.A1(_06195_),
    .A2(_06198_),
    .B(net5604),
    .Y(_06199_));
 OAI21x1_ASAP7_75t_R _28644_ (.A1(net5605),
    .A2(_06192_),
    .B(_06199_),
    .Y(_06200_));
 OAI21x1_ASAP7_75t_R _28645_ (.A1(_06179_),
    .A2(_06187_),
    .B(_06200_),
    .Y(_06201_));
 NOR2x1_ASAP7_75t_R _28646_ (.A(net6041),
    .B(_06103_),
    .Y(_06202_));
 NOR2x1_ASAP7_75t_R _28647_ (.A(net5606),
    .B(_06202_),
    .Y(_06203_));
 NAND2x1_ASAP7_75t_R _28648_ (.A(_06203_),
    .B(_06099_),
    .Y(_06204_));
 INVx1_ASAP7_75t_R _28649_ (.A(_06105_),
    .Y(_06205_));
 AO21x1_ASAP7_75t_R _28650_ (.A1(net4829),
    .A2(_06205_),
    .B(net6041),
    .Y(_06206_));
 AOI21x1_ASAP7_75t_R _28651_ (.A1(_05915_),
    .A2(_05908_),
    .B(net5355),
    .Y(_06207_));
 NAND2x1_ASAP7_75t_R _28652_ (.A(_06206_),
    .B(_06207_),
    .Y(_06208_));
 NAND2x1_ASAP7_75t_R _28653_ (.A(_06204_),
    .B(_06208_),
    .Y(_06209_));
 NAND2x1_ASAP7_75t_R _28654_ (.A(_05977_),
    .B(_05893_),
    .Y(_06210_));
 AOI21x1_ASAP7_75t_R _28655_ (.A1(_05884_),
    .A2(_06210_),
    .B(net5355),
    .Y(_06211_));
 NAND2x1_ASAP7_75t_R _28656_ (.A(net4729),
    .B(net6041),
    .Y(_06212_));
 OAI21x1_ASAP7_75t_R _28657_ (.A1(net5605),
    .A2(_06212_),
    .B(_05973_),
    .Y(_06213_));
 OAI21x1_ASAP7_75t_R _28658_ (.A1(_06211_),
    .A2(_06213_),
    .B(net5604),
    .Y(_06214_));
 AOI21x1_ASAP7_75t_R _28659_ (.A1(net6045),
    .A2(_06209_),
    .B(_06214_),
    .Y(_06215_));
 NAND3x1_ASAP7_75t_R _28660_ (.A(net5617),
    .B(net6047),
    .C(net5623),
    .Y(_06216_));
 AOI21x1_ASAP7_75t_R _28661_ (.A1(net5090),
    .A2(net6047),
    .B(net6045),
    .Y(_06217_));
 OAI21x1_ASAP7_75t_R _28662_ (.A1(net4994),
    .A2(_06105_),
    .B(net6043),
    .Y(_06218_));
 NAND3x1_ASAP7_75t_R _28663_ (.A(_06216_),
    .B(_06217_),
    .C(_06218_),
    .Y(_06219_));
 NAND2x1_ASAP7_75t_R _28664_ (.A(_06032_),
    .B(_05963_),
    .Y(_06220_));
 AOI21x1_ASAP7_75t_R _28665_ (.A1(_06219_),
    .A2(_06220_),
    .B(net5605),
    .Y(_06221_));
 AO21x1_ASAP7_75t_R _28666_ (.A1(_06098_),
    .A2(_06142_),
    .B(net6041),
    .Y(_06222_));
 AOI21x1_ASAP7_75t_R _28667_ (.A1(_06222_),
    .A2(_06082_),
    .B(net5614),
    .Y(_06223_));
 NAND2x1_ASAP7_75t_R _28668_ (.A(net5605),
    .B(_06106_),
    .Y(_06224_));
 OAI21x1_ASAP7_75t_R _28669_ (.A1(_06223_),
    .A2(_06224_),
    .B(net6039),
    .Y(_06225_));
 NOR2x1_ASAP7_75t_R _28670_ (.A(_06221_),
    .B(_06225_),
    .Y(_06226_));
 OAI21x1_ASAP7_75t_R _28671_ (.A1(_06215_),
    .A2(_06226_),
    .B(net6038),
    .Y(_06227_));
 OAI21x1_ASAP7_75t_R _28672_ (.A1(net6038),
    .A2(_06201_),
    .B(_06227_),
    .Y(_00139_));
 NAND2x1_ASAP7_75t_R _28673_ (.A(_05824_),
    .B(_06165_),
    .Y(_06228_));
 NAND2x1_ASAP7_75t_R _28674_ (.A(net5360),
    .B(_05885_),
    .Y(_06229_));
 AOI21x1_ASAP7_75t_R _28675_ (.A1(_06228_),
    .A2(net5084),
    .B(net6045),
    .Y(_06230_));
 OA21x2_ASAP7_75t_R _28676_ (.A1(_06086_),
    .A2(_06065_),
    .B(_06166_),
    .Y(_06231_));
 OAI21x1_ASAP7_75t_R _28677_ (.A1(_06230_),
    .A2(_06231_),
    .B(net6039),
    .Y(_06232_));
 INVx1_ASAP7_75t_R _28678_ (.A(_06128_),
    .Y(_06233_));
 AOI21x1_ASAP7_75t_R _28679_ (.A1(net6045),
    .A2(_05959_),
    .B(_06233_),
    .Y(_06234_));
 AO21x1_ASAP7_75t_R _28680_ (.A1(_05981_),
    .A2(net5618),
    .B(net6045),
    .Y(_06235_));
 NAND2x1_ASAP7_75t_R _28681_ (.A(net6045),
    .B(_05890_),
    .Y(_06236_));
 AO21x1_ASAP7_75t_R _28682_ (.A1(_06235_),
    .A2(_06236_),
    .B(_06088_),
    .Y(_06237_));
 NAND2x1_ASAP7_75t_R _28683_ (.A(_06234_),
    .B(_06237_),
    .Y(_06238_));
 AOI21x1_ASAP7_75t_R _28684_ (.A1(_06232_),
    .A2(_06238_),
    .B(net5355),
    .Y(_06239_));
 OAI22x1_ASAP7_75t_R _28685_ (.A1(_05917_),
    .A2(_06064_),
    .B1(_06016_),
    .B2(_06044_),
    .Y(_06240_));
 NAND2x1_ASAP7_75t_R _28686_ (.A(net4837),
    .B(net5609),
    .Y(_06241_));
 OA21x2_ASAP7_75t_R _28687_ (.A1(net4833),
    .A2(_06241_),
    .B(net6039),
    .Y(_06242_));
 OAI21x1_ASAP7_75t_R _28688_ (.A1(net5609),
    .A2(_06240_),
    .B(_06242_),
    .Y(_06243_));
 NAND2x1_ASAP7_75t_R _28689_ (.A(net5355),
    .B(_06243_),
    .Y(_06244_));
 AOI21x1_ASAP7_75t_R _28690_ (.A1(net4833),
    .A2(_05982_),
    .B(net5610),
    .Y(_06245_));
 AO21x1_ASAP7_75t_R _28691_ (.A1(net5086),
    .A2(_05995_),
    .B(net6052),
    .Y(_06246_));
 NAND2x1_ASAP7_75t_R _28692_ (.A(_05966_),
    .B(net6052),
    .Y(_06247_));
 AND3x1_ASAP7_75t_R _28693_ (.A(_06005_),
    .B(_06217_),
    .C(_06247_),
    .Y(_06248_));
 AOI211x1_ASAP7_75t_R _28694_ (.A1(_06245_),
    .A2(_06246_),
    .B(_06248_),
    .C(net6039),
    .Y(_06249_));
 OAI21x1_ASAP7_75t_R _28695_ (.A1(_06244_),
    .A2(_06249_),
    .B(_06036_),
    .Y(_06250_));
 NAND2x1_ASAP7_75t_R _28696_ (.A(_05851_),
    .B(_05855_),
    .Y(_06251_));
 AOI21x1_ASAP7_75t_R _28697_ (.A1(_05999_),
    .A2(_06251_),
    .B(net5610),
    .Y(_06252_));
 NAND2x1_ASAP7_75t_R _28698_ (.A(_05989_),
    .B(_05984_),
    .Y(_06253_));
 AOI21x1_ASAP7_75t_R _28699_ (.A1(_06229_),
    .A2(_06253_),
    .B(net6045),
    .Y(_06254_));
 OAI21x1_ASAP7_75t_R _28700_ (.A1(_06252_),
    .A2(_06254_),
    .B(net5606),
    .Y(_06255_));
 OAI21x1_ASAP7_75t_R _28701_ (.A1(_01352_),
    .A2(net6052),
    .B(_06247_),
    .Y(_06256_));
 AOI21x1_ASAP7_75t_R _28702_ (.A1(net6045),
    .A2(_06256_),
    .B(net5606),
    .Y(_06257_));
 NAND2x1_ASAP7_75t_R _28703_ (.A(_05944_),
    .B(_05984_),
    .Y(_06258_));
 AOI21x1_ASAP7_75t_R _28704_ (.A1(_05989_),
    .A2(_05944_),
    .B(net6052),
    .Y(_06259_));
 NOR2x1_ASAP7_75t_R _28705_ (.A(net6045),
    .B(_06259_),
    .Y(_06260_));
 NAND2x1_ASAP7_75t_R _28706_ (.A(_06258_),
    .B(_06260_),
    .Y(_06261_));
 AOI21x1_ASAP7_75t_R _28707_ (.A1(_06257_),
    .A2(_06261_),
    .B(net6039),
    .Y(_06262_));
 NAND2x1_ASAP7_75t_R _28708_ (.A(_06255_),
    .B(_06262_),
    .Y(_06263_));
 AOI21x1_ASAP7_75t_R _28709_ (.A1(_06126_),
    .A2(_05995_),
    .B(net5609),
    .Y(_06264_));
 NAND2x1_ASAP7_75t_R _28710_ (.A(_05934_),
    .B(_06264_),
    .Y(_06265_));
 OAI21x1_ASAP7_75t_R _28711_ (.A1(net5618),
    .A2(net5364),
    .B(net6051),
    .Y(_06266_));
 OA21x2_ASAP7_75t_R _28712_ (.A1(net5092),
    .A2(net5616),
    .B(net6042),
    .Y(_06267_));
 NOR2x1_ASAP7_75t_R _28713_ (.A(net6045),
    .B(_06267_),
    .Y(_06268_));
 AOI21x1_ASAP7_75t_R _28714_ (.A1(_06266_),
    .A2(_06268_),
    .B(net5606),
    .Y(_06269_));
 NAND2x1_ASAP7_75t_R _28715_ (.A(_06269_),
    .B(_06265_),
    .Y(_06270_));
 NAND2x1_ASAP7_75t_R _28716_ (.A(_05890_),
    .B(net5364),
    .Y(_06271_));
 AOI21x1_ASAP7_75t_R _28717_ (.A1(_05912_),
    .A2(_06067_),
    .B(net6045),
    .Y(_06272_));
 OAI21x1_ASAP7_75t_R _28718_ (.A1(net6051),
    .A2(_06271_),
    .B(_06272_),
    .Y(_06273_));
 NOR2x1_ASAP7_75t_R _28719_ (.A(net5609),
    .B(_06030_),
    .Y(_06274_));
 NAND2x1_ASAP7_75t_R _28720_ (.A(_06056_),
    .B(_05849_),
    .Y(_06275_));
 AOI21x1_ASAP7_75t_R _28721_ (.A1(_06274_),
    .A2(_06275_),
    .B(net5355),
    .Y(_06276_));
 AOI21x1_ASAP7_75t_R _28722_ (.A1(_06273_),
    .A2(_06276_),
    .B(net5604),
    .Y(_06277_));
 AOI21x1_ASAP7_75t_R _28723_ (.A1(_06277_),
    .A2(_06270_),
    .B(_06036_),
    .Y(_06278_));
 NAND2x1_ASAP7_75t_R _28724_ (.A(_06278_),
    .B(_06263_),
    .Y(_06279_));
 OAI21x1_ASAP7_75t_R _28725_ (.A1(_06239_),
    .A2(_06250_),
    .B(_06279_),
    .Y(_00140_));
 OA21x2_ASAP7_75t_R _28726_ (.A1(net5617),
    .A2(net6043),
    .B(net6045),
    .Y(_06280_));
 AO21x1_ASAP7_75t_R _28727_ (.A1(_05850_),
    .A2(_06280_),
    .B(net5605),
    .Y(_06281_));
 AO21x1_ASAP7_75t_R _28728_ (.A1(_06086_),
    .A2(net5617),
    .B(_06038_),
    .Y(_06282_));
 OA21x2_ASAP7_75t_R _28729_ (.A1(_05983_),
    .A2(net5616),
    .B(net6042),
    .Y(_06283_));
 AOI21x1_ASAP7_75t_R _28730_ (.A1(net5356),
    .A2(_06283_),
    .B(net6045),
    .Y(_06284_));
 AND2x2_ASAP7_75t_R _28731_ (.A(_06282_),
    .B(_06284_),
    .Y(_06285_));
 OAI21x1_ASAP7_75t_R _28732_ (.A1(_06281_),
    .A2(_06285_),
    .B(net6039),
    .Y(_06286_));
 NOR2x1_ASAP7_75t_R _28733_ (.A(net6047),
    .B(_05958_),
    .Y(_06287_));
 NOR2x1_ASAP7_75t_R _28734_ (.A(_06287_),
    .B(_05935_),
    .Y(_06288_));
 AO21x1_ASAP7_75t_R _28735_ (.A1(_06054_),
    .A2(_06205_),
    .B(net6048),
    .Y(_06289_));
 AOI21x1_ASAP7_75t_R _28736_ (.A1(net6048),
    .A2(net4832),
    .B(net6045),
    .Y(_06290_));
 AO21x1_ASAP7_75t_R _28737_ (.A1(_06289_),
    .A2(_06290_),
    .B(net5355),
    .Y(_06291_));
 NOR2x1_ASAP7_75t_R _28738_ (.A(_06288_),
    .B(_06291_),
    .Y(_06292_));
 NAND2x1_ASAP7_75t_R _28739_ (.A(net5085),
    .B(net5616),
    .Y(_06293_));
 AO21x1_ASAP7_75t_R _28740_ (.A1(_06293_),
    .A2(net6052),
    .B(_05839_),
    .Y(_06294_));
 AOI21x1_ASAP7_75t_R _28741_ (.A1(net5352),
    .A2(_06092_),
    .B(net6050),
    .Y(_06295_));
 AOI21x1_ASAP7_75t_R _28742_ (.A1(_06057_),
    .A2(_06018_),
    .B(net5605),
    .Y(_06296_));
 OAI21x1_ASAP7_75t_R _28743_ (.A1(_06294_),
    .A2(_06295_),
    .B(_06296_),
    .Y(_06297_));
 OA21x2_ASAP7_75t_R _28744_ (.A1(net6040),
    .A2(_05826_),
    .B(net6045),
    .Y(_06298_));
 OAI21x1_ASAP7_75t_R _28745_ (.A1(net5607),
    .A2(_05989_),
    .B(net6040),
    .Y(_06299_));
 AOI21x1_ASAP7_75t_R _28746_ (.A1(_06298_),
    .A2(_06299_),
    .B(net5355),
    .Y(_06300_));
 OAI21x1_ASAP7_75t_R _28747_ (.A1(net4994),
    .A2(net4832),
    .B(net6050),
    .Y(_06301_));
 OAI21x1_ASAP7_75t_R _28748_ (.A1(net4729),
    .A2(_06105_),
    .B(_05853_),
    .Y(_06302_));
 NAND3x1_ASAP7_75t_R _28749_ (.A(_06301_),
    .B(_05839_),
    .C(_06302_),
    .Y(_06303_));
 AOI21x1_ASAP7_75t_R _28750_ (.A1(_06300_),
    .A2(_06303_),
    .B(net6039),
    .Y(_06304_));
 AOI21x1_ASAP7_75t_R _28751_ (.A1(_06297_),
    .A2(_06304_),
    .B(_06036_),
    .Y(_06305_));
 OAI21x1_ASAP7_75t_R _28752_ (.A1(_06286_),
    .A2(_06292_),
    .B(_06305_),
    .Y(_06306_));
 NOR2x1_ASAP7_75t_R _28753_ (.A(net6043),
    .B(net4832),
    .Y(_06307_));
 AOI22x1_ASAP7_75t_R _28754_ (.A1(_06307_),
    .A2(net5353),
    .B1(net5358),
    .B2(_05908_),
    .Y(_06308_));
 NAND2x1_ASAP7_75t_R _28755_ (.A(net5606),
    .B(_06247_),
    .Y(_06309_));
 AO21x1_ASAP7_75t_R _28756_ (.A1(net5354),
    .A2(_06267_),
    .B(_06309_),
    .Y(_06310_));
 OAI21x1_ASAP7_75t_R _28757_ (.A1(net5606),
    .A2(_06308_),
    .B(_06310_),
    .Y(_06311_));
 OAI21x1_ASAP7_75t_R _28758_ (.A1(net6052),
    .A2(_06105_),
    .B(net5606),
    .Y(_06312_));
 AOI211x1_ASAP7_75t_R _28759_ (.A1(net5620),
    .A2(net5276),
    .B(net4729),
    .C(net6041),
    .Y(_06313_));
 OAI21x1_ASAP7_75t_R _28760_ (.A1(_06312_),
    .A2(_06313_),
    .B(net6045),
    .Y(_06314_));
 AO21x1_ASAP7_75t_R _28761_ (.A1(net5607),
    .A2(net6050),
    .B(net5606),
    .Y(_06315_));
 AOI21x1_ASAP7_75t_R _28762_ (.A1(net5359),
    .A2(net5361),
    .B(_06315_),
    .Y(_06316_));
 OAI21x1_ASAP7_75t_R _28763_ (.A1(_06314_),
    .A2(_06316_),
    .B(net5604),
    .Y(_06317_));
 AOI21x1_ASAP7_75t_R _28764_ (.A1(net5611),
    .A2(_06311_),
    .B(_06317_),
    .Y(_06318_));
 AOI21x1_ASAP7_75t_R _28765_ (.A1(net5622),
    .A2(net5618),
    .B(net5090),
    .Y(_06319_));
 NOR2x1_ASAP7_75t_R _28766_ (.A(net6043),
    .B(_06319_),
    .Y(_06320_));
 AO21x1_ASAP7_75t_R _28767_ (.A1(net6043),
    .A2(_05915_),
    .B(net5611),
    .Y(_06321_));
 NOR2x1_ASAP7_75t_R _28768_ (.A(net6045),
    .B(_06126_),
    .Y(_06322_));
 AOI21x1_ASAP7_75t_R _28769_ (.A1(_06322_),
    .A2(_06031_),
    .B(net5355),
    .Y(_06323_));
 OAI21x1_ASAP7_75t_R _28770_ (.A1(_06320_),
    .A2(_06321_),
    .B(_06323_),
    .Y(_06324_));
 OAI21x1_ASAP7_75t_R _28771_ (.A1(net5625),
    .A2(_05977_),
    .B(_06283_),
    .Y(_06325_));
 INVx1_ASAP7_75t_R _28772_ (.A(_05928_),
    .Y(_06326_));
 NOR2x1_ASAP7_75t_R _28773_ (.A(net5273),
    .B(net6042),
    .Y(_06327_));
 AOI211x1_ASAP7_75t_R _28774_ (.A1(_06326_),
    .A2(net6052),
    .B(_06327_),
    .C(net6045),
    .Y(_06328_));
 NAND2x1_ASAP7_75t_R _28775_ (.A(_06325_),
    .B(_06328_),
    .Y(_06329_));
 NAND2x1_ASAP7_75t_R _28776_ (.A(_06027_),
    .B(_05916_),
    .Y(_06330_));
 AOI21x1_ASAP7_75t_R _28777_ (.A1(net6042),
    .A2(_05929_),
    .B(net5609),
    .Y(_06331_));
 AOI21x1_ASAP7_75t_R _28778_ (.A1(_06330_),
    .A2(_06331_),
    .B(net5606),
    .Y(_06332_));
 NAND2x1_ASAP7_75t_R _28779_ (.A(_06329_),
    .B(_06332_),
    .Y(_06333_));
 AOI21x1_ASAP7_75t_R _28780_ (.A1(_06324_),
    .A2(_06333_),
    .B(net5604),
    .Y(_06334_));
 OAI21x1_ASAP7_75t_R _28781_ (.A1(_06318_),
    .A2(_06334_),
    .B(_06036_),
    .Y(_06335_));
 NAND2x1_ASAP7_75t_R _28782_ (.A(_06335_),
    .B(_06306_),
    .Y(_00141_));
 OAI21x1_ASAP7_75t_R _28783_ (.A1(net6042),
    .A2(net4836),
    .B(net5606),
    .Y(_06336_));
 AOI21x1_ASAP7_75t_R _28784_ (.A1(_06071_),
    .A2(_06098_),
    .B(net6049),
    .Y(_06337_));
 AOI211x1_ASAP7_75t_R _28785_ (.A1(net5358),
    .A2(_06030_),
    .B(_06336_),
    .C(_06337_),
    .Y(_06338_));
 NAND2x1_ASAP7_75t_R _28786_ (.A(_01355_),
    .B(_01359_),
    .Y(_06339_));
 AO21x1_ASAP7_75t_R _28787_ (.A1(net6042),
    .A2(_06339_),
    .B(net5606),
    .Y(_06340_));
 NOR2x1_ASAP7_75t_R _28788_ (.A(_06088_),
    .B(_05919_),
    .Y(_06341_));
 OAI21x1_ASAP7_75t_R _28789_ (.A1(_06340_),
    .A2(_06341_),
    .B(net6045),
    .Y(_06342_));
 OAI21x1_ASAP7_75t_R _28790_ (.A1(_06338_),
    .A2(_06342_),
    .B(net6039),
    .Y(_06343_));
 OAI21x1_ASAP7_75t_R _28791_ (.A1(net4618),
    .A2(_06146_),
    .B(net5355),
    .Y(_06344_));
 AOI21x1_ASAP7_75t_R _28792_ (.A1(net5088),
    .A2(net4831),
    .B(_06081_),
    .Y(_06345_));
 INVx1_ASAP7_75t_R _28793_ (.A(_05967_),
    .Y(_06346_));
 NAND2x1_ASAP7_75t_R _28794_ (.A(net5606),
    .B(_05989_),
    .Y(_06347_));
 NAND2x1_ASAP7_75t_R _28795_ (.A(net6049),
    .B(_05961_),
    .Y(_06348_));
 OAI21x1_ASAP7_75t_R _28796_ (.A1(_06346_),
    .A2(_06347_),
    .B(_06348_),
    .Y(_06349_));
 NOR2x1_ASAP7_75t_R _28797_ (.A(_06345_),
    .B(_06349_),
    .Y(_06350_));
 AOI21x1_ASAP7_75t_R _28798_ (.A1(_06344_),
    .A2(_06350_),
    .B(net6045),
    .Y(_06351_));
 OAI21x1_ASAP7_75t_R _28799_ (.A1(_06343_),
    .A2(_06351_),
    .B(_06036_),
    .Y(_06352_));
 INVx1_ASAP7_75t_R _28800_ (.A(_06161_),
    .Y(_06353_));
 INVx1_ASAP7_75t_R _28801_ (.A(_05888_),
    .Y(_06354_));
 OAI21x1_ASAP7_75t_R _28802_ (.A1(_06353_),
    .A2(_06114_),
    .B(_06354_),
    .Y(_06355_));
 AOI21x1_ASAP7_75t_R _28803_ (.A1(net5354),
    .A2(_06092_),
    .B(net6043),
    .Y(_06356_));
 AOI21x1_ASAP7_75t_R _28804_ (.A1(net4994),
    .A2(net6043),
    .B(net5611),
    .Y(_06357_));
 OAI21x1_ASAP7_75t_R _28805_ (.A1(_06267_),
    .A2(_06356_),
    .B(_06357_),
    .Y(_06358_));
 AOI21x1_ASAP7_75t_R _28806_ (.A1(_06355_),
    .A2(_06358_),
    .B(net5605),
    .Y(_06359_));
 AO21x1_ASAP7_75t_R _28807_ (.A1(net4832),
    .A2(net6043),
    .B(net6045),
    .Y(_06360_));
 NOR2x1_ASAP7_75t_R _28808_ (.A(_06016_),
    .B(_05919_),
    .Y(_06361_));
 OAI21x1_ASAP7_75t_R _28809_ (.A1(_06360_),
    .A2(_06361_),
    .B(net5606),
    .Y(_06362_));
 AOI21x1_ASAP7_75t_R _28810_ (.A1(net4540),
    .A2(net4830),
    .B(net6047),
    .Y(_06363_));
 NAND2x1_ASAP7_75t_R _28811_ (.A(net5620),
    .B(net6049),
    .Y(_06364_));
 OAI21x1_ASAP7_75t_R _28812_ (.A1(net5624),
    .A2(_06364_),
    .B(net6045),
    .Y(_06365_));
 AOI211x1_ASAP7_75t_R _28813_ (.A1(net5362),
    .A2(_05855_),
    .B(_06363_),
    .C(_06365_),
    .Y(_06366_));
 OAI21x1_ASAP7_75t_R _28814_ (.A1(_06362_),
    .A2(_06366_),
    .B(net5604),
    .Y(_06367_));
 NOR2x1_ASAP7_75t_R _28815_ (.A(_06367_),
    .B(_06359_),
    .Y(_06368_));
 OA21x2_ASAP7_75t_R _28816_ (.A1(_06319_),
    .A2(net6043),
    .B(_06357_),
    .Y(_06369_));
 INVx1_ASAP7_75t_R _28817_ (.A(_06016_),
    .Y(_06370_));
 NOR2x1_ASAP7_75t_R _28818_ (.A(_06370_),
    .B(_05920_),
    .Y(_06371_));
 OAI21x1_ASAP7_75t_R _28819_ (.A1(_06369_),
    .A2(_06371_),
    .B(net6039),
    .Y(_06372_));
 AND2x2_ASAP7_75t_R _28820_ (.A(_06122_),
    .B(net5604),
    .Y(_06373_));
 INVx1_ASAP7_75t_R _28821_ (.A(_06258_),
    .Y(_06374_));
 OAI21x1_ASAP7_75t_R _28822_ (.A1(net4839),
    .A2(_06374_),
    .B(_05839_),
    .Y(_06375_));
 NAND2x1_ASAP7_75t_R _28823_ (.A(_06373_),
    .B(_06375_),
    .Y(_06376_));
 AOI21x1_ASAP7_75t_R _28824_ (.A1(_06372_),
    .A2(_06376_),
    .B(net5355),
    .Y(_06377_));
 AO21x1_ASAP7_75t_R _28825_ (.A1(net6052),
    .A2(_01356_),
    .B(net5609),
    .Y(_06378_));
 AOI21x1_ASAP7_75t_R _28826_ (.A1(net5356),
    .A2(_06283_),
    .B(_06378_),
    .Y(_06379_));
 NOR2x1_ASAP7_75t_R _28827_ (.A(net4994),
    .B(_06057_),
    .Y(_06380_));
 OAI21x1_ASAP7_75t_R _28828_ (.A1(_06062_),
    .A2(_06380_),
    .B(net5604),
    .Y(_06381_));
 OAI21x1_ASAP7_75t_R _28829_ (.A1(_06379_),
    .A2(_06381_),
    .B(net5355),
    .Y(_06382_));
 NAND2x1_ASAP7_75t_R _28830_ (.A(_05853_),
    .B(_05938_),
    .Y(_06383_));
 NOR2x1_ASAP7_75t_R _28831_ (.A(_06180_),
    .B(_06383_),
    .Y(_06384_));
 AOI21x1_ASAP7_75t_R _28832_ (.A1(_05989_),
    .A2(net5360),
    .B(net6040),
    .Y(_06385_));
 OAI21x1_ASAP7_75t_R _28833_ (.A1(_06384_),
    .A2(_06385_),
    .B(net5612),
    .Y(_06386_));
 AND2x2_ASAP7_75t_R _28834_ (.A(_06124_),
    .B(net6045),
    .Y(_06387_));
 INVx1_ASAP7_75t_R _28835_ (.A(_06385_),
    .Y(_06388_));
 NAND2x1_ASAP7_75t_R _28836_ (.A(_06387_),
    .B(_06388_),
    .Y(_06389_));
 AOI21x1_ASAP7_75t_R _28837_ (.A1(_06386_),
    .A2(_06389_),
    .B(net5604),
    .Y(_06390_));
 OAI21x1_ASAP7_75t_R _28838_ (.A1(_06382_),
    .A2(_06390_),
    .B(net6038),
    .Y(_06391_));
 OAI22x1_ASAP7_75t_R _28839_ (.A1(_06368_),
    .A2(_06352_),
    .B1(_06377_),
    .B2(_06391_),
    .Y(_00142_));
 INVx1_ASAP7_75t_R _28840_ (.A(_06267_),
    .Y(_06392_));
 AO21x1_ASAP7_75t_R _28841_ (.A1(_06392_),
    .A2(_06016_),
    .B(_06236_),
    .Y(_06393_));
 OAI21x1_ASAP7_75t_R _28842_ (.A1(_06049_),
    .A2(_06341_),
    .B(net5609),
    .Y(_06394_));
 AOI21x1_ASAP7_75t_R _28843_ (.A1(_06393_),
    .A2(_06394_),
    .B(net5355),
    .Y(_06395_));
 AND2x2_ASAP7_75t_R _28844_ (.A(_05994_),
    .B(net5358),
    .Y(_06396_));
 NAND2x1_ASAP7_75t_R _28845_ (.A(net5614),
    .B(_06222_),
    .Y(_06397_));
 OAI21x1_ASAP7_75t_R _28846_ (.A1(_06396_),
    .A2(_06397_),
    .B(net5355),
    .Y(_06398_));
 OR3x1_ASAP7_75t_R _28847_ (.A(net4832),
    .B(net6043),
    .C(_05810_),
    .Y(_06399_));
 OAI21x1_ASAP7_75t_R _28848_ (.A1(net5618),
    .A2(net5364),
    .B(_05890_),
    .Y(_06400_));
 NAND2x1_ASAP7_75t_R _28849_ (.A(net6043),
    .B(_06400_),
    .Y(_06401_));
 AOI21x1_ASAP7_75t_R _28850_ (.A1(_06399_),
    .A2(_06401_),
    .B(net5611),
    .Y(_06402_));
 OAI21x1_ASAP7_75t_R _28851_ (.A1(_06398_),
    .A2(_06402_),
    .B(net6039),
    .Y(_06403_));
 INVx1_ASAP7_75t_R _28852_ (.A(_06272_),
    .Y(_06404_));
 AND3x1_ASAP7_75t_R _28853_ (.A(_05918_),
    .B(net5364),
    .C(net6042),
    .Y(_06405_));
 AOI21x1_ASAP7_75t_R _28854_ (.A1(_01352_),
    .A2(net6052),
    .B(net5610),
    .Y(_06406_));
 AOI21x1_ASAP7_75t_R _28855_ (.A1(_05962_),
    .A2(_06406_),
    .B(net5606),
    .Y(_06407_));
 OAI21x1_ASAP7_75t_R _28856_ (.A1(_06404_),
    .A2(_06405_),
    .B(_06407_),
    .Y(_06408_));
 OA21x2_ASAP7_75t_R _28857_ (.A1(net6042),
    .A2(_01359_),
    .B(net6045),
    .Y(_06409_));
 AO21x1_ASAP7_75t_R _28858_ (.A1(_06100_),
    .A2(_06103_),
    .B(net6049),
    .Y(_06410_));
 AOI21x1_ASAP7_75t_R _28859_ (.A1(_06409_),
    .A2(_06410_),
    .B(net5355),
    .Y(_06411_));
 AO21x1_ASAP7_75t_R _28860_ (.A1(_05995_),
    .A2(_05915_),
    .B(net6043),
    .Y(_06412_));
 AOI21x1_ASAP7_75t_R _28861_ (.A1(_05944_),
    .A2(_05908_),
    .B(net6045),
    .Y(_06413_));
 NAND2x1_ASAP7_75t_R _28862_ (.A(_06412_),
    .B(_06413_),
    .Y(_06414_));
 AOI21x1_ASAP7_75t_R _28863_ (.A1(_06411_),
    .A2(_06414_),
    .B(net6039),
    .Y(_06415_));
 AOI21x1_ASAP7_75t_R _28864_ (.A1(_06408_),
    .A2(_06415_),
    .B(net6038),
    .Y(_06416_));
 OAI21x1_ASAP7_75t_R _28865_ (.A1(_06395_),
    .A2(_06403_),
    .B(_06416_),
    .Y(_06417_));
 AO21x1_ASAP7_75t_R _28866_ (.A1(_06045_),
    .A2(_06104_),
    .B(_06337_),
    .Y(_06418_));
 AOI21x1_ASAP7_75t_R _28867_ (.A1(net4834),
    .A2(_06021_),
    .B(net6045),
    .Y(_06419_));
 NAND2x1_ASAP7_75t_R _28868_ (.A(_05915_),
    .B(_05908_),
    .Y(_06420_));
 AOI21x1_ASAP7_75t_R _28869_ (.A1(_06419_),
    .A2(_06420_),
    .B(net5355),
    .Y(_06421_));
 OAI21x1_ASAP7_75t_R _28870_ (.A1(net5611),
    .A2(_06418_),
    .B(_06421_),
    .Y(_06422_));
 AND2x2_ASAP7_75t_R _28871_ (.A(_06383_),
    .B(net6045),
    .Y(_06423_));
 AOI21x1_ASAP7_75t_R _28872_ (.A1(_06258_),
    .A2(_06423_),
    .B(net5606),
    .Y(_06424_));
 NOR2x1_ASAP7_75t_R _28873_ (.A(_06062_),
    .B(_06259_),
    .Y(_06425_));
 OAI21x1_ASAP7_75t_R _28874_ (.A1(net6042),
    .A2(_06400_),
    .B(_06425_),
    .Y(_06426_));
 AOI21x1_ASAP7_75t_R _28875_ (.A1(_06424_),
    .A2(_06426_),
    .B(net5604),
    .Y(_06427_));
 NAND2x1_ASAP7_75t_R _28876_ (.A(_06422_),
    .B(_06427_),
    .Y(_06428_));
 AOI21x1_ASAP7_75t_R _28877_ (.A1(net6047),
    .A2(net5353),
    .B(_06321_),
    .Y(_06429_));
 OAI21x1_ASAP7_75t_R _28878_ (.A1(net5624),
    .A2(net5354),
    .B(net6047),
    .Y(_06430_));
 OAI21x1_ASAP7_75t_R _28879_ (.A1(net5618),
    .A2(net5364),
    .B(net6043),
    .Y(_06431_));
 AO21x1_ASAP7_75t_R _28880_ (.A1(net6043),
    .A2(net4994),
    .B(net6045),
    .Y(_06432_));
 AOI21x1_ASAP7_75t_R _28881_ (.A1(_06430_),
    .A2(_06431_),
    .B(_06432_),
    .Y(_06433_));
 OAI21x1_ASAP7_75t_R _28882_ (.A1(_06433_),
    .A2(_06429_),
    .B(net5606),
    .Y(_06434_));
 OAI21x1_ASAP7_75t_R _28883_ (.A1(_05945_),
    .A2(_06431_),
    .B(_06166_),
    .Y(_06435_));
 NAND2x1_ASAP7_75t_R _28884_ (.A(net6043),
    .B(net5618),
    .Y(_06436_));
 OAI21x1_ASAP7_75t_R _28885_ (.A1(_06044_),
    .A2(_06016_),
    .B(_06436_),
    .Y(_06437_));
 AOI21x1_ASAP7_75t_R _28886_ (.A1(net5611),
    .A2(_06437_),
    .B(net5606),
    .Y(_06438_));
 AOI21x1_ASAP7_75t_R _28887_ (.A1(_06435_),
    .A2(_06438_),
    .B(net6039),
    .Y(_06439_));
 AOI21x1_ASAP7_75t_R _28888_ (.A1(_06439_),
    .A2(_06434_),
    .B(_06036_),
    .Y(_06440_));
 NAND2x1_ASAP7_75t_R _28889_ (.A(_06440_),
    .B(_06428_),
    .Y(_06441_));
 NAND2x1_ASAP7_75t_R _28890_ (.A(_06417_),
    .B(_06441_),
    .Y(_00143_));
 NOR2x1_ASAP7_75t_R _28891_ (.A(net6657),
    .B(_00405_),
    .Y(_06442_));
 XOR2x2_ASAP7_75t_R _28892_ (.A(_12123_),
    .B(net6584),
    .Y(_06443_));
 XOR2x2_ASAP7_75t_R _28893_ (.A(_12160_),
    .B(_03665_),
    .Y(_06444_));
 NAND2x1_ASAP7_75t_R _28894_ (.A(_06443_),
    .B(_06444_),
    .Y(_06445_));
 XNOR2x2_ASAP7_75t_R _28895_ (.A(net6584),
    .B(_12123_),
    .Y(_06446_));
 XOR2x2_ASAP7_75t_R _28896_ (.A(_12162_),
    .B(_03665_),
    .Y(_06447_));
 NAND2x1_ASAP7_75t_R _28897_ (.A(_06446_),
    .B(_06447_),
    .Y(_06448_));
 AOI21x1_ASAP7_75t_R _28898_ (.A1(_06445_),
    .A2(_06448_),
    .B(net6454),
    .Y(_06449_));
 OAI21x1_ASAP7_75t_R _28899_ (.A1(net6392),
    .A2(_06449_),
    .B(net6487),
    .Y(_06450_));
 AND2x2_ASAP7_75t_R _28900_ (.A(net6454),
    .B(_00405_),
    .Y(_06451_));
 NAND2x1_ASAP7_75t_R _28901_ (.A(_06443_),
    .B(_06447_),
    .Y(_06452_));
 NAND2x1_ASAP7_75t_R _28902_ (.A(_06444_),
    .B(_06446_),
    .Y(_06453_));
 AOI21x1_ASAP7_75t_R _28903_ (.A1(_06452_),
    .A2(_06453_),
    .B(net6454),
    .Y(_06454_));
 INVx1_ASAP7_75t_R _28904_ (.A(net6487),
    .Y(_06455_));
 OAI21x1_ASAP7_75t_R _28905_ (.A1(_06451_),
    .A2(net6343),
    .B(_06455_),
    .Y(_06456_));
 NAND2x2_ASAP7_75t_R _28906_ (.A(_06450_),
    .B(_06456_),
    .Y(_06457_));
 OR2x2_ASAP7_75t_R _28908_ (.A(net6660),
    .B(_00406_),
    .Y(_06458_));
 NOR2x1_ASAP7_75t_R _28909_ (.A(_12319_),
    .B(_12145_),
    .Y(_06459_));
 NOR2x1p5_ASAP7_75t_R _28910_ (.A(net6549),
    .B(_12146_),
    .Y(_06460_));
 OAI21x1_ASAP7_75t_R _28911_ (.A1(_06460_),
    .A2(_06459_),
    .B(net6438),
    .Y(_06461_));
 INVx1_ASAP7_75t_R _28912_ (.A(_06461_),
    .Y(_06462_));
 NOR3x1_ASAP7_75t_R _28913_ (.A(_06460_),
    .B(_06459_),
    .C(net6438),
    .Y(_06463_));
 OAI21x1_ASAP7_75t_R _28914_ (.A1(_06463_),
    .A2(_06462_),
    .B(net6657),
    .Y(_06464_));
 AOI21x1_ASAP7_75t_R _28915_ (.A1(net6391),
    .A2(net5601),
    .B(net6492),
    .Y(_06465_));
 NAND2x1_ASAP7_75t_R _28916_ (.A(_00406_),
    .B(net6459),
    .Y(_06466_));
 XOR2x2_ASAP7_75t_R _28917_ (.A(_12145_),
    .B(_12319_),
    .Y(_06467_));
 NAND2x1_ASAP7_75t_R _28918_ (.A(net6435),
    .B(_06467_),
    .Y(_06468_));
 NAND3x1_ASAP7_75t_R _28919_ (.A(_06468_),
    .B(net6657),
    .C(_06461_),
    .Y(_06469_));
 INVx1_ASAP7_75t_R _28920_ (.A(net6492),
    .Y(_06470_));
 AOI21x1_ASAP7_75t_R _28921_ (.A1(_06466_),
    .A2(net6037),
    .B(_06470_),
    .Y(_06471_));
 NOR2x1_ASAP7_75t_R _28922_ (.A(_06465_),
    .B(_06471_),
    .Y(_06472_));
 XOR2x2_ASAP7_75t_R _28924_ (.A(net6635),
    .B(net6583),
    .Y(_06473_));
 NAND2x1_ASAP7_75t_R _28925_ (.A(net6436),
    .B(_06473_),
    .Y(_06474_));
 XNOR2x2_ASAP7_75t_R _28926_ (.A(net6635),
    .B(net6583),
    .Y(_06475_));
 NAND2x1_ASAP7_75t_R _28927_ (.A(net6552),
    .B(_06475_),
    .Y(_06476_));
 AOI21x1_ASAP7_75t_R _28928_ (.A1(_06474_),
    .A2(_06476_),
    .B(_03708_),
    .Y(_06477_));
 XOR2x2_ASAP7_75t_R _28929_ (.A(net6583),
    .B(net6552),
    .Y(_06478_));
 NAND2x1_ASAP7_75t_R _28930_ (.A(net6635),
    .B(_06478_),
    .Y(_06479_));
 XNOR2x2_ASAP7_75t_R _28931_ (.A(net6582),
    .B(net6552),
    .Y(_06480_));
 NAND2x1_ASAP7_75t_R _28932_ (.A(net6413),
    .B(_06480_),
    .Y(_06481_));
 AOI21x1_ASAP7_75t_R _28933_ (.A1(_06479_),
    .A2(_06481_),
    .B(_03697_),
    .Y(_06482_));
 OAI21x1_ASAP7_75t_R _28934_ (.A1(_06477_),
    .A2(_06482_),
    .B(net6656),
    .Y(_06483_));
 NOR2x1_ASAP7_75t_R _28935_ (.A(net6657),
    .B(_00407_),
    .Y(_06484_));
 INVx1_ASAP7_75t_R _28936_ (.A(_06484_),
    .Y(_06485_));
 NAND3x1_ASAP7_75t_R _28937_ (.A(_06483_),
    .B(net6480),
    .C(_06485_),
    .Y(_06486_));
 AO21x1_ASAP7_75t_R _28938_ (.A1(_06483_),
    .A2(_06485_),
    .B(net6480),
    .Y(_06487_));
 NAND2x1_ASAP7_75t_R _28940_ (.A(_06486_),
    .B(_06487_),
    .Y(_06489_));
 AOI21x1_ASAP7_75t_R _28942_ (.A1(_06464_),
    .A2(_06458_),
    .B(_06470_),
    .Y(_06490_));
 AOI21x1_ASAP7_75t_R _28943_ (.A1(_06466_),
    .A2(_06469_),
    .B(net6492),
    .Y(_06491_));
 NOR2x2_ASAP7_75t_R _28944_ (.A(_06491_),
    .B(_06490_),
    .Y(_06492_));
 NAND3x1_ASAP7_75t_R _28946_ (.A(_06483_),
    .B(_08822_),
    .C(_06485_),
    .Y(_06493_));
 AO21x1_ASAP7_75t_R _28947_ (.A1(_06483_),
    .A2(_06485_),
    .B(_08822_),
    .Y(_06494_));
 NAND2x2_ASAP7_75t_R _28949_ (.A(_06493_),
    .B(_06494_),
    .Y(_06496_));
 XOR2x2_ASAP7_75t_R _28951_ (.A(net6632),
    .B(_00597_),
    .Y(_06497_));
 XOR2x2_ASAP7_75t_R _28952_ (.A(_06497_),
    .B(_00692_),
    .Y(_06498_));
 XOR2x2_ASAP7_75t_R _28953_ (.A(_06498_),
    .B(_12270_),
    .Y(_06499_));
 NOR2x1_ASAP7_75t_R _28954_ (.A(net6657),
    .B(_00531_),
    .Y(_06500_));
 AO21x1_ASAP7_75t_R _28955_ (.A1(_06499_),
    .A2(net6657),
    .B(_06500_),
    .Y(_06501_));
 XOR2x2_ASAP7_75t_R _28956_ (.A(_06501_),
    .B(_00930_),
    .Y(_06502_));
 AO21x1_ASAP7_75t_R _28958_ (.A1(net6033),
    .A2(net6034),
    .B(_01365_),
    .Y(_06504_));
 INVx1_ASAP7_75t_R _28959_ (.A(_01369_),
    .Y(_06505_));
 XNOR2x2_ASAP7_75t_R _28961_ (.A(_00658_),
    .B(_12189_),
    .Y(_06507_));
 NOR2x1_ASAP7_75t_R _28962_ (.A(_06507_),
    .B(_03725_),
    .Y(_06508_));
 XOR2x2_ASAP7_75t_R _28963_ (.A(_12189_),
    .B(_00658_),
    .Y(_06509_));
 XNOR2x2_ASAP7_75t_R _28964_ (.A(_03724_),
    .B(_03723_),
    .Y(_06510_));
 OAI21x1_ASAP7_75t_R _28965_ (.A1(_06509_),
    .A2(_06510_),
    .B(net6657),
    .Y(_06511_));
 NAND2x1_ASAP7_75t_R _28966_ (.A(_00534_),
    .B(net6459),
    .Y(_06512_));
 OAI21x1_ASAP7_75t_R _28967_ (.A1(_06508_),
    .A2(_06511_),
    .B(_06512_),
    .Y(_06513_));
 XOR2x2_ASAP7_75t_R _28968_ (.A(_06513_),
    .B(_00927_),
    .Y(_06514_));
 AOI21x1_ASAP7_75t_R _28969_ (.A1(_06505_),
    .A2(net5600),
    .B(net6025),
    .Y(_06515_));
 NAND2x1_ASAP7_75t_R _28970_ (.A(_06504_),
    .B(net4492),
    .Y(_06516_));
 INVx1_ASAP7_75t_R _28971_ (.A(_01365_),
    .Y(_06517_));
 AO21x1_ASAP7_75t_R _28972_ (.A1(net6035),
    .A2(net6036),
    .B(_06517_),
    .Y(_06518_));
 AO21x1_ASAP7_75t_R _28974_ (.A1(net6033),
    .A2(net6034),
    .B(net4720),
    .Y(_06520_));
 XNOR2x2_ASAP7_75t_R _28976_ (.A(_00927_),
    .B(_06513_),
    .Y(_06522_));
 AO21x1_ASAP7_75t_R _28978_ (.A1(_06518_),
    .A2(net4539),
    .B(net6019),
    .Y(_06524_));
 XOR2x2_ASAP7_75t_R _28979_ (.A(_12215_),
    .B(_00659_),
    .Y(_06525_));
 XOR2x2_ASAP7_75t_R _28980_ (.A(_03748_),
    .B(_06525_),
    .Y(_06526_));
 NOR2x1_ASAP7_75t_R _28981_ (.A(net6659),
    .B(_00533_),
    .Y(_06527_));
 AOI21x1_ASAP7_75t_R _28982_ (.A1(net6659),
    .A2(_06526_),
    .B(_06527_),
    .Y(_06528_));
 XOR2x2_ASAP7_75t_R _28983_ (.A(_06528_),
    .B(_00928_),
    .Y(_06529_));
 AOI21x1_ASAP7_75t_R _28985_ (.A1(_06516_),
    .A2(_06524_),
    .B(net6016),
    .Y(_06531_));
 OAI21x1_ASAP7_75t_R _28986_ (.A1(net4720),
    .A2(net5600),
    .B(net6023),
    .Y(_06532_));
 INVx1_ASAP7_75t_R _28987_ (.A(net4537),
    .Y(_06533_));
 NAND2x1_ASAP7_75t_R _28988_ (.A(net5600),
    .B(net5602),
    .Y(_06534_));
 INVx1_ASAP7_75t_R _28989_ (.A(_01366_),
    .Y(_06535_));
 AOI21x1_ASAP7_75t_R _28990_ (.A1(net6036),
    .A2(net6035),
    .B(_06535_),
    .Y(_06536_));
 NOR2x2_ASAP7_75t_R _28991_ (.A(_06536_),
    .B(net6024),
    .Y(_06537_));
 INVx2_ASAP7_75t_R _28992_ (.A(_06529_),
    .Y(_06538_));
 AOI211x1_ASAP7_75t_R _28994_ (.A1(_06533_),
    .A2(net5351),
    .B(net5594),
    .C(_06537_),
    .Y(_06540_));
 NOR2x1_ASAP7_75t_R _28995_ (.A(net6659),
    .B(_00532_),
    .Y(_06541_));
 INVx1_ASAP7_75t_R _28996_ (.A(_06541_),
    .Y(_06542_));
 XOR2x2_ASAP7_75t_R _28997_ (.A(_00595_),
    .B(_00596_),
    .Y(_06543_));
 XOR2x2_ASAP7_75t_R _28998_ (.A(_06543_),
    .B(_15009_),
    .Y(_06544_));
 XOR2x2_ASAP7_75t_R _28999_ (.A(_06544_),
    .B(_12238_),
    .Y(_06545_));
 NAND2x1_ASAP7_75t_R _29000_ (.A(net6659),
    .B(_06545_),
    .Y(_06546_));
 AOI21x1_ASAP7_75t_R _29001_ (.A1(_06542_),
    .A2(_06546_),
    .B(_00929_),
    .Y(_06547_));
 INVx1_ASAP7_75t_R _29002_ (.A(_00929_),
    .Y(_06548_));
 AOI211x1_ASAP7_75t_R _29003_ (.A1(_06545_),
    .A2(net6659),
    .B(_06541_),
    .C(_06548_),
    .Y(_06549_));
 NOR2x1_ASAP7_75t_R _29004_ (.A(_06547_),
    .B(_06549_),
    .Y(_06550_));
 INVx1_ASAP7_75t_R _29005_ (.A(_06550_),
    .Y(_06551_));
 OAI21x1_ASAP7_75t_R _29007_ (.A1(_06531_),
    .A2(_06540_),
    .B(net5350),
    .Y(_06553_));
 NAND2x1_ASAP7_75t_R _29008_ (.A(net6032),
    .B(_06553_),
    .Y(_06554_));
 NOR2x1_ASAP7_75t_R _29009_ (.A(_06505_),
    .B(net5600),
    .Y(_06555_));
 INVx1_ASAP7_75t_R _29010_ (.A(_06555_),
    .Y(_06556_));
 AOI21x1_ASAP7_75t_R _29012_ (.A1(_06518_),
    .A2(_06556_),
    .B(net6019),
    .Y(_06558_));
 AO21x1_ASAP7_75t_R _29014_ (.A1(net5082),
    .A2(net5602),
    .B(net5595),
    .Y(_06560_));
 AOI21x1_ASAP7_75t_R _29017_ (.A1(net4539),
    .A2(_06560_),
    .B(net6028),
    .Y(_06563_));
 OAI21x1_ASAP7_75t_R _29020_ (.A1(_06558_),
    .A2(_06563_),
    .B(net5594),
    .Y(_06566_));
 NAND2x1_ASAP7_75t_R _29021_ (.A(net5600),
    .B(net5083),
    .Y(_06567_));
 NAND2x1_ASAP7_75t_R _29022_ (.A(net5602),
    .B(net5079),
    .Y(_06568_));
 AO21x1_ASAP7_75t_R _29025_ (.A1(net4827),
    .A2(net4826),
    .B(net6027),
    .Y(_06571_));
 NOR2x1_ASAP7_75t_R _29026_ (.A(net5603),
    .B(net5083),
    .Y(_06572_));
 NOR2x1_ASAP7_75t_R _29027_ (.A(net5600),
    .B(net5079),
    .Y(_06573_));
 OAI21x1_ASAP7_75t_R _29029_ (.A1(_06572_),
    .A2(_06573_),
    .B(net6025),
    .Y(_06575_));
 AO21x1_ASAP7_75t_R _29031_ (.A1(_06571_),
    .A2(_06575_),
    .B(net5594),
    .Y(_06577_));
 AOI21x1_ASAP7_75t_R _29032_ (.A1(_06566_),
    .A2(_06577_),
    .B(net5350),
    .Y(_06578_));
 NOR2x1_ASAP7_75t_R _29033_ (.A(_06578_),
    .B(_06554_),
    .Y(_06579_));
 OAI21x1_ASAP7_75t_R _29034_ (.A1(_06442_),
    .A2(_06449_),
    .B(_06455_),
    .Y(_06580_));
 OAI21x1_ASAP7_75t_R _29035_ (.A1(_06451_),
    .A2(_06454_),
    .B(net6487),
    .Y(_06581_));
 NAND2x1_ASAP7_75t_R _29036_ (.A(_06580_),
    .B(_06581_),
    .Y(_06582_));
 NAND2x1_ASAP7_75t_R _29038_ (.A(net5600),
    .B(net5590),
    .Y(_06583_));
 AO21x1_ASAP7_75t_R _29039_ (.A1(net6033),
    .A2(net6034),
    .B(net4798),
    .Y(_06584_));
 AO21x1_ASAP7_75t_R _29041_ (.A1(net5347),
    .A2(net4617),
    .B(net6027),
    .Y(_06586_));
 NAND2x1_ASAP7_75t_R _29042_ (.A(net5603),
    .B(net5083),
    .Y(_06587_));
 AOI21x1_ASAP7_75t_R _29043_ (.A1(net5600),
    .A2(net5079),
    .B(net6021),
    .Y(_06588_));
 OAI21x1_ASAP7_75t_R _29044_ (.A1(net5600),
    .A2(_06587_),
    .B(_06588_),
    .Y(_06589_));
 AO21x1_ASAP7_75t_R _29047_ (.A1(_06586_),
    .A2(_06589_),
    .B(net6017),
    .Y(_06592_));
 OA21x2_ASAP7_75t_R _29049_ (.A1(net5603),
    .A2(net5600),
    .B(net6018),
    .Y(_06594_));
 NOR2x1_ASAP7_75t_R _29050_ (.A(net5599),
    .B(net5590),
    .Y(_06595_));
 NAND2x1_ASAP7_75t_R _29051_ (.A(net5079),
    .B(_06595_),
    .Y(_06596_));
 NAND2x1_ASAP7_75t_R _29052_ (.A(_06594_),
    .B(_06596_),
    .Y(_06597_));
 INVx1_ASAP7_75t_R _29053_ (.A(_01374_),
    .Y(_06598_));
 AO21x1_ASAP7_75t_R _29054_ (.A1(net6033),
    .A2(net6034),
    .B(_06598_),
    .Y(_06599_));
 NAND2x1_ASAP7_75t_R _29056_ (.A(net4491),
    .B(_06588_),
    .Y(_06601_));
 AO21x1_ASAP7_75t_R _29057_ (.A1(_06597_),
    .A2(_06601_),
    .B(net5594),
    .Y(_06602_));
 AOI21x1_ASAP7_75t_R _29060_ (.A1(_06592_),
    .A2(_06602_),
    .B(net5591),
    .Y(_06605_));
 AO21x1_ASAP7_75t_R _29061_ (.A1(net6035),
    .A2(net6036),
    .B(net4793),
    .Y(_06606_));
 AO21x1_ASAP7_75t_R _29064_ (.A1(net4538),
    .A2(_06606_),
    .B(net6023),
    .Y(_06609_));
 OAI21x1_ASAP7_75t_R _29066_ (.A1(net5602),
    .A2(net5595),
    .B(net5079),
    .Y(_06611_));
 NAND2x1_ASAP7_75t_R _29067_ (.A(net6023),
    .B(_06611_),
    .Y(_06612_));
 AND3x1_ASAP7_75t_R _29068_ (.A(_06609_),
    .B(_06612_),
    .C(net6015),
    .Y(_06613_));
 INVx1_ASAP7_75t_R _29069_ (.A(net4794),
    .Y(_06614_));
 OA21x2_ASAP7_75t_R _29070_ (.A1(net5600),
    .A2(_06614_),
    .B(net6031),
    .Y(_06615_));
 NAND2x1_ASAP7_75t_R _29071_ (.A(_06615_),
    .B(_06596_),
    .Y(_06616_));
 AOI21x1_ASAP7_75t_R _29073_ (.A1(net5600),
    .A2(net5079),
    .B(net6031),
    .Y(_06618_));
 NOR2x1_ASAP7_75t_R _29074_ (.A(net6017),
    .B(net4823),
    .Y(_06619_));
 AO21x1_ASAP7_75t_R _29076_ (.A1(_06616_),
    .A2(_06619_),
    .B(net5348),
    .Y(_06621_));
 INVx1_ASAP7_75t_R _29077_ (.A(_06502_),
    .Y(_06622_));
 OAI21x1_ASAP7_75t_R _29079_ (.A1(_06613_),
    .A2(_06621_),
    .B(net5588),
    .Y(_06624_));
 XOR2x2_ASAP7_75t_R _29080_ (.A(_00597_),
    .B(net6630),
    .Y(_06625_));
 XOR2x2_ASAP7_75t_R _29081_ (.A(_06625_),
    .B(_00693_),
    .Y(_06626_));
 XOR2x2_ASAP7_75t_R _29082_ (.A(_06626_),
    .B(_12321_),
    .Y(_06627_));
 NOR2x1_ASAP7_75t_R _29083_ (.A(net6659),
    .B(_00530_),
    .Y(_06628_));
 AO21x1_ASAP7_75t_R _29084_ (.A1(_06627_),
    .A2(net6659),
    .B(_06628_),
    .Y(_06629_));
 XOR2x2_ASAP7_75t_R _29085_ (.A(_06629_),
    .B(_00931_),
    .Y(_06630_));
 OAI21x1_ASAP7_75t_R _29086_ (.A1(_06605_),
    .A2(_06624_),
    .B(net6014),
    .Y(_06631_));
 NAND2x1_ASAP7_75t_R _29087_ (.A(net5597),
    .B(net5602),
    .Y(_06632_));
 NOR2x1_ASAP7_75t_R _29088_ (.A(net5083),
    .B(net5343),
    .Y(_06633_));
 AOI21x1_ASAP7_75t_R _29089_ (.A1(net4796),
    .A2(net5600),
    .B(net6023),
    .Y(_06634_));
 INVx1_ASAP7_75t_R _29090_ (.A(_06634_),
    .Y(_06635_));
 OA21x2_ASAP7_75t_R _29093_ (.A1(net4617),
    .A2(net6031),
    .B(net5592),
    .Y(_06638_));
 OAI21x1_ASAP7_75t_R _29094_ (.A1(_06633_),
    .A2(_06635_),
    .B(_06638_),
    .Y(_06639_));
 INVx1_ASAP7_75t_R _29095_ (.A(_06584_),
    .Y(_06640_));
 AOI21x1_ASAP7_75t_R _29096_ (.A1(net6029),
    .A2(_06640_),
    .B(net5592),
    .Y(_06641_));
 OAI21x1_ASAP7_75t_R _29097_ (.A1(net5083),
    .A2(net5344),
    .B(_06515_),
    .Y(_06642_));
 AOI21x1_ASAP7_75t_R _29098_ (.A1(_06641_),
    .A2(_06642_),
    .B(net5350),
    .Y(_06643_));
 AOI21x1_ASAP7_75t_R _29099_ (.A1(_06639_),
    .A2(_06643_),
    .B(net5588),
    .Y(_06644_));
 AOI21x1_ASAP7_75t_R _29100_ (.A1(net6036),
    .A2(net6035),
    .B(net4795),
    .Y(_06645_));
 AOI21x1_ASAP7_75t_R _29101_ (.A1(net5596),
    .A2(net4826),
    .B(net4612),
    .Y(_06646_));
 NOR2x1_ASAP7_75t_R _29102_ (.A(net6029),
    .B(_06646_),
    .Y(_06647_));
 AO21x1_ASAP7_75t_R _29103_ (.A1(net6035),
    .A2(net6036),
    .B(net4798),
    .Y(_06648_));
 OA21x2_ASAP7_75t_R _29104_ (.A1(_06648_),
    .A2(net6029),
    .B(net5592),
    .Y(_06649_));
 NAND2x1_ASAP7_75t_R _29105_ (.A(_06504_),
    .B(_06588_),
    .Y(_06650_));
 NAND2x1_ASAP7_75t_R _29106_ (.A(_06649_),
    .B(_06650_),
    .Y(_06651_));
 INVx1_ASAP7_75t_R _29107_ (.A(_01382_),
    .Y(_06652_));
 AO21x1_ASAP7_75t_R _29109_ (.A1(net6035),
    .A2(net6036),
    .B(net4720),
    .Y(_06654_));
 NAND2x1p5_ASAP7_75t_R _29111_ (.A(_06654_),
    .B(net6021),
    .Y(_06656_));
 OAI21x1_ASAP7_75t_R _29112_ (.A1(_06652_),
    .A2(net6021),
    .B(_06656_),
    .Y(_06657_));
 AOI21x1_ASAP7_75t_R _29114_ (.A1(net6017),
    .A2(_06657_),
    .B(net5591),
    .Y(_06659_));
 OAI21x1_ASAP7_75t_R _29115_ (.A1(_06647_),
    .A2(_06651_),
    .B(_06659_),
    .Y(_06660_));
 AOI21x1_ASAP7_75t_R _29116_ (.A1(_06644_),
    .A2(_06660_),
    .B(net6014),
    .Y(_06661_));
 AO21x1_ASAP7_75t_R _29117_ (.A1(net6033),
    .A2(net6034),
    .B(_06535_),
    .Y(_06662_));
 NAND2x1p5_ASAP7_75t_R _29119_ (.A(net6026),
    .B(net4451),
    .Y(_06664_));
 INVx2_ASAP7_75t_R _29120_ (.A(_06664_),
    .Y(_06665_));
 AOI21x1_ASAP7_75t_R _29121_ (.A1(net6034),
    .A2(net6033),
    .B(_01370_),
    .Y(_06666_));
 OAI21x1_ASAP7_75t_R _29123_ (.A1(net4612),
    .A2(net4610),
    .B(net6022),
    .Y(_06668_));
 NAND2x1_ASAP7_75t_R _29124_ (.A(net6016),
    .B(_06668_),
    .Y(_06669_));
 INVx2_ASAP7_75t_R _29125_ (.A(_06645_),
    .Y(_06670_));
 OA21x2_ASAP7_75t_R _29126_ (.A1(_06670_),
    .A2(net6027),
    .B(net5594),
    .Y(_06671_));
 AOI21x1_ASAP7_75t_R _29127_ (.A1(_06671_),
    .A2(_06589_),
    .B(net5591),
    .Y(_06672_));
 OAI21x1_ASAP7_75t_R _29128_ (.A1(net4424),
    .A2(_06669_),
    .B(_06672_),
    .Y(_06673_));
 AO21x1_ASAP7_75t_R _29129_ (.A1(_06518_),
    .A2(net4617),
    .B(net6027),
    .Y(_06674_));
 NOR2x1_ASAP7_75t_R _29130_ (.A(net5594),
    .B(_06615_),
    .Y(_06675_));
 AOI21x1_ASAP7_75t_R _29132_ (.A1(_06674_),
    .A2(_06675_),
    .B(net5350),
    .Y(_06677_));
 AOI21x1_ASAP7_75t_R _29133_ (.A1(net5599),
    .A2(net5603),
    .B(net6031),
    .Y(_06678_));
 NAND2x1_ASAP7_75t_R _29134_ (.A(net4535),
    .B(_06678_),
    .Y(_06679_));
 AO21x1_ASAP7_75t_R _29135_ (.A1(net6035),
    .A2(net6036),
    .B(_06505_),
    .Y(_06680_));
 NAND2x1_ASAP7_75t_R _29136_ (.A(net5597),
    .B(net5082),
    .Y(_06681_));
 NAND2x1_ASAP7_75t_R _29137_ (.A(_06680_),
    .B(_06681_),
    .Y(_06682_));
 AOI21x1_ASAP7_75t_R _29138_ (.A1(net6026),
    .A2(_06682_),
    .B(net6016),
    .Y(_06683_));
 NAND2x1_ASAP7_75t_R _29139_ (.A(_06679_),
    .B(_06683_),
    .Y(_06684_));
 AOI21x1_ASAP7_75t_R _29140_ (.A1(_06677_),
    .A2(_06684_),
    .B(net6032),
    .Y(_06685_));
 NAND2x1_ASAP7_75t_R _29141_ (.A(_06673_),
    .B(_06685_),
    .Y(_06686_));
 NAND2x1_ASAP7_75t_R _29142_ (.A(_06661_),
    .B(_06686_),
    .Y(_06687_));
 OAI21x1_ASAP7_75t_R _29143_ (.A1(_06631_),
    .A2(_06579_),
    .B(_06687_),
    .Y(_00144_));
 NOR2x1_ASAP7_75t_R _29144_ (.A(_06517_),
    .B(net5600),
    .Y(_06688_));
 INVx1_ASAP7_75t_R _29145_ (.A(_06688_),
    .Y(_06689_));
 AOI21x1_ASAP7_75t_R _29146_ (.A1(net5600),
    .A2(net5083),
    .B(net6026),
    .Y(_06690_));
 AOI22x1_ASAP7_75t_R _29147_ (.A1(_06665_),
    .A2(net4488),
    .B1(_06689_),
    .B2(_06690_),
    .Y(_06691_));
 NOR2x1_ASAP7_75t_R _29148_ (.A(net5593),
    .B(_06691_),
    .Y(_06692_));
 NAND2x1_ASAP7_75t_R _29149_ (.A(net5599),
    .B(net5079),
    .Y(_06693_));
 INVx1_ASAP7_75t_R _29150_ (.A(_06693_),
    .Y(_06694_));
 NOR2x1_ASAP7_75t_R _29151_ (.A(_06694_),
    .B(_06656_),
    .Y(_06695_));
 NAND2x1_ASAP7_75t_R _29152_ (.A(net5598),
    .B(net6027),
    .Y(_06696_));
 OA21x2_ASAP7_75t_R _29153_ (.A1(_06696_),
    .A2(net5083),
    .B(net5593),
    .Y(_06697_));
 OAI21x1_ASAP7_75t_R _29154_ (.A1(net6018),
    .A2(net4824),
    .B(_06697_),
    .Y(_06698_));
 OAI21x1_ASAP7_75t_R _29155_ (.A1(_06695_),
    .A2(_06698_),
    .B(net5348),
    .Y(_06699_));
 NOR2x1_ASAP7_75t_R _29156_ (.A(net4720),
    .B(net5600),
    .Y(_06700_));
 AO21x1_ASAP7_75t_R _29157_ (.A1(net5346),
    .A2(net5083),
    .B(net6019),
    .Y(_06701_));
 AO21x1_ASAP7_75t_R _29158_ (.A1(net6033),
    .A2(net6034),
    .B(net4795),
    .Y(_06702_));
 OA21x2_ASAP7_75t_R _29159_ (.A1(_06702_),
    .A2(net6028),
    .B(net5594),
    .Y(_06703_));
 OAI21x1_ASAP7_75t_R _29160_ (.A1(_06700_),
    .A2(_06701_),
    .B(_06703_),
    .Y(_06704_));
 AOI21x1_ASAP7_75t_R _29161_ (.A1(net5603),
    .A2(net5083),
    .B(net5600),
    .Y(_06705_));
 NAND2x1_ASAP7_75t_R _29162_ (.A(net6018),
    .B(_06705_),
    .Y(_06706_));
 NAND2x1_ASAP7_75t_R _29163_ (.A(net5599),
    .B(net5590),
    .Y(_06707_));
 OA21x2_ASAP7_75t_R _29164_ (.A1(net5599),
    .A2(net4616),
    .B(net6025),
    .Y(_06708_));
 AOI21x1_ASAP7_75t_R _29165_ (.A1(net5341),
    .A2(_06708_),
    .B(net5594),
    .Y(_06709_));
 AOI21x1_ASAP7_75t_R _29166_ (.A1(_06706_),
    .A2(_06709_),
    .B(net5348),
    .Y(_06710_));
 NAND2x1_ASAP7_75t_R _29167_ (.A(_06704_),
    .B(_06710_),
    .Y(_06711_));
 OAI21x1_ASAP7_75t_R _29168_ (.A1(_06692_),
    .A2(_06699_),
    .B(_06711_),
    .Y(_06712_));
 NAND2x1_ASAP7_75t_R _29170_ (.A(_06583_),
    .B(_06567_),
    .Y(_06714_));
 INVx1_ASAP7_75t_R _29171_ (.A(_06714_),
    .Y(_06715_));
 NAND2x1_ASAP7_75t_R _29172_ (.A(net5590),
    .B(net5079),
    .Y(_06716_));
 AOI21x1_ASAP7_75t_R _29173_ (.A1(_06716_),
    .A2(_06678_),
    .B(net6017),
    .Y(_06717_));
 OAI21x1_ASAP7_75t_R _29174_ (.A1(net6018),
    .A2(_06715_),
    .B(_06717_),
    .Y(_06718_));
 AOI21x1_ASAP7_75t_R _29175_ (.A1(net4452),
    .A2(_06588_),
    .B(net5593),
    .Y(_06719_));
 NAND2x1_ASAP7_75t_R _29176_ (.A(net5600),
    .B(net5079),
    .Y(_06720_));
 AO21x1_ASAP7_75t_R _29177_ (.A1(_06720_),
    .A2(_06702_),
    .B(net6027),
    .Y(_06721_));
 AOI21x1_ASAP7_75t_R _29178_ (.A1(_06719_),
    .A2(_06721_),
    .B(net5350),
    .Y(_06722_));
 NAND2x1_ASAP7_75t_R _29179_ (.A(_06718_),
    .B(_06722_),
    .Y(_06723_));
 AOI21x1_ASAP7_75t_R _29180_ (.A1(_06599_),
    .A2(_06537_),
    .B(net6016),
    .Y(_06724_));
 OAI21x1_ASAP7_75t_R _29181_ (.A1(net6031),
    .A2(_06646_),
    .B(_06724_),
    .Y(_06725_));
 AOI21x1_ASAP7_75t_R _29182_ (.A1(net6028),
    .A2(net5351),
    .B(net5594),
    .Y(_06726_));
 OA21x2_ASAP7_75t_R _29183_ (.A1(net6028),
    .A2(_06670_),
    .B(net5340),
    .Y(_06727_));
 AOI21x1_ASAP7_75t_R _29184_ (.A1(_06726_),
    .A2(_06727_),
    .B(net5591),
    .Y(_06728_));
 AOI21x1_ASAP7_75t_R _29185_ (.A1(_06725_),
    .A2(_06728_),
    .B(net5588),
    .Y(_06729_));
 AOI21x1_ASAP7_75t_R _29186_ (.A1(_06723_),
    .A2(_06729_),
    .B(net6014),
    .Y(_06730_));
 OAI21x1_ASAP7_75t_R _29187_ (.A1(net6032),
    .A2(_06712_),
    .B(_06730_),
    .Y(_06731_));
 AO21x1_ASAP7_75t_R _29188_ (.A1(net5083),
    .A2(net5598),
    .B(net6031),
    .Y(_06732_));
 NOR2x1_ASAP7_75t_R _29189_ (.A(net5346),
    .B(_06732_),
    .Y(_06733_));
 AO21x1_ASAP7_75t_R _29190_ (.A1(_06615_),
    .A2(net5347),
    .B(net5591),
    .Y(_06734_));
 OAI21x1_ASAP7_75t_R _29192_ (.A1(_06733_),
    .A2(_06734_),
    .B(net6017),
    .Y(_06736_));
 NOR2x1_ASAP7_75t_R _29193_ (.A(_06705_),
    .B(_06714_),
    .Y(_06737_));
 AO21x1_ASAP7_75t_R _29194_ (.A1(net5600),
    .A2(_06517_),
    .B(net6029),
    .Y(_06738_));
 OA21x2_ASAP7_75t_R _29195_ (.A1(_06738_),
    .A2(_06694_),
    .B(net5591),
    .Y(_06739_));
 OA21x2_ASAP7_75t_R _29196_ (.A1(net6018),
    .A2(_06737_),
    .B(_06739_),
    .Y(_06740_));
 NAND2x1_ASAP7_75t_R _29197_ (.A(_01379_),
    .B(net6031),
    .Y(_06741_));
 OAI21x1_ASAP7_75t_R _29198_ (.A1(net5080),
    .A2(_06632_),
    .B(_06515_),
    .Y(_06742_));
 OAI21x1_ASAP7_75t_R _29199_ (.A1(net5591),
    .A2(_06741_),
    .B(net4437),
    .Y(_06743_));
 AOI21x1_ASAP7_75t_R _29200_ (.A1(net5593),
    .A2(_06743_),
    .B(net5588),
    .Y(_06744_));
 OAI21x1_ASAP7_75t_R _29201_ (.A1(_06736_),
    .A2(_06740_),
    .B(_06744_),
    .Y(_06745_));
 AOI21x1_ASAP7_75t_R _29202_ (.A1(net5347),
    .A2(_06615_),
    .B(net5350),
    .Y(_06746_));
 AO21x1_ASAP7_75t_R _29203_ (.A1(_06693_),
    .A2(_06518_),
    .B(net6031),
    .Y(_06747_));
 NAND2x1_ASAP7_75t_R _29204_ (.A(_06746_),
    .B(_06747_),
    .Y(_06748_));
 NOR2x1_ASAP7_75t_R _29205_ (.A(net6026),
    .B(net5083),
    .Y(_06749_));
 OAI21x1_ASAP7_75t_R _29206_ (.A1(_06749_),
    .A2(_06678_),
    .B(_06720_),
    .Y(_06750_));
 NOR2x1p5_ASAP7_75t_R _29207_ (.A(net5591),
    .B(_06665_),
    .Y(_06751_));
 AOI21x1_ASAP7_75t_R _29208_ (.A1(_06751_),
    .A2(_06750_),
    .B(net6017),
    .Y(_06752_));
 AOI21x1_ASAP7_75t_R _29209_ (.A1(_06748_),
    .A2(_06752_),
    .B(net6032),
    .Y(_06753_));
 AO21x1_ASAP7_75t_R _29210_ (.A1(net6033),
    .A2(net6034),
    .B(net4793),
    .Y(_06754_));
 NAND2x1_ASAP7_75t_R _29211_ (.A(_06754_),
    .B(_06648_),
    .Y(_06755_));
 AOI21x1_ASAP7_75t_R _29212_ (.A1(net6023),
    .A2(_06755_),
    .B(net5591),
    .Y(_06756_));
 OAI21x1_ASAP7_75t_R _29213_ (.A1(_06700_),
    .A2(_06701_),
    .B(_06756_),
    .Y(_06757_));
 NAND2x1_ASAP7_75t_R _29214_ (.A(_06504_),
    .B(_06537_),
    .Y(_06758_));
 INVx1_ASAP7_75t_R _29215_ (.A(net4827),
    .Y(_06759_));
 OAI21x1_ASAP7_75t_R _29216_ (.A1(net6027),
    .A2(net4617),
    .B(net5591),
    .Y(_06760_));
 AOI21x1_ASAP7_75t_R _29217_ (.A1(net6018),
    .A2(_06759_),
    .B(_06760_),
    .Y(_06761_));
 AOI21x1_ASAP7_75t_R _29218_ (.A1(_06758_),
    .A2(_06761_),
    .B(net5593),
    .Y(_06762_));
 NAND2x1_ASAP7_75t_R _29219_ (.A(_06757_),
    .B(_06762_),
    .Y(_06763_));
 INVx1_ASAP7_75t_R _29220_ (.A(_06630_),
    .Y(_06764_));
 AOI21x1_ASAP7_75t_R _29221_ (.A1(_06753_),
    .A2(_06763_),
    .B(_06764_),
    .Y(_06765_));
 NAND2x1_ASAP7_75t_R _29222_ (.A(_06765_),
    .B(_06745_),
    .Y(_06766_));
 NAND2x1_ASAP7_75t_R _29223_ (.A(_06731_),
    .B(_06766_),
    .Y(_00145_));
 INVx1_ASAP7_75t_R _29224_ (.A(_06668_),
    .Y(_06767_));
 AOI21x1_ASAP7_75t_R _29225_ (.A1(net4490),
    .A2(net5343),
    .B(net6022),
    .Y(_06768_));
 OAI21x1_ASAP7_75t_R _29226_ (.A1(_06767_),
    .A2(_06768_),
    .B(net5592),
    .Y(_06769_));
 AOI21x1_ASAP7_75t_R _29227_ (.A1(net4489),
    .A2(_06681_),
    .B(net6023),
    .Y(_06770_));
 INVx1_ASAP7_75t_R _29228_ (.A(_06606_),
    .Y(_06771_));
 OA21x2_ASAP7_75t_R _29229_ (.A1(_06771_),
    .A2(net4610),
    .B(net6022),
    .Y(_06772_));
 OAI21x1_ASAP7_75t_R _29230_ (.A1(_06770_),
    .A2(_06772_),
    .B(net6015),
    .Y(_06773_));
 NAND2x1_ASAP7_75t_R _29231_ (.A(_06769_),
    .B(_06773_),
    .Y(_06774_));
 INVx2_ASAP7_75t_R _29232_ (.A(net4454),
    .Y(_06775_));
 AO21x1_ASAP7_75t_R _29233_ (.A1(net4538),
    .A2(_06775_),
    .B(net6022),
    .Y(_06776_));
 AOI21x1_ASAP7_75t_R _29234_ (.A1(net4796),
    .A2(net5600),
    .B(net6025),
    .Y(_06777_));
 NAND2x1_ASAP7_75t_R _29235_ (.A(net4822),
    .B(_06777_),
    .Y(_06778_));
 AO21x1_ASAP7_75t_R _29236_ (.A1(_06776_),
    .A2(_06778_),
    .B(net6016),
    .Y(_06779_));
 AOI21x1_ASAP7_75t_R _29237_ (.A1(net4614),
    .A2(_06681_),
    .B(net6030),
    .Y(_06780_));
 NOR2x1_ASAP7_75t_R _29238_ (.A(net5595),
    .B(net5602),
    .Y(_06781_));
 OA21x2_ASAP7_75t_R _29239_ (.A1(net5339),
    .A2(net4610),
    .B(net6030),
    .Y(_06782_));
 OAI21x1_ASAP7_75t_R _29240_ (.A1(_06780_),
    .A2(_06782_),
    .B(net6015),
    .Y(_06783_));
 AOI21x1_ASAP7_75t_R _29241_ (.A1(_06779_),
    .A2(_06783_),
    .B(net5349),
    .Y(_06784_));
 AOI211x1_ASAP7_75t_R _29242_ (.A1(_06774_),
    .A2(net5349),
    .B(_06784_),
    .C(net6032),
    .Y(_06785_));
 OAI21x1_ASAP7_75t_R _29243_ (.A1(net5083),
    .A2(net5351),
    .B(net6022),
    .Y(_06786_));
 NAND2x1_ASAP7_75t_R _29244_ (.A(net5592),
    .B(_06786_),
    .Y(_06787_));
 AOI21x1_ASAP7_75t_R _29245_ (.A1(_06754_),
    .A2(_06560_),
    .B(net6023),
    .Y(_06788_));
 OAI21x1_ASAP7_75t_R _29246_ (.A1(_06787_),
    .A2(_06788_),
    .B(net5591),
    .Y(_06789_));
 AOI21x1_ASAP7_75t_R _29247_ (.A1(net5595),
    .A2(net5082),
    .B(net6023),
    .Y(_06790_));
 AND2x2_ASAP7_75t_R _29248_ (.A(_06790_),
    .B(_06648_),
    .Y(_06791_));
 NOR2x1_ASAP7_75t_R _29249_ (.A(_06781_),
    .B(_06532_),
    .Y(_06792_));
 OA21x2_ASAP7_75t_R _29250_ (.A1(_06791_),
    .A2(_06792_),
    .B(net6015),
    .Y(_06793_));
 OAI21x1_ASAP7_75t_R _29251_ (.A1(_06789_),
    .A2(_06793_),
    .B(net6032),
    .Y(_06794_));
 OAI21x1_ASAP7_75t_R _29252_ (.A1(net5597),
    .A2(net5079),
    .B(net5602),
    .Y(_06795_));
 NAND2x1_ASAP7_75t_R _29253_ (.A(net6025),
    .B(_06795_),
    .Y(_06796_));
 AO21x1_ASAP7_75t_R _29254_ (.A1(net4614),
    .A2(_06702_),
    .B(net6025),
    .Y(_06797_));
 AO21x1_ASAP7_75t_R _29255_ (.A1(_06796_),
    .A2(_06797_),
    .B(net5594),
    .Y(_06798_));
 NAND3x1_ASAP7_75t_R _29256_ (.A(_06790_),
    .B(net5341),
    .C(_06670_),
    .Y(_06799_));
 NAND3x1_ASAP7_75t_R _29257_ (.A(_06799_),
    .B(net5594),
    .C(_06679_),
    .Y(_06800_));
 AOI21x1_ASAP7_75t_R _29258_ (.A1(_06798_),
    .A2(_06800_),
    .B(net5591),
    .Y(_06801_));
 OAI21x1_ASAP7_75t_R _29259_ (.A1(_06794_),
    .A2(_06801_),
    .B(net6014),
    .Y(_06802_));
 AND2x2_ASAP7_75t_R _29260_ (.A(_01367_),
    .B(net4795),
    .Y(_06803_));
 AO21x1_ASAP7_75t_R _29261_ (.A1(net6033),
    .A2(net6034),
    .B(_06803_),
    .Y(_06804_));
 AOI21x1_ASAP7_75t_R _29262_ (.A1(net4486),
    .A2(_06560_),
    .B(net6022),
    .Y(_06805_));
 NAND2x1_ASAP7_75t_R _29263_ (.A(net6016),
    .B(_06742_),
    .Y(_06806_));
 AOI21x1_ASAP7_75t_R _29264_ (.A1(net6024),
    .A2(_06688_),
    .B(net6016),
    .Y(_06807_));
 AO21x1_ASAP7_75t_R _29265_ (.A1(net4538),
    .A2(_06670_),
    .B(net6022),
    .Y(_06808_));
 AOI21x1_ASAP7_75t_R _29266_ (.A1(_06807_),
    .A2(_06808_),
    .B(net5350),
    .Y(_06809_));
 OAI21x1_ASAP7_75t_R _29267_ (.A1(_06805_),
    .A2(_06806_),
    .B(_06809_),
    .Y(_06810_));
 NAND2x1_ASAP7_75t_R _29268_ (.A(_01381_),
    .B(net6030),
    .Y(_06811_));
 NAND2x1_ASAP7_75t_R _29269_ (.A(_06811_),
    .B(_06786_),
    .Y(_06812_));
 OA21x2_ASAP7_75t_R _29270_ (.A1(_01383_),
    .A2(net6030),
    .B(net6015),
    .Y(_06813_));
 AOI21x1_ASAP7_75t_R _29271_ (.A1(_06813_),
    .A2(_06796_),
    .B(net5591),
    .Y(_06814_));
 OAI21x1_ASAP7_75t_R _29272_ (.A1(net6015),
    .A2(_06812_),
    .B(_06814_),
    .Y(_06815_));
 AOI21x1_ASAP7_75t_R _29273_ (.A1(_06810_),
    .A2(_06815_),
    .B(net5589),
    .Y(_06816_));
 AO21x1_ASAP7_75t_R _29274_ (.A1(net5590),
    .A2(net5600),
    .B(net6021),
    .Y(_06817_));
 NOR2x1_ASAP7_75t_R _29275_ (.A(_06694_),
    .B(_06817_),
    .Y(_06818_));
 AO21x1_ASAP7_75t_R _29276_ (.A1(_06678_),
    .A2(net4536),
    .B(net5593),
    .Y(_06819_));
 OAI21x1_ASAP7_75t_R _29277_ (.A1(net5083),
    .A2(net5343),
    .B(_06537_),
    .Y(_06820_));
 OA21x2_ASAP7_75t_R _29278_ (.A1(_01382_),
    .A2(net6029),
    .B(net5592),
    .Y(_06821_));
 AOI21x1_ASAP7_75t_R _29279_ (.A1(_06820_),
    .A2(_06821_),
    .B(net5350),
    .Y(_06822_));
 OAI21x1_ASAP7_75t_R _29280_ (.A1(_06818_),
    .A2(_06819_),
    .B(_06822_),
    .Y(_06823_));
 NOR2x1_ASAP7_75t_R _29281_ (.A(net6020),
    .B(_06555_),
    .Y(_06824_));
 AOI22x1_ASAP7_75t_R _29282_ (.A1(_06824_),
    .A2(net4536),
    .B1(_06518_),
    .B2(net5342),
    .Y(_06825_));
 NAND2x1_ASAP7_75t_R _29283_ (.A(_01379_),
    .B(net6018),
    .Y(_06826_));
 AOI21x1_ASAP7_75t_R _29284_ (.A1(net5598),
    .A2(net5603),
    .B(net6018),
    .Y(_06827_));
 AOI21x1_ASAP7_75t_R _29285_ (.A1(_06716_),
    .A2(_06827_),
    .B(net6017),
    .Y(_06828_));
 AOI21x1_ASAP7_75t_R _29286_ (.A1(_06826_),
    .A2(_06828_),
    .B(net5591),
    .Y(_06829_));
 OAI21x1_ASAP7_75t_R _29287_ (.A1(net5593),
    .A2(_06825_),
    .B(_06829_),
    .Y(_06830_));
 AOI21x1_ASAP7_75t_R _29288_ (.A1(_06823_),
    .A2(_06830_),
    .B(net6032),
    .Y(_06831_));
 OAI21x1_ASAP7_75t_R _29289_ (.A1(_06816_),
    .A2(_06831_),
    .B(_06764_),
    .Y(_06832_));
 OAI21x1_ASAP7_75t_R _29290_ (.A1(_06785_),
    .A2(_06802_),
    .B(_06832_),
    .Y(_00146_));
 AND3x1_ASAP7_75t_R _29291_ (.A(net5347),
    .B(net6026),
    .C(net4451),
    .Y(_06833_));
 NAND2x1_ASAP7_75t_R _29292_ (.A(_06716_),
    .B(net4827),
    .Y(_06834_));
 AO21x1_ASAP7_75t_R _29293_ (.A1(_06834_),
    .A2(net6018),
    .B(net5591),
    .Y(_06835_));
 AO21x1_ASAP7_75t_R _29294_ (.A1(_06754_),
    .A2(_06670_),
    .B(net6023),
    .Y(_06836_));
 NOR2x1_ASAP7_75t_R _29295_ (.A(net5350),
    .B(_06792_),
    .Y(_06837_));
 AOI21x1_ASAP7_75t_R _29296_ (.A1(_06836_),
    .A2(_06837_),
    .B(net6015),
    .Y(_06838_));
 OA21x2_ASAP7_75t_R _29297_ (.A1(_06833_),
    .A2(_06835_),
    .B(_06838_),
    .Y(_06839_));
 AND2x2_ASAP7_75t_R _29298_ (.A(_06689_),
    .B(_06537_),
    .Y(_06840_));
 AO21x1_ASAP7_75t_R _29299_ (.A1(_06690_),
    .A2(_06556_),
    .B(net5350),
    .Y(_06841_));
 AOI21x1_ASAP7_75t_R _29300_ (.A1(net6028),
    .A2(net4453),
    .B(net5591),
    .Y(_06842_));
 OAI21x1_ASAP7_75t_R _29301_ (.A1(net5346),
    .A2(_06732_),
    .B(_06842_),
    .Y(_06843_));
 OAI21x1_ASAP7_75t_R _29302_ (.A1(_06840_),
    .A2(_06841_),
    .B(_06843_),
    .Y(_06844_));
 AO21x1_ASAP7_75t_R _29303_ (.A1(_06844_),
    .A2(net6016),
    .B(net5588),
    .Y(_06845_));
 NOR2x1_ASAP7_75t_R _29304_ (.A(_06839_),
    .B(_06845_),
    .Y(_06846_));
 NAND2x1_ASAP7_75t_R _29305_ (.A(net5593),
    .B(_06696_),
    .Y(_06847_));
 OA21x2_ASAP7_75t_R _29306_ (.A1(_06834_),
    .A2(_06847_),
    .B(net5348),
    .Y(_06848_));
 AO21x1_ASAP7_75t_R _29307_ (.A1(net6035),
    .A2(net6036),
    .B(net4796),
    .Y(_06849_));
 AO21x1_ASAP7_75t_R _29308_ (.A1(net4452),
    .A2(_06849_),
    .B(net6028),
    .Y(_06850_));
 NAND2x1_ASAP7_75t_R _29309_ (.A(_06850_),
    .B(_06709_),
    .Y(_06851_));
 AO21x1_ASAP7_75t_R _29310_ (.A1(_06848_),
    .A2(_06851_),
    .B(net6032),
    .Y(_06852_));
 AO21x1_ASAP7_75t_R _29311_ (.A1(net4451),
    .A2(net4487),
    .B(net6026),
    .Y(_06853_));
 AO21x1_ASAP7_75t_R _29312_ (.A1(net4827),
    .A2(net4826),
    .B(net6018),
    .Y(_06854_));
 AOI21x1_ASAP7_75t_R _29313_ (.A1(_06853_),
    .A2(_06854_),
    .B(net5594),
    .Y(_06855_));
 OAI21x1_ASAP7_75t_R _29314_ (.A1(_06705_),
    .A2(_06656_),
    .B(net5593),
    .Y(_06856_));
 AOI21x1_ASAP7_75t_R _29315_ (.A1(_06715_),
    .A2(net4436),
    .B(_06856_),
    .Y(_06857_));
 OA21x2_ASAP7_75t_R _29316_ (.A1(_06855_),
    .A2(_06857_),
    .B(net5591),
    .Y(_06858_));
 OAI21x1_ASAP7_75t_R _29317_ (.A1(_06852_),
    .A2(_06858_),
    .B(_06764_),
    .Y(_06859_));
 AO21x1_ASAP7_75t_R _29318_ (.A1(_06849_),
    .A2(_06804_),
    .B(net6022),
    .Y(_06860_));
 AOI21x1_ASAP7_75t_R _29319_ (.A1(_06742_),
    .A2(_06860_),
    .B(net6016),
    .Y(_06861_));
 OA21x2_ASAP7_75t_R _29320_ (.A1(_06732_),
    .A2(_06771_),
    .B(net6016),
    .Y(_06862_));
 OAI21x1_ASAP7_75t_R _29321_ (.A1(_06861_),
    .A2(_06862_),
    .B(net5350),
    .Y(_06863_));
 AOI21x1_ASAP7_75t_R _29322_ (.A1(_06650_),
    .A2(_06717_),
    .B(net5350),
    .Y(_06864_));
 AO21x1_ASAP7_75t_R _29323_ (.A1(net4538),
    .A2(_06606_),
    .B(net6030),
    .Y(_06865_));
 NOR2x1_ASAP7_75t_R _29324_ (.A(net5597),
    .B(_06522_),
    .Y(_06866_));
 NAND2x1_ASAP7_75t_R _29325_ (.A(net5080),
    .B(_06866_),
    .Y(_06867_));
 INVx1_ASAP7_75t_R _29326_ (.A(_06666_),
    .Y(_06868_));
 OAI21x1_ASAP7_75t_R _29327_ (.A1(net6024),
    .A2(_06868_),
    .B(net6016),
    .Y(_06869_));
 INVx1_ASAP7_75t_R _29328_ (.A(_06869_),
    .Y(_06870_));
 NAND3x1_ASAP7_75t_R _29329_ (.A(_06865_),
    .B(_06867_),
    .C(_06870_),
    .Y(_06871_));
 AOI21x1_ASAP7_75t_R _29330_ (.A1(_06864_),
    .A2(_06871_),
    .B(net6032),
    .Y(_06872_));
 NAND2x1_ASAP7_75t_R _29331_ (.A(_06863_),
    .B(_06872_),
    .Y(_06873_));
 OA21x2_ASAP7_75t_R _29332_ (.A1(net4485),
    .A2(net6022),
    .B(net5591),
    .Y(_06874_));
 AOI21x1_ASAP7_75t_R _29333_ (.A1(_06778_),
    .A2(_06874_),
    .B(net6016),
    .Y(_06875_));
 AO21x1_ASAP7_75t_R _29334_ (.A1(_06606_),
    .A2(_06804_),
    .B(net6022),
    .Y(_06876_));
 AOI21x1_ASAP7_75t_R _29335_ (.A1(net4452),
    .A2(_06618_),
    .B(net5591),
    .Y(_06877_));
 NAND2x1_ASAP7_75t_R _29336_ (.A(_06876_),
    .B(_06877_),
    .Y(_06878_));
 AOI21x1_ASAP7_75t_R _29337_ (.A1(_06875_),
    .A2(_06878_),
    .B(net5589),
    .Y(_06879_));
 NAND2x1_ASAP7_75t_R _29338_ (.A(net6030),
    .B(net4453),
    .Y(_06880_));
 NAND2x1_ASAP7_75t_R _29339_ (.A(net5344),
    .B(_06515_),
    .Y(_06881_));
 AOI21x1_ASAP7_75t_R _29340_ (.A1(_06880_),
    .A2(_06881_),
    .B(net5591),
    .Y(_06882_));
 NOR2x1_ASAP7_75t_R _29341_ (.A(net6030),
    .B(net4452),
    .Y(_06883_));
 AO22x1_ASAP7_75t_R _29342_ (.A1(net6030),
    .A2(_06640_),
    .B1(_06883_),
    .B2(net5591),
    .Y(_06884_));
 OAI21x1_ASAP7_75t_R _29343_ (.A1(_06882_),
    .A2(_06884_),
    .B(net6016),
    .Y(_06885_));
 AOI21x1_ASAP7_75t_R _29344_ (.A1(_06879_),
    .A2(_06885_),
    .B(_06764_),
    .Y(_06886_));
 NAND2x1_ASAP7_75t_R _29345_ (.A(_06873_),
    .B(_06886_),
    .Y(_06887_));
 OAI21x1_ASAP7_75t_R _29346_ (.A1(_06846_),
    .A2(_06859_),
    .B(_06887_),
    .Y(_00147_));
 INVx1_ASAP7_75t_R _29347_ (.A(_01373_),
    .Y(_06888_));
 NAND2x1_ASAP7_75t_R _29348_ (.A(_06888_),
    .B(net6020),
    .Y(_06889_));
 OAI21x1_ASAP7_75t_R _29349_ (.A1(net6020),
    .A2(net4536),
    .B(_06889_),
    .Y(_06890_));
 AO21x1_ASAP7_75t_R _29350_ (.A1(_06890_),
    .A2(net5593),
    .B(net5350),
    .Y(_06891_));
 NAND2x1_ASAP7_75t_R _29351_ (.A(net5340),
    .B(_06634_),
    .Y(_06892_));
 INVx1_ASAP7_75t_R _29352_ (.A(_06892_),
    .Y(_06893_));
 AO21x1_ASAP7_75t_R _29353_ (.A1(net5079),
    .A2(net5603),
    .B(net5600),
    .Y(_06894_));
 OAI21x1_ASAP7_75t_R _29354_ (.A1(net6026),
    .A2(_06894_),
    .B(net6017),
    .Y(_06895_));
 NOR2x1_ASAP7_75t_R _29355_ (.A(_06893_),
    .B(_06895_),
    .Y(_06896_));
 OAI21x1_ASAP7_75t_R _29356_ (.A1(_06891_),
    .A2(_06896_),
    .B(net6032),
    .Y(_06897_));
 AOI21x1_ASAP7_75t_R _29357_ (.A1(net5340),
    .A2(_06587_),
    .B(net6027),
    .Y(_06898_));
 NOR2x1_ASAP7_75t_R _29358_ (.A(_06573_),
    .B(_06635_),
    .Y(_06899_));
 OAI21x1_ASAP7_75t_R _29359_ (.A1(_06898_),
    .A2(_06899_),
    .B(net6017),
    .Y(_06900_));
 AO21x1_ASAP7_75t_R _29360_ (.A1(_06575_),
    .A2(_06674_),
    .B(net6017),
    .Y(_06901_));
 AOI21x1_ASAP7_75t_R _29361_ (.A1(_06900_),
    .A2(_06901_),
    .B(net5591),
    .Y(_06902_));
 OAI21x1_ASAP7_75t_R _29362_ (.A1(_06897_),
    .A2(_06902_),
    .B(net6014),
    .Y(_06903_));
 AO21x1_ASAP7_75t_R _29363_ (.A1(net5600),
    .A2(net4797),
    .B(net6029),
    .Y(_06904_));
 NAND2x1_ASAP7_75t_R _29364_ (.A(net6017),
    .B(_06904_),
    .Y(_06905_));
 OA21x2_ASAP7_75t_R _29365_ (.A1(net5351),
    .A2(net5079),
    .B(net6029),
    .Y(_06906_));
 OAI21x1_ASAP7_75t_R _29366_ (.A1(_06905_),
    .A2(_06906_),
    .B(net5591),
    .Y(_06907_));
 OA21x2_ASAP7_75t_R _29367_ (.A1(net5600),
    .A2(net4613),
    .B(net6021),
    .Y(_06908_));
 AOI21x1_ASAP7_75t_R _29368_ (.A1(net4536),
    .A2(_06908_),
    .B(net6017),
    .Y(_06909_));
 AND2x2_ASAP7_75t_R _29369_ (.A(_06909_),
    .B(_06589_),
    .Y(_06910_));
 OAI21x1_ASAP7_75t_R _29370_ (.A1(_06907_),
    .A2(_06910_),
    .B(net5588),
    .Y(_06911_));
 AND3x1_ASAP7_75t_R _29371_ (.A(net5351),
    .B(net6021),
    .C(_06504_),
    .Y(_06912_));
 AO21x1_ASAP7_75t_R _29372_ (.A1(_06615_),
    .A2(net5347),
    .B(net5593),
    .Y(_06913_));
 NOR2x1_ASAP7_75t_R _29373_ (.A(_06912_),
    .B(_06913_),
    .Y(_06914_));
 AO21x1_ASAP7_75t_R _29374_ (.A1(net4822),
    .A2(net4615),
    .B(net6029),
    .Y(_06915_));
 NOR2x1_ASAP7_75t_R _29375_ (.A(net6017),
    .B(net5338),
    .Y(_06916_));
 AO21x1_ASAP7_75t_R _29376_ (.A1(_06915_),
    .A2(_06916_),
    .B(net5591),
    .Y(_06917_));
 NOR2x1_ASAP7_75t_R _29377_ (.A(_06914_),
    .B(_06917_),
    .Y(_06918_));
 NOR2x1_ASAP7_75t_R _29378_ (.A(_06911_),
    .B(_06918_),
    .Y(_06919_));
 INVx1_ASAP7_75t_R _29379_ (.A(_06828_),
    .Y(_06920_));
 OAI21x1_ASAP7_75t_R _29380_ (.A1(_06920_),
    .A2(_06733_),
    .B(net5350),
    .Y(_06921_));
 AND2x2_ASAP7_75t_R _29381_ (.A(_06827_),
    .B(_06518_),
    .Y(_06922_));
 OA21x2_ASAP7_75t_R _29382_ (.A1(_06922_),
    .A2(_06898_),
    .B(net6017),
    .Y(_06923_));
 AO21x1_ASAP7_75t_R _29383_ (.A1(net5603),
    .A2(net5600),
    .B(net6018),
    .Y(_06924_));
 AOI21x1_ASAP7_75t_R _29384_ (.A1(_06738_),
    .A2(_06924_),
    .B(_06694_),
    .Y(_06925_));
 NOR2x1_ASAP7_75t_R _29385_ (.A(_06640_),
    .B(_06634_),
    .Y(_06926_));
 AOI21x1_ASAP7_75t_R _29386_ (.A1(net6017),
    .A2(_06926_),
    .B(net5350),
    .Y(_06927_));
 OAI21x1_ASAP7_75t_R _29387_ (.A1(net6017),
    .A2(_06925_),
    .B(_06927_),
    .Y(_06928_));
 OAI21x1_ASAP7_75t_R _29388_ (.A1(_06921_),
    .A2(_06923_),
    .B(_06928_),
    .Y(_06929_));
 NOR2x1_ASAP7_75t_R _29389_ (.A(net6032),
    .B(_06929_),
    .Y(_06930_));
 AOI21x1_ASAP7_75t_R _29390_ (.A1(net4484),
    .A2(net4536),
    .B(net6021),
    .Y(_06931_));
 OAI21x1_ASAP7_75t_R _29391_ (.A1(_06931_),
    .A2(_06669_),
    .B(net5591),
    .Y(_06932_));
 NAND2x1_ASAP7_75t_R _29392_ (.A(net6019),
    .B(_06599_),
    .Y(_06933_));
 OAI21x1_ASAP7_75t_R _29393_ (.A1(_06933_),
    .A2(net4453),
    .B(net5592),
    .Y(_06934_));
 NOR2x1_ASAP7_75t_R _29394_ (.A(_06635_),
    .B(_06633_),
    .Y(_06935_));
 NOR2x1_ASAP7_75t_R _29395_ (.A(_06934_),
    .B(_06935_),
    .Y(_06936_));
 OAI21x1_ASAP7_75t_R _29396_ (.A1(_06932_),
    .A2(_06936_),
    .B(net6032),
    .Y(_06937_));
 AO21x1_ASAP7_75t_R _29397_ (.A1(net6035),
    .A2(net6036),
    .B(net4616),
    .Y(_06938_));
 INVx1_ASAP7_75t_R _29398_ (.A(_06938_),
    .Y(_06939_));
 AO21x1_ASAP7_75t_R _29399_ (.A1(net5596),
    .A2(net4794),
    .B(net6029),
    .Y(_06940_));
 OAI21x1_ASAP7_75t_R _29400_ (.A1(_06939_),
    .A2(_06940_),
    .B(net6016),
    .Y(_06941_));
 NOR2x1_ASAP7_75t_R _29401_ (.A(_06817_),
    .B(_06633_),
    .Y(_06942_));
 OAI21x1_ASAP7_75t_R _29402_ (.A1(_06941_),
    .A2(_06942_),
    .B(net5350),
    .Y(_06943_));
 INVx1_ASAP7_75t_R _29403_ (.A(_06504_),
    .Y(_06944_));
 OAI21x1_ASAP7_75t_R _29404_ (.A1(net4483),
    .A2(_06817_),
    .B(net5593),
    .Y(_06945_));
 NOR2x1_ASAP7_75t_R _29405_ (.A(_06945_),
    .B(_06647_),
    .Y(_06946_));
 NOR2x1_ASAP7_75t_R _29406_ (.A(_06943_),
    .B(_06946_),
    .Y(_06947_));
 OAI21x1_ASAP7_75t_R _29407_ (.A1(_06937_),
    .A2(_06947_),
    .B(_06764_),
    .Y(_06948_));
 OAI22x1_ASAP7_75t_R _29408_ (.A1(_06903_),
    .A2(_06919_),
    .B1(_06930_),
    .B2(_06948_),
    .Y(_00148_));
 AOI21x1_ASAP7_75t_R _29409_ (.A1(_06518_),
    .A2(net4452),
    .B(net6023),
    .Y(_06949_));
 AOI211x1_ASAP7_75t_R _29410_ (.A1(net6023),
    .A2(_06771_),
    .B(_06949_),
    .C(net6016),
    .Y(_06950_));
 AO21x1_ASAP7_75t_R _29411_ (.A1(net5340),
    .A2(net4611),
    .B(net6028),
    .Y(_06951_));
 OA21x2_ASAP7_75t_R _29412_ (.A1(net4535),
    .A2(net6019),
    .B(net6016),
    .Y(_06952_));
 AND2x2_ASAP7_75t_R _29413_ (.A(_06951_),
    .B(_06952_),
    .Y(_06953_));
 OAI21x1_ASAP7_75t_R _29414_ (.A1(_06950_),
    .A2(_06953_),
    .B(net5349),
    .Y(_06954_));
 INVx1_ASAP7_75t_R _29415_ (.A(_06705_),
    .Y(_06955_));
 AND3x1_ASAP7_75t_R _29416_ (.A(_06955_),
    .B(net6026),
    .C(net4487),
    .Y(_06956_));
 AO21x1_ASAP7_75t_R _29417_ (.A1(net4823),
    .A2(net4824),
    .B(net5594),
    .Y(_06957_));
 AO21x1_ASAP7_75t_R _29418_ (.A1(net5590),
    .A2(net6026),
    .B(net6017),
    .Y(_06958_));
 OA21x2_ASAP7_75t_R _29419_ (.A1(_06898_),
    .A2(_06958_),
    .B(net5591),
    .Y(_06959_));
 OAI21x1_ASAP7_75t_R _29420_ (.A1(_06956_),
    .A2(_06957_),
    .B(_06959_),
    .Y(_06960_));
 AOI21x1_ASAP7_75t_R _29421_ (.A1(_06954_),
    .A2(_06960_),
    .B(_06622_),
    .Y(_06961_));
 AOI211x1_ASAP7_75t_R _29422_ (.A1(net4826),
    .A2(net5338),
    .B(_06908_),
    .C(net5593),
    .Y(_06962_));
 AO21x1_ASAP7_75t_R _29423_ (.A1(net4451),
    .A2(net6018),
    .B(net6017),
    .Y(_06963_));
 AOI21x1_ASAP7_75t_R _29424_ (.A1(net4484),
    .A2(_06720_),
    .B(net6020),
    .Y(_06964_));
 OAI21x1_ASAP7_75t_R _29425_ (.A1(_06963_),
    .A2(_06964_),
    .B(net5350),
    .Y(_06965_));
 OAI21x1_ASAP7_75t_R _29426_ (.A1(_06962_),
    .A2(_06965_),
    .B(net5588),
    .Y(_06966_));
 NAND2x1_ASAP7_75t_R _29427_ (.A(net4617),
    .B(net5347),
    .Y(_06967_));
 AOI21x1_ASAP7_75t_R _29428_ (.A1(net4615),
    .A2(net4609),
    .B(net6019),
    .Y(_06968_));
 AOI211x1_ASAP7_75t_R _29429_ (.A1(_06967_),
    .A2(net6019),
    .B(_06968_),
    .C(net6016),
    .Y(_06969_));
 OA21x2_ASAP7_75t_R _29430_ (.A1(net5083),
    .A2(net5344),
    .B(_06777_),
    .Y(_06970_));
 NAND2x1_ASAP7_75t_R _29431_ (.A(net4613),
    .B(net6029),
    .Y(_06971_));
 NAND2x1_ASAP7_75t_R _29432_ (.A(_06971_),
    .B(_06641_),
    .Y(_06972_));
 OAI21x1_ASAP7_75t_R _29433_ (.A1(_06970_),
    .A2(_06972_),
    .B(net5591),
    .Y(_06973_));
 NOR2x1_ASAP7_75t_R _29434_ (.A(_06969_),
    .B(_06973_),
    .Y(_06974_));
 OAI21x1_ASAP7_75t_R _29435_ (.A1(_06966_),
    .A2(_06974_),
    .B(_06764_),
    .Y(_06975_));
 AO21x1_ASAP7_75t_R _29436_ (.A1(_06681_),
    .A2(_06670_),
    .B(net6027),
    .Y(_06976_));
 AND2x2_ASAP7_75t_R _29437_ (.A(_06976_),
    .B(_06589_),
    .Y(_06977_));
 INVx1_ASAP7_75t_R _29438_ (.A(_06680_),
    .Y(_06978_));
 AO21x1_ASAP7_75t_R _29439_ (.A1(_06978_),
    .A2(net6026),
    .B(net5594),
    .Y(_06979_));
 OA21x2_ASAP7_75t_R _29440_ (.A1(_06678_),
    .A2(_06749_),
    .B(_06938_),
    .Y(_06980_));
 OAI21x1_ASAP7_75t_R _29441_ (.A1(_06979_),
    .A2(_06980_),
    .B(net5350),
    .Y(_06981_));
 AOI21x1_ASAP7_75t_R _29442_ (.A1(net5594),
    .A2(_06977_),
    .B(_06981_),
    .Y(_06982_));
 AO21x1_ASAP7_75t_R _29443_ (.A1(net5083),
    .A2(net6025),
    .B(net6015),
    .Y(_06983_));
 NOR2x1_ASAP7_75t_R _29444_ (.A(_06572_),
    .B(_06732_),
    .Y(_06984_));
 OAI21x1_ASAP7_75t_R _29445_ (.A1(_06983_),
    .A2(_06984_),
    .B(net5591),
    .Y(_06985_));
 AND2x2_ASAP7_75t_R _29446_ (.A(_06777_),
    .B(net5341),
    .Y(_06986_));
 AOI211x1_ASAP7_75t_R _29447_ (.A1(net4424),
    .A2(_06596_),
    .B(_06986_),
    .C(net5594),
    .Y(_06987_));
 OAI21x1_ASAP7_75t_R _29448_ (.A1(_06985_),
    .A2(_06987_),
    .B(_06622_),
    .Y(_06988_));
 NOR2x1_ASAP7_75t_R _29449_ (.A(_06982_),
    .B(_06988_),
    .Y(_06989_));
 AO21x1_ASAP7_75t_R _29450_ (.A1(net6023),
    .A2(net4612),
    .B(net5594),
    .Y(_06990_));
 OAI21x1_ASAP7_75t_R _29451_ (.A1(_06708_),
    .A2(_06990_),
    .B(net5591),
    .Y(_06991_));
 OA21x2_ASAP7_75t_R _29452_ (.A1(net5345),
    .A2(net5079),
    .B(net6023),
    .Y(_06992_));
 AO21x1_ASAP7_75t_R _29453_ (.A1(net5599),
    .A2(net4608),
    .B(net6023),
    .Y(_06993_));
 NAND2x1_ASAP7_75t_R _29454_ (.A(net5594),
    .B(_06993_),
    .Y(_06994_));
 AOI21x1_ASAP7_75t_R _29455_ (.A1(_06596_),
    .A2(_06992_),
    .B(_06994_),
    .Y(_06995_));
 OAI21x1_ASAP7_75t_R _29456_ (.A1(_06991_),
    .A2(_06995_),
    .B(net6032),
    .Y(_06996_));
 AO21x1_ASAP7_75t_R _29457_ (.A1(net4539),
    .A2(_06680_),
    .B(net6023),
    .Y(_06997_));
 OA21x2_ASAP7_75t_R _29458_ (.A1(_06532_),
    .A2(_06939_),
    .B(_06997_),
    .Y(_06998_));
 AO21x1_ASAP7_75t_R _29459_ (.A1(_01369_),
    .A2(net6025),
    .B(net6015),
    .Y(_06999_));
 OAI21x1_ASAP7_75t_R _29460_ (.A1(_06999_),
    .A2(_06992_),
    .B(net5350),
    .Y(_07000_));
 AOI21x1_ASAP7_75t_R _29461_ (.A1(net6015),
    .A2(_06998_),
    .B(_07000_),
    .Y(_07001_));
 OAI21x1_ASAP7_75t_R _29462_ (.A1(_06996_),
    .A2(_07001_),
    .B(net6014),
    .Y(_07002_));
 OAI22x1_ASAP7_75t_R _29463_ (.A1(_06961_),
    .A2(_06975_),
    .B1(_06989_),
    .B2(_07002_),
    .Y(_00149_));
 INVx1_ASAP7_75t_R _29464_ (.A(net4492),
    .Y(_07003_));
 AOI21x1_ASAP7_75t_R _29465_ (.A1(_07003_),
    .A2(_06892_),
    .B(net5594),
    .Y(_07004_));
 AOI211x1_ASAP7_75t_R _29466_ (.A1(_06799_),
    .A2(net5594),
    .B(_07004_),
    .C(net5589),
    .Y(_07005_));
 OAI21x1_ASAP7_75t_R _29467_ (.A1(net6022),
    .A2(net4610),
    .B(net4537),
    .Y(_07006_));
 AOI21x1_ASAP7_75t_R _29468_ (.A1(net5080),
    .A2(_06866_),
    .B(net6016),
    .Y(_07007_));
 AOI22x1_ASAP7_75t_R _29469_ (.A1(_06612_),
    .A2(_06726_),
    .B1(_07006_),
    .B2(_07007_),
    .Y(_07008_));
 OAI21x1_ASAP7_75t_R _29470_ (.A1(net6032),
    .A2(_07008_),
    .B(net5349),
    .Y(_07009_));
 NOR2x1_ASAP7_75t_R _29471_ (.A(_07005_),
    .B(_07009_),
    .Y(_07010_));
 NAND2x1_ASAP7_75t_R _29472_ (.A(net5594),
    .B(_06795_),
    .Y(_07011_));
 AOI21x1_ASAP7_75t_R _29473_ (.A1(_06681_),
    .A2(net4825),
    .B(net6023),
    .Y(_07012_));
 OAI21x1_ASAP7_75t_R _29474_ (.A1(_07011_),
    .A2(_07012_),
    .B(net5589),
    .Y(_07013_));
 NAND2x1_ASAP7_75t_R _29475_ (.A(net4491),
    .B(_06690_),
    .Y(_07014_));
 NOR2x1_ASAP7_75t_R _29476_ (.A(net5590),
    .B(net5083),
    .Y(_07015_));
 OAI21x1_ASAP7_75t_R _29477_ (.A1(_06573_),
    .A2(_07015_),
    .B(net6025),
    .Y(_07016_));
 AOI21x1_ASAP7_75t_R _29478_ (.A1(_07014_),
    .A2(_07016_),
    .B(net5594),
    .Y(_07017_));
 OAI21x1_ASAP7_75t_R _29479_ (.A1(_07013_),
    .A2(_07017_),
    .B(net5591),
    .Y(_07018_));
 NAND2x1_ASAP7_75t_R _29480_ (.A(_01377_),
    .B(net6030),
    .Y(_07019_));
 INVx1_ASAP7_75t_R _29481_ (.A(_06986_),
    .Y(_07020_));
 AOI21x1_ASAP7_75t_R _29482_ (.A1(_07019_),
    .A2(_07020_),
    .B(net6015),
    .Y(_07021_));
 NOR2x1_ASAP7_75t_R _29483_ (.A(net5594),
    .B(_06690_),
    .Y(_07022_));
 AO21x1_ASAP7_75t_R _29484_ (.A1(net4539),
    .A2(_06938_),
    .B(net6019),
    .Y(_07023_));
 AO21x1_ASAP7_75t_R _29485_ (.A1(_07022_),
    .A2(_07023_),
    .B(_06622_),
    .Y(_07024_));
 NOR2x1_ASAP7_75t_R _29486_ (.A(_07021_),
    .B(_07024_),
    .Y(_07025_));
 OAI21x1_ASAP7_75t_R _29487_ (.A1(_07018_),
    .A2(_07025_),
    .B(net6014),
    .Y(_07026_));
 NOR2x1_ASAP7_75t_R _29488_ (.A(_07010_),
    .B(_07026_),
    .Y(_07027_));
 OAI21x1_ASAP7_75t_R _29489_ (.A1(_06640_),
    .A2(net5339),
    .B(net6030),
    .Y(_07028_));
 NAND2x1_ASAP7_75t_R _29490_ (.A(_06599_),
    .B(_06777_),
    .Y(_07029_));
 NAND3x1_ASAP7_75t_R _29491_ (.A(_07028_),
    .B(_07007_),
    .C(_07029_),
    .Y(_07030_));
 AOI21x1_ASAP7_75t_R _29492_ (.A1(_06670_),
    .A2(_06648_),
    .B(net6024),
    .Y(_07031_));
 NOR2x1_ASAP7_75t_R _29493_ (.A(_06869_),
    .B(_07031_),
    .Y(_07032_));
 AO21x1_ASAP7_75t_R _29494_ (.A1(net4822),
    .A2(_06775_),
    .B(net6030),
    .Y(_07033_));
 AOI21x1_ASAP7_75t_R _29495_ (.A1(_07032_),
    .A2(_07033_),
    .B(net5591),
    .Y(_07034_));
 NAND2x1_ASAP7_75t_R _29496_ (.A(_07030_),
    .B(_07034_),
    .Y(_07035_));
 OA21x2_ASAP7_75t_R _29497_ (.A1(net5602),
    .A2(net5596),
    .B(net6029),
    .Y(_07036_));
 NAND2x1_ASAP7_75t_R _29498_ (.A(net4826),
    .B(_07036_),
    .Y(_07037_));
 AO21x1_ASAP7_75t_R _29499_ (.A1(_01376_),
    .A2(_01380_),
    .B(net6029),
    .Y(_07038_));
 AND2x2_ASAP7_75t_R _29500_ (.A(_07038_),
    .B(net5592),
    .Y(_07039_));
 NAND2x1_ASAP7_75t_R _29501_ (.A(_07037_),
    .B(_07039_),
    .Y(_07040_));
 INVx1_ASAP7_75t_R _29502_ (.A(net4797),
    .Y(_07041_));
 AOI22x1_ASAP7_75t_R _29503_ (.A1(_06866_),
    .A2(net4607),
    .B1(_06688_),
    .B2(net6024),
    .Y(_07042_));
 AOI21x1_ASAP7_75t_R _29504_ (.A1(_06870_),
    .A2(_07042_),
    .B(net5350),
    .Y(_07043_));
 AOI21x1_ASAP7_75t_R _29505_ (.A1(_07040_),
    .A2(_07043_),
    .B(net6032),
    .Y(_07044_));
 NAND2x1_ASAP7_75t_R _29506_ (.A(_07035_),
    .B(_07044_),
    .Y(_07045_));
 AOI21x1_ASAP7_75t_R _29507_ (.A1(_06811_),
    .A2(_06786_),
    .B(net4427),
    .Y(_07046_));
 AOI21x1_ASAP7_75t_R _29508_ (.A1(net5595),
    .A2(net5590),
    .B(net6022),
    .Y(_07047_));
 OAI21x1_ASAP7_75t_R _29509_ (.A1(net5595),
    .A2(net4826),
    .B(_07047_),
    .Y(_07048_));
 NOR2x1_ASAP7_75t_R _29510_ (.A(_07041_),
    .B(net5597),
    .Y(_07049_));
 OA21x2_ASAP7_75t_R _29511_ (.A1(_06532_),
    .A2(_07049_),
    .B(net5592),
    .Y(_07050_));
 AOI21x1_ASAP7_75t_R _29512_ (.A1(_07048_),
    .A2(_07050_),
    .B(net5350),
    .Y(_07051_));
 OAI21x1_ASAP7_75t_R _29513_ (.A1(net5592),
    .A2(_07046_),
    .B(_07051_),
    .Y(_07052_));
 OA21x2_ASAP7_75t_R _29514_ (.A1(_06680_),
    .A2(net6025),
    .B(net6015),
    .Y(_07053_));
 OAI21x1_ASAP7_75t_R _29515_ (.A1(net5590),
    .A2(_06573_),
    .B(net6025),
    .Y(_07054_));
 AOI21x1_ASAP7_75t_R _29516_ (.A1(_07053_),
    .A2(_07054_),
    .B(net5591),
    .Y(_07055_));
 AO21x1_ASAP7_75t_R _29517_ (.A1(_06804_),
    .A2(_06775_),
    .B(net6030),
    .Y(_07056_));
 NAND3x1_ASAP7_75t_R _29518_ (.A(_06575_),
    .B(_07056_),
    .C(_07007_),
    .Y(_07057_));
 AOI21x1_ASAP7_75t_R _29519_ (.A1(_07055_),
    .A2(_07057_),
    .B(net5589),
    .Y(_07058_));
 NAND2x1_ASAP7_75t_R _29520_ (.A(_07052_),
    .B(_07058_),
    .Y(_07059_));
 AOI21x1_ASAP7_75t_R _29521_ (.A1(_07045_),
    .A2(_07059_),
    .B(net6014),
    .Y(_07060_));
 NOR2x1_ASAP7_75t_R _29522_ (.A(_07027_),
    .B(_07060_),
    .Y(_00150_));
 AOI21x1_ASAP7_75t_R _29523_ (.A1(net6026),
    .A2(_06955_),
    .B(_06963_),
    .Y(_07061_));
 AO21x1_ASAP7_75t_R _29524_ (.A1(net5346),
    .A2(net5083),
    .B(_06532_),
    .Y(_07062_));
 AO21x1_ASAP7_75t_R _29525_ (.A1(_07015_),
    .A2(net5599),
    .B(net6019),
    .Y(_07063_));
 AOI21x1_ASAP7_75t_R _29526_ (.A1(_07062_),
    .A2(_07063_),
    .B(net5594),
    .Y(_07064_));
 OAI21x1_ASAP7_75t_R _29527_ (.A1(_07061_),
    .A2(_07064_),
    .B(net5348),
    .Y(_07065_));
 NOR2x1_ASAP7_75t_R _29528_ (.A(_06694_),
    .B(_06924_),
    .Y(_07066_));
 OAI21x1_ASAP7_75t_R _29529_ (.A1(_06749_),
    .A2(_07066_),
    .B(net6017),
    .Y(_07067_));
 OAI21x1_ASAP7_75t_R _29530_ (.A1(net5598),
    .A2(_06587_),
    .B(_06594_),
    .Y(_07068_));
 AOI21x1_ASAP7_75t_R _29531_ (.A1(_06828_),
    .A2(_07068_),
    .B(net5348),
    .Y(_07069_));
 AOI21x1_ASAP7_75t_R _29532_ (.A1(_07067_),
    .A2(_07069_),
    .B(net5588),
    .Y(_07070_));
 NAND2x1_ASAP7_75t_R _29533_ (.A(_07065_),
    .B(_07070_),
    .Y(_07071_));
 AO21x1_ASAP7_75t_R _29534_ (.A1(net5590),
    .A2(net5598),
    .B(net5083),
    .Y(_07072_));
 AO21x1_ASAP7_75t_R _29535_ (.A1(_07072_),
    .A2(net6020),
    .B(net5350),
    .Y(_07073_));
 AO21x1_ASAP7_75t_R _29536_ (.A1(net5346),
    .A2(net5083),
    .B(_06944_),
    .Y(_07074_));
 NOR2x1_ASAP7_75t_R _29537_ (.A(net6020),
    .B(_07074_),
    .Y(_07075_));
 NAND2x1p5_ASAP7_75t_R _29538_ (.A(_06537_),
    .B(net4491),
    .Y(_07076_));
 AOI21x1_ASAP7_75t_R _29539_ (.A1(_07076_),
    .A2(net4428),
    .B(net5594),
    .Y(_07077_));
 OAI21x1_ASAP7_75t_R _29540_ (.A1(_07073_),
    .A2(_07075_),
    .B(_07077_),
    .Y(_07078_));
 AOI21x1_ASAP7_75t_R _29541_ (.A1(net6019),
    .A2(net4491),
    .B(net5350),
    .Y(_07079_));
 AOI21x1_ASAP7_75t_R _29542_ (.A1(_06892_),
    .A2(_07079_),
    .B(net6016),
    .Y(_07080_));
 AOI21x1_ASAP7_75t_R _29543_ (.A1(net4822),
    .A2(_07036_),
    .B(net5591),
    .Y(_07081_));
 NAND2x1_ASAP7_75t_R _29544_ (.A(_07029_),
    .B(_07081_),
    .Y(_07082_));
 AOI21x1_ASAP7_75t_R _29545_ (.A1(_07080_),
    .A2(_07082_),
    .B(net6032),
    .Y(_07083_));
 AOI21x1_ASAP7_75t_R _29546_ (.A1(_07078_),
    .A2(_07083_),
    .B(_06764_),
    .Y(_07084_));
 NAND2x1_ASAP7_75t_R _29547_ (.A(_07071_),
    .B(_07084_),
    .Y(_07085_));
 AOI211x1_ASAP7_75t_R _29548_ (.A1(_06924_),
    .A2(_06904_),
    .B(net4483),
    .C(net6017),
    .Y(_07086_));
 NAND2x1_ASAP7_75t_R _29549_ (.A(net4613),
    .B(net6019),
    .Y(_07087_));
 AOI21x1_ASAP7_75t_R _29550_ (.A1(_07087_),
    .A2(_07037_),
    .B(net5592),
    .Y(_07088_));
 OAI21x1_ASAP7_75t_R _29551_ (.A1(_07086_),
    .A2(_07088_),
    .B(net5350),
    .Y(_07089_));
 NAND2x1_ASAP7_75t_R _29552_ (.A(_06587_),
    .B(_06678_),
    .Y(_07090_));
 AOI21x1_ASAP7_75t_R _29553_ (.A1(_07090_),
    .A2(_06860_),
    .B(net5593),
    .Y(_07091_));
 OAI21x1_ASAP7_75t_R _29554_ (.A1(_06978_),
    .A2(_06664_),
    .B(net5594),
    .Y(_07092_));
 AOI21x1_ASAP7_75t_R _29555_ (.A1(net6020),
    .A2(_07074_),
    .B(_07092_),
    .Y(_07093_));
 OAI21x1_ASAP7_75t_R _29556_ (.A1(_07091_),
    .A2(_07093_),
    .B(net5591),
    .Y(_07094_));
 NAND2x1_ASAP7_75t_R _29557_ (.A(_07089_),
    .B(_07094_),
    .Y(_07095_));
 AND3x1_ASAP7_75t_R _29558_ (.A(net4826),
    .B(net6021),
    .C(net5351),
    .Y(_07096_));
 NAND2x1_ASAP7_75t_R _29559_ (.A(_01373_),
    .B(net6031),
    .Y(_07097_));
 AOI21x1_ASAP7_75t_R _29560_ (.A1(_07097_),
    .A2(_06649_),
    .B(net5350),
    .Y(_07098_));
 OAI21x1_ASAP7_75t_R _29561_ (.A1(_06913_),
    .A2(_07096_),
    .B(_07098_),
    .Y(_07099_));
 AOI21x1_ASAP7_75t_R _29562_ (.A1(net4539),
    .A2(_06537_),
    .B(net5592),
    .Y(_07100_));
 NAND2x1_ASAP7_75t_R _29563_ (.A(net5340),
    .B(_06618_),
    .Y(_07101_));
 NAND2x1_ASAP7_75t_R _29564_ (.A(_07101_),
    .B(_07100_),
    .Y(_07102_));
 AO21x1_ASAP7_75t_R _29565_ (.A1(_06775_),
    .A2(_06868_),
    .B(net6030),
    .Y(_07103_));
 OA21x2_ASAP7_75t_R _29566_ (.A1(_01380_),
    .A2(net6024),
    .B(net5592),
    .Y(_07104_));
 AOI21x1_ASAP7_75t_R _29567_ (.A1(_07103_),
    .A2(_07104_),
    .B(net5591),
    .Y(_07105_));
 AOI21x1_ASAP7_75t_R _29568_ (.A1(_07102_),
    .A2(_07105_),
    .B(net5588),
    .Y(_07106_));
 AOI21x1_ASAP7_75t_R _29569_ (.A1(_07099_),
    .A2(_07106_),
    .B(net6014),
    .Y(_07107_));
 OAI21x1_ASAP7_75t_R _29570_ (.A1(net6032),
    .A2(_07095_),
    .B(_07107_),
    .Y(_07108_));
 NAND2x1_ASAP7_75t_R _29571_ (.A(_07085_),
    .B(_07108_),
    .Y(_00151_));
 NOR2x1_ASAP7_75t_R _29572_ (.A(net6660),
    .B(_00408_),
    .Y(_07109_));
 XOR2x2_ASAP7_75t_R _29573_ (.A(_12814_),
    .B(net6575),
    .Y(_07110_));
 XOR2x2_ASAP7_75t_R _29574_ (.A(_04380_),
    .B(_12851_),
    .Y(_07111_));
 NAND2x1_ASAP7_75t_R _29575_ (.A(_07110_),
    .B(_07111_),
    .Y(_07112_));
 XNOR2x2_ASAP7_75t_R _29576_ (.A(net6575),
    .B(_12814_),
    .Y(_07113_));
 XOR2x2_ASAP7_75t_R _29577_ (.A(_04380_),
    .B(_12853_),
    .Y(_07114_));
 NAND2x1_ASAP7_75t_R _29578_ (.A(_07113_),
    .B(_07114_),
    .Y(_07115_));
 AOI21x1_ASAP7_75t_R _29579_ (.A1(_07112_),
    .A2(_07115_),
    .B(net6459),
    .Y(_07116_));
 OAI21x1_ASAP7_75t_R _29580_ (.A1(_07109_),
    .A2(net6342),
    .B(net6473),
    .Y(_07117_));
 AND2x2_ASAP7_75t_R _29581_ (.A(net6459),
    .B(_00408_),
    .Y(_07118_));
 NAND2x1_ASAP7_75t_R _29582_ (.A(_07110_),
    .B(_07114_),
    .Y(_07119_));
 NAND2x1_ASAP7_75t_R _29583_ (.A(_07111_),
    .B(_07113_),
    .Y(_07120_));
 AOI21x1_ASAP7_75t_R _29584_ (.A1(_07120_),
    .A2(_07119_),
    .B(net6459),
    .Y(_07121_));
 OAI21x1_ASAP7_75t_R _29585_ (.A1(_07118_),
    .A2(net6341),
    .B(_08913_),
    .Y(_07122_));
 NAND2x1p5_ASAP7_75t_R _29586_ (.A(_07117_),
    .B(_07122_),
    .Y(_07123_));
 AND2x2_ASAP7_75t_R _29588_ (.A(net6459),
    .B(_00409_),
    .Y(_07124_));
 XOR2x2_ASAP7_75t_R _29589_ (.A(_12814_),
    .B(_12838_),
    .Y(_07125_));
 NAND2x1_ASAP7_75t_R _29590_ (.A(_04574_),
    .B(_07125_),
    .Y(_07126_));
 XOR2x2_ASAP7_75t_R _29591_ (.A(_12820_),
    .B(_12838_),
    .Y(_07127_));
 NAND2x1_ASAP7_75t_R _29592_ (.A(net6542),
    .B(_07127_),
    .Y(_07128_));
 AOI21x1_ASAP7_75t_R _29593_ (.A1(_07126_),
    .A2(_07128_),
    .B(net6459),
    .Y(_07129_));
 OAI21x1_ASAP7_75t_R _29594_ (.A1(_07124_),
    .A2(_07129_),
    .B(net6477),
    .Y(_07130_));
 NOR2x1_ASAP7_75t_R _29595_ (.A(net6660),
    .B(_00409_),
    .Y(_07131_));
 NAND2x1_ASAP7_75t_R _29596_ (.A(net6542),
    .B(_07125_),
    .Y(_07132_));
 NAND2x1_ASAP7_75t_R _29597_ (.A(_04574_),
    .B(_07127_),
    .Y(_07133_));
 AOI21x1_ASAP7_75t_R _29598_ (.A1(_07132_),
    .A2(_07133_),
    .B(net6459),
    .Y(_07134_));
 OAI21x1_ASAP7_75t_R _29599_ (.A1(_07131_),
    .A2(_07134_),
    .B(_08908_),
    .Y(_07135_));
 NAND2x1_ASAP7_75t_R _29600_ (.A(_07130_),
    .B(_07135_),
    .Y(_07136_));
 INVx2_ASAP7_75t_R _29601_ (.A(net5585),
    .Y(_01389_));
 XOR2x2_ASAP7_75t_R _29602_ (.A(net6627),
    .B(net6574),
    .Y(_07137_));
 NAND2x1_ASAP7_75t_R _29603_ (.A(net6425),
    .B(_07137_),
    .Y(_07138_));
 XNOR2x2_ASAP7_75t_R _29604_ (.A(net6627),
    .B(net6574),
    .Y(_07139_));
 NAND2x1_ASAP7_75t_R _29605_ (.A(net6546),
    .B(_07139_),
    .Y(_07140_));
 AOI21x1_ASAP7_75t_R _29606_ (.A1(_07138_),
    .A2(_07140_),
    .B(_04423_),
    .Y(_07141_));
 XOR2x2_ASAP7_75t_R _29607_ (.A(net6574),
    .B(net6546),
    .Y(_07142_));
 NAND2x1_ASAP7_75t_R _29608_ (.A(net6627),
    .B(_07142_),
    .Y(_07143_));
 XNOR2x2_ASAP7_75t_R _29609_ (.A(net6574),
    .B(net6546),
    .Y(_07144_));
 NAND2x1_ASAP7_75t_R _29610_ (.A(_01582_),
    .B(_07144_),
    .Y(_07145_));
 AOI21x1_ASAP7_75t_R _29611_ (.A1(_07143_),
    .A2(_07145_),
    .B(net6395),
    .Y(_07146_));
 OAI21x1_ASAP7_75t_R _29612_ (.A1(_07141_),
    .A2(_07146_),
    .B(net6661),
    .Y(_07147_));
 NOR2x1_ASAP7_75t_R _29613_ (.A(net6657),
    .B(_00410_),
    .Y(_07148_));
 INVx1_ASAP7_75t_R _29614_ (.A(_07148_),
    .Y(_07149_));
 NAND3x1_ASAP7_75t_R _29615_ (.A(_07147_),
    .B(_00956_),
    .C(_07149_),
    .Y(_07150_));
 AO21x1_ASAP7_75t_R _29616_ (.A1(_07147_),
    .A2(_07149_),
    .B(_00956_),
    .Y(_07151_));
 NAND2x2_ASAP7_75t_R _29618_ (.A(_07150_),
    .B(_07151_),
    .Y(_07153_));
 INVx1_ASAP7_75t_R _29621_ (.A(_00956_),
    .Y(_07154_));
 NAND3x2_ASAP7_75t_R _29622_ (.B(_07154_),
    .C(_07149_),
    .Y(_07155_),
    .A(_07147_));
 AO21x1_ASAP7_75t_R _29623_ (.A1(_07147_),
    .A2(_07149_),
    .B(_07154_),
    .Y(_07156_));
 NAND2x2_ASAP7_75t_R _29625_ (.A(_07155_),
    .B(_07156_),
    .Y(_07158_));
 XNOR2x2_ASAP7_75t_R _29627_ (.A(net6573),
    .B(_12882_),
    .Y(_07159_));
 NOR2x1_ASAP7_75t_R _29628_ (.A(_07159_),
    .B(_04439_),
    .Y(_07160_));
 XOR2x2_ASAP7_75t_R _29629_ (.A(_12882_),
    .B(net6573),
    .Y(_07161_));
 XNOR2x2_ASAP7_75t_R _29630_ (.A(_04438_),
    .B(_04437_),
    .Y(_07162_));
 OAI21x1_ASAP7_75t_R _29631_ (.A1(_07161_),
    .A2(_07162_),
    .B(net6663),
    .Y(_07163_));
 NAND2x1_ASAP7_75t_R _29632_ (.A(_00529_),
    .B(net6458),
    .Y(_07164_));
 OAI21x1_ASAP7_75t_R _29633_ (.A1(_07160_),
    .A2(_07163_),
    .B(_07164_),
    .Y(_07165_));
 XOR2x2_ASAP7_75t_R _29634_ (.A(_07165_),
    .B(_00959_),
    .Y(_07166_));
 NOR2x1_ASAP7_75t_R _29637_ (.A(net5576),
    .B(net5586),
    .Y(_07169_));
 INVx1_ASAP7_75t_R _29638_ (.A(_07169_),
    .Y(_07170_));
 XOR2x2_ASAP7_75t_R _29639_ (.A(_07165_),
    .B(_08924_),
    .Y(_07171_));
 AOI21x1_ASAP7_75t_R _29642_ (.A1(net6011),
    .A2(net6010),
    .B(_01388_),
    .Y(_07174_));
 XOR2x2_ASAP7_75t_R _29643_ (.A(_12910_),
    .B(net6572),
    .Y(_07175_));
 XOR2x2_ASAP7_75t_R _29644_ (.A(_04449_),
    .B(_07175_),
    .Y(_07176_));
 NOR2x1_ASAP7_75t_R _29645_ (.A(net6657),
    .B(_00523_),
    .Y(_07177_));
 AOI21x1_ASAP7_75t_R _29646_ (.A1(net6659),
    .A2(_07176_),
    .B(_07177_),
    .Y(_07178_));
 XOR2x2_ASAP7_75t_R _29647_ (.A(_07178_),
    .B(_00960_),
    .Y(_07179_));
 AOI21x1_ASAP7_75t_R _29649_ (.A1(net6000),
    .A2(net5077),
    .B(net5997),
    .Y(_07181_));
 OAI21x1_ASAP7_75t_R _29650_ (.A1(net6005),
    .A2(net5078),
    .B(_07181_),
    .Y(_07182_));
 AO21x1_ASAP7_75t_R _29651_ (.A1(net5583),
    .A2(net5582),
    .B(net6001),
    .Y(_07183_));
 NAND2x1_ASAP7_75t_R _29654_ (.A(net5580),
    .B(net5586),
    .Y(_07186_));
 NOR2x1_ASAP7_75t_R _29655_ (.A(net5583),
    .B(_07186_),
    .Y(_07187_));
 NOR2x1_ASAP7_75t_R _29656_ (.A(_07183_),
    .B(_07187_),
    .Y(_07188_));
 XOR2x2_ASAP7_75t_R _29657_ (.A(_00603_),
    .B(_00604_),
    .Y(_07189_));
 XNOR2x2_ASAP7_75t_R _29658_ (.A(net6543),
    .B(_07189_),
    .Y(_07190_));
 XOR2x2_ASAP7_75t_R _29659_ (.A(_07190_),
    .B(_12959_),
    .Y(_07191_));
 NOR2x1_ASAP7_75t_R _29660_ (.A(net6658),
    .B(_00516_),
    .Y(_07192_));
 AO21x1_ASAP7_75t_R _29661_ (.A1(_07191_),
    .A2(net6658),
    .B(_07192_),
    .Y(_07193_));
 XOR2x2_ASAP7_75t_R _29662_ (.A(_07193_),
    .B(_00961_),
    .Y(_07194_));
 OAI21x1_ASAP7_75t_R _29664_ (.A1(_07182_),
    .A2(_07188_),
    .B(net5993),
    .Y(_07196_));
 OAI21x1_ASAP7_75t_R _29666_ (.A1(_07109_),
    .A2(_07116_),
    .B(_08913_),
    .Y(_07198_));
 OAI21x1_ASAP7_75t_R _29667_ (.A1(_07121_),
    .A2(_07118_),
    .B(net6473),
    .Y(_07199_));
 NAND2x2_ASAP7_75t_R _29668_ (.A(_07199_),
    .B(_07198_),
    .Y(_01384_));
 NAND2x2_ASAP7_75t_R _29669_ (.A(net5576),
    .B(net5575),
    .Y(_07200_));
 NOR2x1_ASAP7_75t_R _29670_ (.A(net5580),
    .B(net5575),
    .Y(_07201_));
 AO21x1_ASAP7_75t_R _29671_ (.A1(_07201_),
    .A2(net5584),
    .B(net6006),
    .Y(_07202_));
 INVx1_ASAP7_75t_R _29672_ (.A(_07202_),
    .Y(_07203_));
 INVx1_ASAP7_75t_R _29673_ (.A(_01395_),
    .Y(_07204_));
 AO21x1_ASAP7_75t_R _29674_ (.A1(net6010),
    .A2(net6011),
    .B(_07204_),
    .Y(_07205_));
 INVx1_ASAP7_75t_R _29675_ (.A(net4606),
    .Y(_07206_));
 OAI21x1_ASAP7_75t_R _29677_ (.A1(_07206_),
    .A2(_07183_),
    .B(net5997),
    .Y(_07208_));
 AOI21x1_ASAP7_75t_R _29678_ (.A1(net5331),
    .A2(_07203_),
    .B(_07208_),
    .Y(_07209_));
 NOR2x1_ASAP7_75t_R _29679_ (.A(_07196_),
    .B(_07209_),
    .Y(_07210_));
 INVx1_ASAP7_75t_R _29680_ (.A(_01387_),
    .Y(_07211_));
 AOI21x1_ASAP7_75t_R _29681_ (.A1(net6011),
    .A2(net6010),
    .B(_07211_),
    .Y(_07212_));
 AO21x1_ASAP7_75t_R _29683_ (.A1(net6012),
    .A2(net6013),
    .B(net4821),
    .Y(_07214_));
 NAND2x1_ASAP7_75t_R _29684_ (.A(net6006),
    .B(_07214_),
    .Y(_07215_));
 OAI21x1_ASAP7_75t_R _29685_ (.A1(net4727),
    .A2(_07215_),
    .B(net5996),
    .Y(_07216_));
 AOI21x1_ASAP7_75t_R _29686_ (.A1(net5584),
    .A2(net5587),
    .B(net5577),
    .Y(_07217_));
 NOR2x2_ASAP7_75t_R _29688_ (.A(net5581),
    .B(net5584),
    .Y(_07219_));
 OA21x2_ASAP7_75t_R _29691_ (.A1(_07217_),
    .A2(_07219_),
    .B(net6002),
    .Y(_07222_));
 NOR2x1_ASAP7_75t_R _29692_ (.A(_07216_),
    .B(_07222_),
    .Y(_07223_));
 XOR2x2_ASAP7_75t_R _29693_ (.A(_07178_),
    .B(_09588_),
    .Y(_07224_));
 AOI21x1_ASAP7_75t_R _29695_ (.A1(net5581),
    .A2(net5583),
    .B(net6007),
    .Y(_07226_));
 INVx1_ASAP7_75t_R _29696_ (.A(_07226_),
    .Y(_07227_));
 NAND2x1_ASAP7_75t_R _29697_ (.A(net5991),
    .B(net5076),
    .Y(_07228_));
 AO21x1_ASAP7_75t_R _29699_ (.A1(net5579),
    .A2(net5270),
    .B(_07171_),
    .Y(_07230_));
 NAND2x1_ASAP7_75t_R _29700_ (.A(net5581),
    .B(net5587),
    .Y(_07231_));
 NOR2x1_ASAP7_75t_R _29701_ (.A(net5337),
    .B(_07231_),
    .Y(_07232_));
 NOR2x1_ASAP7_75t_R _29702_ (.A(net5075),
    .B(_07232_),
    .Y(_07233_));
 XNOR2x2_ASAP7_75t_R _29703_ (.A(_00961_),
    .B(_07193_),
    .Y(_07234_));
 OAI21x1_ASAP7_75t_R _29705_ (.A1(_07228_),
    .A2(_07233_),
    .B(net5987),
    .Y(_07236_));
 XOR2x2_ASAP7_75t_R _29706_ (.A(_00604_),
    .B(_00605_),
    .Y(_07237_));
 XOR2x2_ASAP7_75t_R _29707_ (.A(_07237_),
    .B(_12957_),
    .Y(_07238_));
 XOR2x2_ASAP7_75t_R _29708_ (.A(_07238_),
    .B(_12929_),
    .Y(_07239_));
 NOR2x1_ASAP7_75t_R _29709_ (.A(net6665),
    .B(_00508_),
    .Y(_07240_));
 AO21x1_ASAP7_75t_R _29710_ (.A1(_07239_),
    .A2(net6658),
    .B(_07240_),
    .Y(_07241_));
 XOR2x2_ASAP7_75t_R _29711_ (.A(_07241_),
    .B(_00962_),
    .Y(_07242_));
 INVx1_ASAP7_75t_R _29712_ (.A(_07242_),
    .Y(_07243_));
 OAI21x1_ASAP7_75t_R _29714_ (.A1(_07223_),
    .A2(_07236_),
    .B(net5574),
    .Y(_07245_));
 XOR2x2_ASAP7_75t_R _29715_ (.A(_00605_),
    .B(net6624),
    .Y(_07246_));
 XOR2x2_ASAP7_75t_R _29716_ (.A(_07246_),
    .B(_00701_),
    .Y(_07247_));
 XOR2x2_ASAP7_75t_R _29717_ (.A(_07247_),
    .B(_13004_),
    .Y(_07248_));
 NOR2x1_ASAP7_75t_R _29718_ (.A(net6666),
    .B(_00500_),
    .Y(_07249_));
 AO21x1_ASAP7_75t_R _29719_ (.A1(_07248_),
    .A2(net6660),
    .B(_07249_),
    .Y(_07250_));
 XOR2x2_ASAP7_75t_R _29720_ (.A(_07250_),
    .B(_00963_),
    .Y(_07251_));
 OAI21x1_ASAP7_75t_R _29721_ (.A1(_07210_),
    .A2(_07245_),
    .B(net5984),
    .Y(_07252_));
 AOI21x1_ASAP7_75t_R _29722_ (.A1(net6013),
    .A2(net6012),
    .B(_07211_),
    .Y(_07253_));
 NAND2x1_ASAP7_75t_R _29723_ (.A(net6006),
    .B(net4726),
    .Y(_07254_));
 INVx1_ASAP7_75t_R _29724_ (.A(_07254_),
    .Y(_07255_));
 AOI21x1_ASAP7_75t_R _29725_ (.A1(net6011),
    .A2(net6010),
    .B(_01387_),
    .Y(_07256_));
 OA21x2_ASAP7_75t_R _29727_ (.A1(_07201_),
    .A2(_07256_),
    .B(net6002),
    .Y(_07258_));
 OAI21x1_ASAP7_75t_R _29729_ (.A1(_07255_),
    .A2(_07258_),
    .B(net5996),
    .Y(_07260_));
 INVx1_ASAP7_75t_R _29730_ (.A(_01390_),
    .Y(_07261_));
 AO21x1_ASAP7_75t_R _29731_ (.A1(net6012),
    .A2(net6013),
    .B(_07261_),
    .Y(_07262_));
 INVx1_ASAP7_75t_R _29732_ (.A(_01386_),
    .Y(_07263_));
 AO21x1_ASAP7_75t_R _29733_ (.A1(net6010),
    .A2(net6011),
    .B(_07263_),
    .Y(_07264_));
 AO21x1_ASAP7_75t_R _29734_ (.A1(_07262_),
    .A2(net4819),
    .B(net6009),
    .Y(_07265_));
 AO21x1_ASAP7_75t_R _29735_ (.A1(net6012),
    .A2(net6013),
    .B(_07263_),
    .Y(_07266_));
 INVx1_ASAP7_75t_R _29736_ (.A(_07256_),
    .Y(_07267_));
 AO21x1_ASAP7_75t_R _29737_ (.A1(_07266_),
    .A2(_07267_),
    .B(net6002),
    .Y(_07268_));
 AO21x1_ASAP7_75t_R _29739_ (.A1(_07265_),
    .A2(_07268_),
    .B(net5996),
    .Y(_07270_));
 AOI21x1_ASAP7_75t_R _29740_ (.A1(_07260_),
    .A2(_07270_),
    .B(net5987),
    .Y(_07271_));
 INVx2_ASAP7_75t_R _29742_ (.A(net4727),
    .Y(_07273_));
 NAND2x1p5_ASAP7_75t_R _29743_ (.A(_07273_),
    .B(net6003),
    .Y(_07274_));
 NOR2x1_ASAP7_75t_R _29744_ (.A(net5583),
    .B(_07231_),
    .Y(_07275_));
 NOR2x1_ASAP7_75t_R _29745_ (.A(_07274_),
    .B(_07275_),
    .Y(_07276_));
 NOR2x1_ASAP7_75t_R _29747_ (.A(net4820),
    .B(net5581),
    .Y(_07278_));
 NOR2x1_ASAP7_75t_R _29748_ (.A(_07263_),
    .B(net5577),
    .Y(_07279_));
 OAI21x1_ASAP7_75t_R _29751_ (.A1(_07278_),
    .A2(_07279_),
    .B(net6009),
    .Y(_07282_));
 NAND2x1_ASAP7_75t_R _29752_ (.A(net5988),
    .B(_07282_),
    .Y(_07283_));
 OAI21x1_ASAP7_75t_R _29754_ (.A1(_07283_),
    .A2(_07276_),
    .B(_07234_),
    .Y(_07285_));
 NAND2x1_ASAP7_75t_R _29755_ (.A(net5584),
    .B(net5575),
    .Y(_07286_));
 OAI21x1_ASAP7_75t_R _29756_ (.A1(net5581),
    .A2(net5584),
    .B(_07171_),
    .Y(_07287_));
 INVx1_ASAP7_75t_R _29757_ (.A(_07287_),
    .Y(_07288_));
 NOR2x1_ASAP7_75t_R _29758_ (.A(net5576),
    .B(net5583),
    .Y(_07289_));
 AO21x1_ASAP7_75t_R _29759_ (.A1(net5586),
    .A2(net5583),
    .B(net6000),
    .Y(_07290_));
 OAI21x1_ASAP7_75t_R _29760_ (.A1(_07289_),
    .A2(_07290_),
    .B(net5994),
    .Y(_07291_));
 AOI21x1_ASAP7_75t_R _29761_ (.A1(_07286_),
    .A2(_07288_),
    .B(_07291_),
    .Y(_07292_));
 OAI21x1_ASAP7_75t_R _29763_ (.A1(_07285_),
    .A2(_07292_),
    .B(net5985),
    .Y(_07294_));
 NOR2x1_ASAP7_75t_R _29764_ (.A(_07271_),
    .B(_07294_),
    .Y(_07295_));
 INVx1_ASAP7_75t_R _29765_ (.A(_07174_),
    .Y(_07296_));
 OA21x2_ASAP7_75t_R _29766_ (.A1(_07296_),
    .A2(net6000),
    .B(net5997),
    .Y(_07297_));
 NAND2x1_ASAP7_75t_R _29767_ (.A(net5583),
    .B(net5586),
    .Y(_07298_));
 INVx1_ASAP7_75t_R _29768_ (.A(net5328),
    .Y(_07299_));
 AOI21x1_ASAP7_75t_R _29769_ (.A1(net4820),
    .A2(net5581),
    .B(net6009),
    .Y(_07300_));
 INVx1_ASAP7_75t_R _29770_ (.A(_07300_),
    .Y(_07301_));
 AO21x1_ASAP7_75t_R _29771_ (.A1(net5579),
    .A2(_07299_),
    .B(_07301_),
    .Y(_07302_));
 NAND2x1_ASAP7_75t_R _29772_ (.A(_07297_),
    .B(_07302_),
    .Y(_07303_));
 AOI21x1_ASAP7_75t_R _29773_ (.A1(net5030),
    .A2(net5582),
    .B(net5999),
    .Y(_07304_));
 OA21x2_ASAP7_75t_R _29774_ (.A1(net5328),
    .A2(net5582),
    .B(net4818),
    .Y(_07305_));
 INVx1_ASAP7_75t_R _29775_ (.A(_07181_),
    .Y(_07306_));
 OA21x2_ASAP7_75t_R _29776_ (.A1(_07305_),
    .A2(_07306_),
    .B(net5987),
    .Y(_07307_));
 AOI21x1_ASAP7_75t_R _29779_ (.A1(net6013),
    .A2(net6012),
    .B(_01387_),
    .Y(_07310_));
 NOR2x1p5_ASAP7_75t_R _29780_ (.A(net6007),
    .B(_07310_),
    .Y(_07311_));
 AOI21x1_ASAP7_75t_R _29781_ (.A1(_01403_),
    .A2(net6004),
    .B(_07311_),
    .Y(_07312_));
 OAI21x1_ASAP7_75t_R _29783_ (.A1(net5989),
    .A2(_07312_),
    .B(net5993),
    .Y(_07314_));
 AO21x1_ASAP7_75t_R _29784_ (.A1(net6010),
    .A2(net6011),
    .B(_01386_),
    .Y(_07315_));
 INVx1_ASAP7_75t_R _29785_ (.A(_07315_),
    .Y(_07316_));
 NOR2x1_ASAP7_75t_R _29786_ (.A(net5271),
    .B(net5576),
    .Y(_07317_));
 NAND2x1_ASAP7_75t_R _29787_ (.A(net5999),
    .B(_07317_),
    .Y(_07318_));
 OAI21x1_ASAP7_75t_R _29788_ (.A1(_07316_),
    .A2(_07183_),
    .B(_07318_),
    .Y(_07319_));
 AO21x1_ASAP7_75t_R _29790_ (.A1(net5586),
    .A2(net5583),
    .B(net5582),
    .Y(_07321_));
 AOI21x1_ASAP7_75t_R _29791_ (.A1(net6013),
    .A2(net6012),
    .B(_01393_),
    .Y(_07322_));
 AOI21x1_ASAP7_75t_R _29792_ (.A1(net6001),
    .A2(net5074),
    .B(net5994),
    .Y(_07323_));
 OAI21x1_ASAP7_75t_R _29793_ (.A1(net6005),
    .A2(_07321_),
    .B(_07323_),
    .Y(_07324_));
 NOR2x1_ASAP7_75t_R _29794_ (.A(_07319_),
    .B(_07324_),
    .Y(_07325_));
 OAI21x1_ASAP7_75t_R _29796_ (.A1(_07314_),
    .A2(_07325_),
    .B(net5985),
    .Y(_07327_));
 AOI21x1_ASAP7_75t_R _29797_ (.A1(_07303_),
    .A2(_07307_),
    .B(_07327_),
    .Y(_07328_));
 OA21x2_ASAP7_75t_R _29798_ (.A1(_07187_),
    .A2(net5334),
    .B(_07323_),
    .Y(_07329_));
 AO21x1_ASAP7_75t_R _29799_ (.A1(net5074),
    .A2(net6003),
    .B(net5991),
    .Y(_07330_));
 AO21x1_ASAP7_75t_R _29800_ (.A1(net6010),
    .A2(net6011),
    .B(_01391_),
    .Y(_07331_));
 INVx1_ASAP7_75t_R _29802_ (.A(net4817),
    .Y(_07333_));
 NOR2x1_ASAP7_75t_R _29803_ (.A(net6003),
    .B(_07212_),
    .Y(_07334_));
 AO21x1_ASAP7_75t_R _29804_ (.A1(net6003),
    .A2(_07333_),
    .B(_07334_),
    .Y(_07335_));
 OAI21x1_ASAP7_75t_R _29805_ (.A1(_07330_),
    .A2(_07335_),
    .B(net5993),
    .Y(_07336_));
 NOR2x1_ASAP7_75t_R _29806_ (.A(_07329_),
    .B(_07336_),
    .Y(_07337_));
 OAI21x1_ASAP7_75t_R _29807_ (.A1(net5077),
    .A2(_07279_),
    .B(net6000),
    .Y(_07338_));
 INVx1_ASAP7_75t_R _29808_ (.A(_07338_),
    .Y(_07339_));
 NAND2x1_ASAP7_75t_R _29809_ (.A(net5997),
    .B(net5075),
    .Y(_07340_));
 OAI21x1_ASAP7_75t_R _29810_ (.A1(_07339_),
    .A2(_07340_),
    .B(net5987),
    .Y(_07341_));
 AOI21x1_ASAP7_75t_R _29811_ (.A1(net5578),
    .A2(net5587),
    .B(net6009),
    .Y(_07342_));
 INVx1_ASAP7_75t_R _29812_ (.A(net5327),
    .Y(_07343_));
 NOR2x1_ASAP7_75t_R _29813_ (.A(net4992),
    .B(_07343_),
    .Y(_07344_));
 NAND2x1_ASAP7_75t_R _29814_ (.A(net5580),
    .B(net5584),
    .Y(_07345_));
 INVx1_ASAP7_75t_R _29815_ (.A(_07345_),
    .Y(_07346_));
 AO21x1_ASAP7_75t_R _29816_ (.A1(net5581),
    .A2(net4820),
    .B(net6002),
    .Y(_07347_));
 OAI21x1_ASAP7_75t_R _29818_ (.A1(_07346_),
    .A2(_07347_),
    .B(net5988),
    .Y(_07349_));
 NOR2x1_ASAP7_75t_R _29819_ (.A(_07344_),
    .B(_07349_),
    .Y(_07350_));
 OAI21x1_ASAP7_75t_R _29820_ (.A1(_07341_),
    .A2(_07350_),
    .B(net5574),
    .Y(_07351_));
 INVx1_ASAP7_75t_R _29821_ (.A(_07251_),
    .Y(_07352_));
 OAI21x1_ASAP7_75t_R _29822_ (.A1(_07337_),
    .A2(_07351_),
    .B(_07352_),
    .Y(_07353_));
 OAI22x1_ASAP7_75t_R _29823_ (.A1(_07252_),
    .A2(_07295_),
    .B1(_07328_),
    .B2(_07353_),
    .Y(_00152_));
 NOR2x1_ASAP7_75t_R _29824_ (.A(net6003),
    .B(_07275_),
    .Y(_07354_));
 NAND2x1_ASAP7_75t_R _29825_ (.A(net6000),
    .B(_07205_),
    .Y(_07355_));
 INVx1_ASAP7_75t_R _29826_ (.A(_07355_),
    .Y(_07356_));
 INVx1_ASAP7_75t_R _29827_ (.A(_01388_),
    .Y(_07357_));
 AO21x1_ASAP7_75t_R _29828_ (.A1(net6012),
    .A2(net6013),
    .B(_07357_),
    .Y(_07358_));
 AO21x1_ASAP7_75t_R _29830_ (.A1(_07356_),
    .A2(net4815),
    .B(net5987),
    .Y(_07360_));
 AO21x1_ASAP7_75t_R _29831_ (.A1(net4725),
    .A2(_07354_),
    .B(_07360_),
    .Y(_07361_));
 NAND2x1_ASAP7_75t_R _29832_ (.A(net6000),
    .B(_07289_),
    .Y(_07362_));
 OA21x2_ASAP7_75t_R _29833_ (.A1(net6005),
    .A2(_07296_),
    .B(net5987),
    .Y(_07363_));
 NAND2x1_ASAP7_75t_R _29834_ (.A(_07362_),
    .B(_07363_),
    .Y(_07364_));
 NOR2x1p5_ASAP7_75t_R _29835_ (.A(net6003),
    .B(_07253_),
    .Y(_07365_));
 AND2x2_ASAP7_75t_R _29836_ (.A(_07365_),
    .B(_07315_),
    .Y(_07366_));
 OA21x2_ASAP7_75t_R _29837_ (.A1(_07364_),
    .A2(_07366_),
    .B(net5994),
    .Y(_07367_));
 INVx1_ASAP7_75t_R _29838_ (.A(net5075),
    .Y(_07368_));
 NOR2x1_ASAP7_75t_R _29839_ (.A(_01386_),
    .B(net5579),
    .Y(_07369_));
 NOR2x1_ASAP7_75t_R _29840_ (.A(_07369_),
    .B(_07287_),
    .Y(_07370_));
 AOI211x1_ASAP7_75t_R _29841_ (.A1(_07368_),
    .A2(net5078),
    .B(_07370_),
    .C(net5993),
    .Y(_07371_));
 INVx2_ASAP7_75t_R _29842_ (.A(_07334_),
    .Y(_07372_));
 NAND2x1p5_ASAP7_75t_R _29843_ (.A(net5993),
    .B(net4450),
    .Y(_07373_));
 NOR2x1_ASAP7_75t_R _29844_ (.A(net5076),
    .B(_07187_),
    .Y(_07374_));
 OAI21x1_ASAP7_75t_R _29845_ (.A1(_07374_),
    .A2(_07373_),
    .B(net5991),
    .Y(_07375_));
 OAI21x1_ASAP7_75t_R _29846_ (.A1(_07371_),
    .A2(_07375_),
    .B(net5574),
    .Y(_07376_));
 AOI21x1_ASAP7_75t_R _29847_ (.A1(_07361_),
    .A2(_07367_),
    .B(_07376_),
    .Y(_07377_));
 NOR2x1_ASAP7_75t_R _29848_ (.A(net5584),
    .B(net5575),
    .Y(_07378_));
 NAND2x1_ASAP7_75t_R _29849_ (.A(net5578),
    .B(_07378_),
    .Y(_07379_));
 AND2x2_ASAP7_75t_R _29850_ (.A(net6008),
    .B(_01400_),
    .Y(_07380_));
 AOI22x1_ASAP7_75t_R _29851_ (.A1(_07379_),
    .A2(net4604),
    .B1(net5992),
    .B2(_07380_),
    .Y(_07381_));
 OAI21x1_ASAP7_75t_R _29852_ (.A1(net5996),
    .A2(_07381_),
    .B(net5985),
    .Y(_07382_));
 AOI21x1_ASAP7_75t_R _29853_ (.A1(net5587),
    .A2(net5336),
    .B(net5581),
    .Y(_07383_));
 OAI21x1_ASAP7_75t_R _29854_ (.A1(_07217_),
    .A2(_07383_),
    .B(net6008),
    .Y(_07384_));
 AO21x1_ASAP7_75t_R _29855_ (.A1(net5581),
    .A2(_07263_),
    .B(net6008),
    .Y(_07385_));
 OA21x2_ASAP7_75t_R _29856_ (.A1(_07385_),
    .A2(_07346_),
    .B(net5986),
    .Y(_07386_));
 NOR2x1_ASAP7_75t_R _29857_ (.A(_07201_),
    .B(_07287_),
    .Y(_07387_));
 OAI21x1_ASAP7_75t_R _29859_ (.A1(net5335),
    .A2(_07230_),
    .B(net5992),
    .Y(_07389_));
 OAI21x1_ASAP7_75t_R _29860_ (.A1(_07387_),
    .A2(_07389_),
    .B(net5995),
    .Y(_07390_));
 AOI21x1_ASAP7_75t_R _29861_ (.A1(_07384_),
    .A2(_07386_),
    .B(_07390_),
    .Y(_07391_));
 OAI21x1_ASAP7_75t_R _29862_ (.A1(_07382_),
    .A2(_07391_),
    .B(net5984),
    .Y(_07392_));
 AO21x1_ASAP7_75t_R _29863_ (.A1(net5587),
    .A2(net5581),
    .B(net5998),
    .Y(_07393_));
 NAND2x1_ASAP7_75t_R _29864_ (.A(net5331),
    .B(_07393_),
    .Y(_07394_));
 OAI21x1_ASAP7_75t_R _29865_ (.A1(_07330_),
    .A2(_07394_),
    .B(net5993),
    .Y(_07395_));
 NAND2x1_ASAP7_75t_R _29866_ (.A(_07205_),
    .B(_07365_),
    .Y(_07396_));
 INVx1_ASAP7_75t_R _29867_ (.A(_07396_),
    .Y(_07397_));
 NOR2x1_ASAP7_75t_R _29868_ (.A(_07397_),
    .B(_07324_),
    .Y(_07398_));
 OAI21x1_ASAP7_75t_R _29869_ (.A1(_07395_),
    .A2(_07398_),
    .B(net5985),
    .Y(_07399_));
 OAI21x1_ASAP7_75t_R _29870_ (.A1(net5577),
    .A2(net5584),
    .B(net6002),
    .Y(_07400_));
 AOI21x1_ASAP7_75t_R _29871_ (.A1(net5270),
    .A2(net5579),
    .B(_07400_),
    .Y(_07401_));
 OAI21x1_ASAP7_75t_R _29872_ (.A1(net4727),
    .A2(_07183_),
    .B(net5994),
    .Y(_07402_));
 OAI21x1_ASAP7_75t_R _29873_ (.A1(_07401_),
    .A2(_07402_),
    .B(net5987),
    .Y(_07403_));
 NOR2x1_ASAP7_75t_R _29874_ (.A(net5580),
    .B(net5998),
    .Y(_07404_));
 AO21x1_ASAP7_75t_R _29875_ (.A1(net5327),
    .A2(_07286_),
    .B(net5994),
    .Y(_07405_));
 AOI21x1_ASAP7_75t_R _29876_ (.A1(net5328),
    .A2(_07404_),
    .B(_07405_),
    .Y(_07406_));
 NOR2x1_ASAP7_75t_R _29877_ (.A(_07403_),
    .B(_07406_),
    .Y(_07407_));
 OAI21x1_ASAP7_75t_R _29878_ (.A1(_07399_),
    .A2(_07407_),
    .B(_07352_),
    .Y(_07408_));
 INVx1_ASAP7_75t_R _29879_ (.A(_07322_),
    .Y(_07409_));
 NAND2x1_ASAP7_75t_R _29880_ (.A(net6007),
    .B(_07409_),
    .Y(_07410_));
 NOR2x1_ASAP7_75t_R _29881_ (.A(net4727),
    .B(_07410_),
    .Y(_07411_));
 INVx1_ASAP7_75t_R _29882_ (.A(_07264_),
    .Y(_07412_));
 NOR2x1_ASAP7_75t_R _29883_ (.A(_07412_),
    .B(_07400_),
    .Y(_07413_));
 OA21x2_ASAP7_75t_R _29884_ (.A1(_07411_),
    .A2(_07413_),
    .B(_07179_),
    .Y(_07414_));
 AO21x1_ASAP7_75t_R _29885_ (.A1(_07311_),
    .A2(net5325),
    .B(_07179_),
    .Y(_07415_));
 OA21x2_ASAP7_75t_R _29886_ (.A1(_07346_),
    .A2(_07378_),
    .B(net6009),
    .Y(_07416_));
 OAI21x1_ASAP7_75t_R _29887_ (.A1(_07415_),
    .A2(_07416_),
    .B(net5992),
    .Y(_07417_));
 NOR2x1_ASAP7_75t_R _29888_ (.A(_07414_),
    .B(_07417_),
    .Y(_07418_));
 INVx1_ASAP7_75t_R _29889_ (.A(net5331),
    .Y(_07419_));
 OAI21x1_ASAP7_75t_R _29890_ (.A1(_07419_),
    .A2(_07215_),
    .B(net5996),
    .Y(_07420_));
 AND2x2_ASAP7_75t_R _29891_ (.A(_07383_),
    .B(net6002),
    .Y(_07421_));
 OAI21x1_ASAP7_75t_R _29892_ (.A1(_07420_),
    .A2(_07421_),
    .B(_07234_),
    .Y(_07422_));
 AO21x1_ASAP7_75t_R _29893_ (.A1(net6010),
    .A2(net6011),
    .B(net5269),
    .Y(_07423_));
 OAI21x1_ASAP7_75t_R _29894_ (.A1(net6006),
    .A2(_07423_),
    .B(net5991),
    .Y(_07424_));
 AOI21x1_ASAP7_75t_R _29895_ (.A1(net4725),
    .A2(_07354_),
    .B(_07424_),
    .Y(_07425_));
 OAI21x1_ASAP7_75t_R _29896_ (.A1(_07422_),
    .A2(_07425_),
    .B(net5574),
    .Y(_07426_));
 NOR2x1_ASAP7_75t_R _29897_ (.A(_07418_),
    .B(_07426_),
    .Y(_07427_));
 OAI22x1_ASAP7_75t_R _29898_ (.A1(_07377_),
    .A2(_07392_),
    .B1(_07408_),
    .B2(_07427_),
    .Y(_00153_));
 AOI21x1_ASAP7_75t_R _29899_ (.A1(net6013),
    .A2(net6012),
    .B(_01395_),
    .Y(_07428_));
 INVx1_ASAP7_75t_R _29900_ (.A(_07428_),
    .Y(_07429_));
 AO21x1_ASAP7_75t_R _29901_ (.A1(_07423_),
    .A2(_07429_),
    .B(net6004),
    .Y(_07430_));
 OAI21x1_ASAP7_75t_R _29902_ (.A1(net5576),
    .A2(net5583),
    .B(net5586),
    .Y(_07431_));
 NAND2x1_ASAP7_75t_R _29903_ (.A(net6004),
    .B(_07431_),
    .Y(_07432_));
 AO21x1_ASAP7_75t_R _29904_ (.A1(_07430_),
    .A2(_07432_),
    .B(net5989),
    .Y(_07433_));
 NOR2x1_ASAP7_75t_R _29905_ (.A(_07219_),
    .B(_07410_),
    .Y(_07434_));
 AOI21x1_ASAP7_75t_R _29907_ (.A1(net5331),
    .A2(_07434_),
    .B(net5994),
    .Y(_07436_));
 OAI21x1_ASAP7_75t_R _29908_ (.A1(net4992),
    .A2(_07343_),
    .B(_07436_),
    .Y(_07437_));
 AOI21x1_ASAP7_75t_R _29909_ (.A1(_07433_),
    .A2(_07437_),
    .B(net5987),
    .Y(_07438_));
 NOR2x1p5_ASAP7_75t_R _29910_ (.A(net6009),
    .B(_07256_),
    .Y(_07439_));
 AND2x2_ASAP7_75t_R _29911_ (.A(_07170_),
    .B(_07439_),
    .Y(_07440_));
 AO21x1_ASAP7_75t_R _29912_ (.A1(net5581),
    .A2(_07357_),
    .B(net5998),
    .Y(_07441_));
 NOR2x1_ASAP7_75t_R _29913_ (.A(_07219_),
    .B(_07441_),
    .Y(_07442_));
 OA21x2_ASAP7_75t_R _29914_ (.A1(_07440_),
    .A2(_07442_),
    .B(net5994),
    .Y(_07443_));
 NAND2x1_ASAP7_75t_R _29915_ (.A(net5990),
    .B(_07202_),
    .Y(_07444_));
 OA211x2_ASAP7_75t_R _29916_ (.A1(net5330),
    .A2(net5584),
    .B(net6007),
    .C(_07205_),
    .Y(_07445_));
 OAI21x1_ASAP7_75t_R _29917_ (.A1(_07444_),
    .A2(_07445_),
    .B(net5987),
    .Y(_07446_));
 OAI21x1_ASAP7_75t_R _29918_ (.A1(_07443_),
    .A2(_07446_),
    .B(net5985),
    .Y(_07447_));
 NOR2x1_ASAP7_75t_R _29919_ (.A(_07438_),
    .B(_07447_),
    .Y(_07448_));
 NAND2x1_ASAP7_75t_R _29920_ (.A(net5999),
    .B(_07429_),
    .Y(_07449_));
 OAI21x1_ASAP7_75t_R _29921_ (.A1(_07219_),
    .A2(_07410_),
    .B(_07449_),
    .Y(_07450_));
 NOR2x1_ASAP7_75t_R _29922_ (.A(_07166_),
    .B(net4817),
    .Y(_07451_));
 NOR2x1_ASAP7_75t_R _29923_ (.A(net5988),
    .B(_07451_),
    .Y(_07452_));
 AO21x1_ASAP7_75t_R _29924_ (.A1(_07450_),
    .A2(_07452_),
    .B(net5986),
    .Y(_07453_));
 AO21x1_ASAP7_75t_R _29925_ (.A1(net5332),
    .A2(net4814),
    .B(net6003),
    .Y(_07454_));
 OAI21x1_ASAP7_75t_R _29926_ (.A1(net5074),
    .A2(_07333_),
    .B(net6003),
    .Y(_07455_));
 AND3x1_ASAP7_75t_R _29927_ (.A(_07454_),
    .B(net5990),
    .C(_07455_),
    .Y(_07456_));
 NOR2x1_ASAP7_75t_R _29928_ (.A(_07453_),
    .B(_07456_),
    .Y(_07457_));
 AOI21x1_ASAP7_75t_R _29929_ (.A1(net5030),
    .A2(net5581),
    .B(_07166_),
    .Y(_07458_));
 NAND2x1_ASAP7_75t_R _29930_ (.A(_07345_),
    .B(_07458_),
    .Y(_07459_));
 INVx1_ASAP7_75t_R _29931_ (.A(net4726),
    .Y(_07460_));
 AO21x1_ASAP7_75t_R _29932_ (.A1(_07460_),
    .A2(_07267_),
    .B(net6002),
    .Y(_07461_));
 AOI21x1_ASAP7_75t_R _29933_ (.A1(_07459_),
    .A2(_07461_),
    .B(net5996),
    .Y(_07462_));
 AOI21x1_ASAP7_75t_R _29934_ (.A1(net5582),
    .A2(net5575),
    .B(_07171_),
    .Y(_07463_));
 OAI21x1_ASAP7_75t_R _29935_ (.A1(net4813),
    .A2(_07287_),
    .B(_07179_),
    .Y(_07464_));
 AOI21x1_ASAP7_75t_R _29936_ (.A1(net4817),
    .A2(net5324),
    .B(_07464_),
    .Y(_07465_));
 OAI21x1_ASAP7_75t_R _29937_ (.A1(_07462_),
    .A2(_07465_),
    .B(net5987),
    .Y(_07466_));
 NAND2x1_ASAP7_75t_R _29938_ (.A(net5574),
    .B(_07466_),
    .Y(_07467_));
 OAI21x1_ASAP7_75t_R _29939_ (.A1(_07457_),
    .A2(_07467_),
    .B(net5984),
    .Y(_07468_));
 NAND2x1_ASAP7_75t_R _29940_ (.A(_01402_),
    .B(net6004),
    .Y(_07469_));
 OAI21x1_ASAP7_75t_R _29941_ (.A1(net6007),
    .A2(_07232_),
    .B(_07469_),
    .Y(_07470_));
 OA21x2_ASAP7_75t_R _29942_ (.A1(_01404_),
    .A2(net6004),
    .B(net5997),
    .Y(_07471_));
 AOI21x1_ASAP7_75t_R _29943_ (.A1(_07471_),
    .A2(_07432_),
    .B(net5987),
    .Y(_07472_));
 OAI21x1_ASAP7_75t_R _29944_ (.A1(net5997),
    .A2(_07470_),
    .B(_07472_),
    .Y(_07473_));
 AND2x2_ASAP7_75t_R _29945_ (.A(_01393_),
    .B(_01388_),
    .Y(_07474_));
 AO21x1_ASAP7_75t_R _29946_ (.A1(net5578),
    .A2(_07474_),
    .B(net6002),
    .Y(_07475_));
 NOR2x1_ASAP7_75t_R _29947_ (.A(net4810),
    .B(_07275_),
    .Y(_07476_));
 OAI21x1_ASAP7_75t_R _29948_ (.A1(_07301_),
    .A2(_07187_),
    .B(net5994),
    .Y(_07477_));
 AO21x1_ASAP7_75t_R _29949_ (.A1(net4814),
    .A2(_07267_),
    .B(net6003),
    .Y(_07478_));
 OA21x2_ASAP7_75t_R _29950_ (.A1(net4819),
    .A2(net6006),
    .B(net5988),
    .Y(_07479_));
 AOI21x1_ASAP7_75t_R _29951_ (.A1(_07478_),
    .A2(_07479_),
    .B(net5992),
    .Y(_07480_));
 OAI21x1_ASAP7_75t_R _29952_ (.A1(_07476_),
    .A2(_07477_),
    .B(_07480_),
    .Y(_07481_));
 AOI21x1_ASAP7_75t_R _29953_ (.A1(_07473_),
    .A2(_07481_),
    .B(net5574),
    .Y(_07482_));
 AND2x2_ASAP7_75t_R _29954_ (.A(net5324),
    .B(net5325),
    .Y(_07483_));
 INVx1_ASAP7_75t_R _29955_ (.A(net4992),
    .Y(_07484_));
 AO21x1_ASAP7_75t_R _29956_ (.A1(net5327),
    .A2(_07484_),
    .B(net5990),
    .Y(_07485_));
 OA21x2_ASAP7_75t_R _29957_ (.A1(_01403_),
    .A2(net6004),
    .B(net5988),
    .Y(_07486_));
 OAI21x1_ASAP7_75t_R _29958_ (.A1(net5582),
    .A2(net5328),
    .B(_07365_),
    .Y(_07487_));
 AOI21x1_ASAP7_75t_R _29959_ (.A1(_07486_),
    .A2(_07487_),
    .B(_07194_),
    .Y(_07488_));
 OAI21x1_ASAP7_75t_R _29960_ (.A1(_07483_),
    .A2(_07485_),
    .B(_07488_),
    .Y(_07489_));
 NOR2x1_ASAP7_75t_R _29961_ (.A(net6002),
    .B(_07278_),
    .Y(_07490_));
 AOI22x1_ASAP7_75t_R _29962_ (.A1(_07490_),
    .A2(_07484_),
    .B1(net5326),
    .B2(_07266_),
    .Y(_07491_));
 NAND2x1_ASAP7_75t_R _29963_ (.A(_01400_),
    .B(net6002),
    .Y(_07492_));
 AOI21x1_ASAP7_75t_R _29964_ (.A1(net5577),
    .A2(net5587),
    .B(net6002),
    .Y(_07493_));
 AOI21x1_ASAP7_75t_R _29965_ (.A1(_07286_),
    .A2(_07493_),
    .B(_07179_),
    .Y(_07494_));
 AOI21x1_ASAP7_75t_R _29966_ (.A1(_07492_),
    .A2(_07494_),
    .B(net5986),
    .Y(_07495_));
 OAI21x1_ASAP7_75t_R _29967_ (.A1(net5988),
    .A2(_07491_),
    .B(_07495_),
    .Y(_07496_));
 AOI21x1_ASAP7_75t_R _29968_ (.A1(_07489_),
    .A2(_07496_),
    .B(net5985),
    .Y(_07497_));
 OAI21x1_ASAP7_75t_R _29969_ (.A1(_07482_),
    .A2(_07497_),
    .B(net5573),
    .Y(_07498_));
 OAI21x1_ASAP7_75t_R _29970_ (.A1(_07448_),
    .A2(_07468_),
    .B(_07498_),
    .Y(_00154_));
 NAND2x1_ASAP7_75t_R _29971_ (.A(net5031),
    .B(net5581),
    .Y(_07499_));
 NAND2x1_ASAP7_75t_R _29972_ (.A(_07474_),
    .B(net5578),
    .Y(_07500_));
 AND3x1_ASAP7_75t_R _29973_ (.A(_07499_),
    .B(_07500_),
    .C(net6009),
    .Y(_07501_));
 AOI21x1_ASAP7_75t_R _29974_ (.A1(net4604),
    .A2(_07379_),
    .B(_07501_),
    .Y(_07502_));
 AND2x2_ASAP7_75t_R _29975_ (.A(_07464_),
    .B(net5992),
    .Y(_07503_));
 OAI21x1_ASAP7_75t_R _29976_ (.A1(net5996),
    .A2(_07502_),
    .B(_07503_),
    .Y(_07504_));
 NOR2x1_ASAP7_75t_R _29977_ (.A(_07316_),
    .B(_07183_),
    .Y(_07505_));
 OA21x2_ASAP7_75t_R _29978_ (.A1(_07331_),
    .A2(net5998),
    .B(_07179_),
    .Y(_07506_));
 INVx1_ASAP7_75t_R _29979_ (.A(_07506_),
    .Y(_07507_));
 INVx1_ASAP7_75t_R _29980_ (.A(_07404_),
    .Y(_07508_));
 OAI21x1_ASAP7_75t_R _29981_ (.A1(_07256_),
    .A2(net4813),
    .B(net5998),
    .Y(_07509_));
 OAI21x1_ASAP7_75t_R _29982_ (.A1(net5337),
    .A2(_07508_),
    .B(_07509_),
    .Y(_07510_));
 OAI22x1_ASAP7_75t_R _29983_ (.A1(_07405_),
    .A2(_07505_),
    .B1(_07507_),
    .B2(_07510_),
    .Y(_07511_));
 AOI21x1_ASAP7_75t_R _29984_ (.A1(net5987),
    .A2(_07511_),
    .B(net5985),
    .Y(_07512_));
 NAND2x1_ASAP7_75t_R _29985_ (.A(net5332),
    .B(_07300_),
    .Y(_07513_));
 AOI21x1_ASAP7_75t_R _29986_ (.A1(_07254_),
    .A2(_07513_),
    .B(_07234_),
    .Y(_07514_));
 NAND2x1_ASAP7_75t_R _29987_ (.A(net6003),
    .B(net4727),
    .Y(_07515_));
 OAI21x1_ASAP7_75t_R _29988_ (.A1(net5992),
    .A2(_07515_),
    .B(_07297_),
    .Y(_07516_));
 OAI21x1_ASAP7_75t_R _29989_ (.A1(_07514_),
    .A2(_07516_),
    .B(net5985),
    .Y(_07517_));
 OA21x2_ASAP7_75t_R _29990_ (.A1(net6002),
    .A2(net4816),
    .B(_07234_),
    .Y(_07518_));
 NAND2x1_ASAP7_75t_R _29991_ (.A(_07459_),
    .B(_07518_),
    .Y(_07519_));
 INVx1_ASAP7_75t_R _29992_ (.A(_07214_),
    .Y(_07520_));
 AOI21x1_ASAP7_75t_R _29993_ (.A1(_07226_),
    .A2(_07273_),
    .B(_07234_),
    .Y(_07521_));
 OAI21x1_ASAP7_75t_R _29994_ (.A1(_07520_),
    .A2(_07475_),
    .B(_07521_),
    .Y(_07522_));
 AOI21x1_ASAP7_75t_R _29995_ (.A1(_07522_),
    .A2(_07519_),
    .B(net5996),
    .Y(_07523_));
 NOR2x1_ASAP7_75t_R _29996_ (.A(_07517_),
    .B(_07523_),
    .Y(_07524_));
 AOI21x1_ASAP7_75t_R _29997_ (.A1(_07504_),
    .A2(_07512_),
    .B(_07524_),
    .Y(_07525_));
 OA21x2_ASAP7_75t_R _29998_ (.A1(_07387_),
    .A2(_07255_),
    .B(net5996),
    .Y(_07526_));
 OA21x2_ASAP7_75t_R _29999_ (.A1(_07299_),
    .A2(_07287_),
    .B(net5990),
    .Y(_07527_));
 NAND2x1_ASAP7_75t_R _30000_ (.A(net4533),
    .B(net5324),
    .Y(_07528_));
 AO21x1_ASAP7_75t_R _30001_ (.A1(_07527_),
    .A2(_07528_),
    .B(net5987),
    .Y(_07529_));
 NOR2x1_ASAP7_75t_R _30002_ (.A(_07278_),
    .B(_07400_),
    .Y(_07530_));
 AND2x2_ASAP7_75t_R _30003_ (.A(_07365_),
    .B(net4819),
    .Y(_07531_));
 OAI21x1_ASAP7_75t_R _30004_ (.A1(_07530_),
    .A2(_07531_),
    .B(_07179_),
    .Y(_07532_));
 AO21x1_ASAP7_75t_R _30005_ (.A1(net6010),
    .A2(net6011),
    .B(_01395_),
    .Y(_07533_));
 AO21x1_ASAP7_75t_R _30006_ (.A1(_07533_),
    .A2(net4814),
    .B(net6002),
    .Y(_07534_));
 AOI21x1_ASAP7_75t_R _30007_ (.A1(_07439_),
    .A2(_07170_),
    .B(net5994),
    .Y(_07535_));
 AOI21x1_ASAP7_75t_R _30008_ (.A1(_07534_),
    .A2(_07535_),
    .B(net5992),
    .Y(_07536_));
 AOI21x1_ASAP7_75t_R _30009_ (.A1(_07532_),
    .A2(_07536_),
    .B(net5574),
    .Y(_07537_));
 OAI21x1_ASAP7_75t_R _30010_ (.A1(_07526_),
    .A2(_07529_),
    .B(_07537_),
    .Y(_07538_));
 OA21x2_ASAP7_75t_R _30011_ (.A1(net5582),
    .A2(net6000),
    .B(net5989),
    .Y(_07539_));
 NAND2x1_ASAP7_75t_R _30012_ (.A(net5579),
    .B(net5337),
    .Y(_07540_));
 NAND2x1_ASAP7_75t_R _30013_ (.A(net5328),
    .B(_07540_),
    .Y(_07541_));
 AOI21x1_ASAP7_75t_R _30014_ (.A1(_07539_),
    .A2(_07541_),
    .B(net5987),
    .Y(_07542_));
 NAND2x1_ASAP7_75t_R _30015_ (.A(_07499_),
    .B(_07439_),
    .Y(_07543_));
 OA21x2_ASAP7_75t_R _30016_ (.A1(net5578),
    .A2(net4821),
    .B(net6009),
    .Y(_07544_));
 AOI21x1_ASAP7_75t_R _30017_ (.A1(net5331),
    .A2(_07544_),
    .B(net5988),
    .Y(_07545_));
 NAND2x1_ASAP7_75t_R _30018_ (.A(_07543_),
    .B(_07545_),
    .Y(_07546_));
 AOI21x1_ASAP7_75t_R _30019_ (.A1(_07542_),
    .A2(_07546_),
    .B(net5985),
    .Y(_07547_));
 INVx1_ASAP7_75t_R _30020_ (.A(_07311_),
    .Y(_07548_));
 NOR2x1_ASAP7_75t_R _30021_ (.A(_07548_),
    .B(_07383_),
    .Y(_07549_));
 AO21x1_ASAP7_75t_R _30022_ (.A1(net5580),
    .A2(_01390_),
    .B(net5998),
    .Y(_07550_));
 OAI21x1_ASAP7_75t_R _30023_ (.A1(_07217_),
    .A2(_07550_),
    .B(net5988),
    .Y(_07551_));
 NOR2x1_ASAP7_75t_R _30024_ (.A(_07549_),
    .B(_07551_),
    .Y(_07552_));
 AO21x1_ASAP7_75t_R _30025_ (.A1(_07262_),
    .A2(_07273_),
    .B(net6009),
    .Y(_07553_));
 OAI21x1_ASAP7_75t_R _30026_ (.A1(_07289_),
    .A2(_07299_),
    .B(net6006),
    .Y(_07554_));
 AOI21x1_ASAP7_75t_R _30027_ (.A1(_07553_),
    .A2(_07554_),
    .B(net5988),
    .Y(_07555_));
 OAI21x1_ASAP7_75t_R _30028_ (.A1(_07552_),
    .A2(_07555_),
    .B(net5987),
    .Y(_07556_));
 AOI21x1_ASAP7_75t_R _30029_ (.A1(_07547_),
    .A2(_07556_),
    .B(net5984),
    .Y(_07557_));
 NAND2x1_ASAP7_75t_R _30030_ (.A(_07538_),
    .B(_07557_),
    .Y(_07558_));
 OAI21x1_ASAP7_75t_R _30031_ (.A1(_07352_),
    .A2(_07525_),
    .B(_07558_),
    .Y(_00155_));
 OAI21x1_ASAP7_75t_R _30032_ (.A1(net5337),
    .A2(net5333),
    .B(net6007),
    .Y(_07559_));
 NOR2x1_ASAP7_75t_R _30033_ (.A(net5335),
    .B(_07559_),
    .Y(_07560_));
 NAND2x1_ASAP7_75t_R _30034_ (.A(net5997),
    .B(_07430_),
    .Y(_07561_));
 NOR2x1_ASAP7_75t_R _30035_ (.A(_07560_),
    .B(_07561_),
    .Y(_07562_));
 AND2x2_ASAP7_75t_R _30036_ (.A(net5324),
    .B(_07315_),
    .Y(_07563_));
 OAI21x1_ASAP7_75t_R _30037_ (.A1(_07563_),
    .A2(_07324_),
    .B(net5993),
    .Y(_07564_));
 NOR2x1_ASAP7_75t_R _30038_ (.A(_07562_),
    .B(_07564_),
    .Y(_07565_));
 NAND2x1p5_ASAP7_75t_R _30039_ (.A(net6007),
    .B(net4992),
    .Y(_07566_));
 NAND2x1_ASAP7_75t_R _30040_ (.A(net4724),
    .B(_07455_),
    .Y(_07567_));
 NOR2x1_ASAP7_75t_R _30041_ (.A(_07507_),
    .B(_07567_),
    .Y(_07568_));
 OAI21x1_ASAP7_75t_R _30042_ (.A1(net4726),
    .A2(_07355_),
    .B(net5991),
    .Y(_07569_));
 OAI21x1_ASAP7_75t_R _30043_ (.A1(_07569_),
    .A2(_07305_),
    .B(net5987),
    .Y(_07570_));
 OAI21x1_ASAP7_75t_R _30044_ (.A1(_07568_),
    .A2(_07570_),
    .B(net5985),
    .Y(_07571_));
 OAI21x1_ASAP7_75t_R _30045_ (.A1(_07565_),
    .A2(_07571_),
    .B(net5573),
    .Y(_07572_));
 INVx1_ASAP7_75t_R _30046_ (.A(_07387_),
    .Y(_07573_));
 AO21x1_ASAP7_75t_R _30047_ (.A1(_07573_),
    .A2(_07494_),
    .B(net5986),
    .Y(_07574_));
 NAND2x1_ASAP7_75t_R _30048_ (.A(_07266_),
    .B(_07493_),
    .Y(_07575_));
 INVx1_ASAP7_75t_R _30049_ (.A(_07378_),
    .Y(_07576_));
 AO21x1_ASAP7_75t_R _30050_ (.A1(_07576_),
    .A2(_07200_),
    .B(net6008),
    .Y(_07577_));
 AOI21x1_ASAP7_75t_R _30051_ (.A1(_07575_),
    .A2(_07577_),
    .B(net5988),
    .Y(_07578_));
 AOI21x1_ASAP7_75t_R _30052_ (.A1(_07385_),
    .A2(_07393_),
    .B(_07346_),
    .Y(_07579_));
 AOI21x1_ASAP7_75t_R _30053_ (.A1(net6009),
    .A2(_07499_),
    .B(net5077),
    .Y(_07580_));
 AOI21x1_ASAP7_75t_R _30054_ (.A1(net5996),
    .A2(_07580_),
    .B(net5992),
    .Y(_07581_));
 OAI21x1_ASAP7_75t_R _30055_ (.A1(net5995),
    .A2(_07579_),
    .B(_07581_),
    .Y(_07582_));
 OAI21x1_ASAP7_75t_R _30056_ (.A1(_07574_),
    .A2(_07578_),
    .B(_07582_),
    .Y(_07583_));
 NOR2x1_ASAP7_75t_R _30057_ (.A(net5985),
    .B(_07583_),
    .Y(_07584_));
 OAI21x1_ASAP7_75t_R _30058_ (.A1(_01394_),
    .A2(net6005),
    .B(net4724),
    .Y(_07585_));
 AO21x1_ASAP7_75t_R _30059_ (.A1(_07585_),
    .A2(net5989),
    .B(net5993),
    .Y(_07586_));
 NAND2x1_ASAP7_75t_R _30060_ (.A(_07200_),
    .B(_07304_),
    .Y(_07587_));
 INVx1_ASAP7_75t_R _30061_ (.A(_07587_),
    .Y(_07588_));
 OAI21x1_ASAP7_75t_R _30062_ (.A1(net6005),
    .A2(_07321_),
    .B(net5997),
    .Y(_07589_));
 NOR2x1_ASAP7_75t_R _30063_ (.A(_07588_),
    .B(_07589_),
    .Y(_07590_));
 OAI21x1_ASAP7_75t_R _30064_ (.A1(_07586_),
    .A2(_07590_),
    .B(net5985),
    .Y(_07591_));
 NOR2x1_ASAP7_75t_R _30065_ (.A(_07289_),
    .B(_07290_),
    .Y(_07592_));
 NAND2x1_ASAP7_75t_R _30066_ (.A(net5989),
    .B(_07338_),
    .Y(_07593_));
 OAI21x1_ASAP7_75t_R _30067_ (.A1(_07592_),
    .A2(_07593_),
    .B(net5993),
    .Y(_07594_));
 AO21x1_ASAP7_75t_R _30068_ (.A1(net5586),
    .A2(net5583),
    .B(net6004),
    .Y(_07595_));
 OAI21x1_ASAP7_75t_R _30069_ (.A1(net5335),
    .A2(_07595_),
    .B(net5997),
    .Y(_07596_));
 AOI21x1_ASAP7_75t_R _30070_ (.A1(net4818),
    .A2(_07540_),
    .B(_07596_),
    .Y(_07597_));
 NOR2x1_ASAP7_75t_R _30071_ (.A(_07594_),
    .B(_07597_),
    .Y(_07598_));
 OAI21x1_ASAP7_75t_R _30072_ (.A1(_07591_),
    .A2(_07598_),
    .B(net5984),
    .Y(_07599_));
 AO21x1_ASAP7_75t_R _30073_ (.A1(net5579),
    .A2(net5270),
    .B(net6007),
    .Y(_07600_));
 OAI21x1_ASAP7_75t_R _30074_ (.A1(net4992),
    .A2(_07600_),
    .B(net5989),
    .Y(_07601_));
 NOR2x1_ASAP7_75t_R _30075_ (.A(_07601_),
    .B(_07188_),
    .Y(_07602_));
 AO21x1_ASAP7_75t_R _30076_ (.A1(net4815),
    .A2(net6003),
    .B(net5991),
    .Y(_07603_));
 OAI21x1_ASAP7_75t_R _30077_ (.A1(_07603_),
    .A2(_07354_),
    .B(net5987),
    .Y(_07604_));
 OAI21x1_ASAP7_75t_R _30078_ (.A1(_07602_),
    .A2(_07604_),
    .B(net5574),
    .Y(_07605_));
 OA21x2_ASAP7_75t_R _30079_ (.A1(_07230_),
    .A2(net5335),
    .B(net5994),
    .Y(_07606_));
 AO21x1_ASAP7_75t_R _30080_ (.A1(net5078),
    .A2(net4819),
    .B(net6006),
    .Y(_07607_));
 AO21x1_ASAP7_75t_R _30081_ (.A1(net5581),
    .A2(net6006),
    .B(net5996),
    .Y(_07608_));
 AOI21x1_ASAP7_75t_R _30082_ (.A1(_07288_),
    .A2(net4605),
    .B(_07608_),
    .Y(_07609_));
 AOI211x1_ASAP7_75t_R _30083_ (.A1(_07606_),
    .A2(_07607_),
    .B(_07609_),
    .C(net5987),
    .Y(_07610_));
 NOR2x1_ASAP7_75t_R _30084_ (.A(_07605_),
    .B(_07610_),
    .Y(_07611_));
 OAI22x1_ASAP7_75t_R _30085_ (.A1(_07572_),
    .A2(_07584_),
    .B1(_07599_),
    .B2(_07611_),
    .Y(_00156_));
 INVx1_ASAP7_75t_R _30086_ (.A(_07347_),
    .Y(_07612_));
 AOI221x1_ASAP7_75t_R _30087_ (.A1(net4605),
    .A2(_07439_),
    .B1(net4534),
    .B2(_07612_),
    .C(net5988),
    .Y(_07613_));
 NOR2x1_ASAP7_75t_R _30088_ (.A(net6009),
    .B(net5336),
    .Y(_07614_));
 NOR2x1_ASAP7_75t_R _30089_ (.A(net5326),
    .B(_07614_),
    .Y(_07615_));
 OA21x2_ASAP7_75t_R _30090_ (.A1(net4820),
    .A2(net6002),
    .B(net5988),
    .Y(_07616_));
 AO21x1_ASAP7_75t_R _30091_ (.A1(_07615_),
    .A2(_07616_),
    .B(_07234_),
    .Y(_07617_));
 OA21x2_ASAP7_75t_R _30092_ (.A1(_07330_),
    .A2(_07544_),
    .B(_07234_),
    .Y(_07618_));
 AND2x2_ASAP7_75t_R _30093_ (.A(_07475_),
    .B(net5988),
    .Y(_07619_));
 OAI21x1_ASAP7_75t_R _30094_ (.A1(_07232_),
    .A2(_07615_),
    .B(_07619_),
    .Y(_07620_));
 AOI21x1_ASAP7_75t_R _30095_ (.A1(_07618_),
    .A2(_07620_),
    .B(net5574),
    .Y(_07621_));
 OAI21x1_ASAP7_75t_R _30096_ (.A1(_07613_),
    .A2(_07617_),
    .B(_07621_),
    .Y(_07622_));
 AOI21x1_ASAP7_75t_R _30097_ (.A1(net5331),
    .A2(net4812),
    .B(net5991),
    .Y(_07623_));
 OAI21x1_ASAP7_75t_R _30098_ (.A1(net4450),
    .A2(_07232_),
    .B(_07623_),
    .Y(_07624_));
 OA21x2_ASAP7_75t_R _30099_ (.A1(net5583),
    .A2(net6001),
    .B(net5989),
    .Y(_07625_));
 NAND2x1_ASAP7_75t_R _30100_ (.A(_07286_),
    .B(_07288_),
    .Y(_07626_));
 AOI21x1_ASAP7_75t_R _30101_ (.A1(_07625_),
    .A2(_07626_),
    .B(net5993),
    .Y(_07627_));
 AOI21x1_ASAP7_75t_R _30102_ (.A1(_07624_),
    .A2(_07627_),
    .B(net5985),
    .Y(_07628_));
 AO21x1_ASAP7_75t_R _30103_ (.A1(_07540_),
    .A2(net4814),
    .B(net6007),
    .Y(_07629_));
 OAI21x1_ASAP7_75t_R _30104_ (.A1(net5334),
    .A2(_07187_),
    .B(_07629_),
    .Y(_07630_));
 OA21x2_ASAP7_75t_R _30105_ (.A1(_07262_),
    .A2(net6002),
    .B(net5996),
    .Y(_07631_));
 OAI21x1_ASAP7_75t_R _30106_ (.A1(net5326),
    .A2(_07614_),
    .B(_07214_),
    .Y(_07632_));
 AOI21x1_ASAP7_75t_R _30107_ (.A1(_07631_),
    .A2(_07632_),
    .B(_07234_),
    .Y(_07633_));
 OAI21x1_ASAP7_75t_R _30108_ (.A1(net5994),
    .A2(_07630_),
    .B(_07633_),
    .Y(_07634_));
 AOI21x1_ASAP7_75t_R _30109_ (.A1(_07628_),
    .A2(_07634_),
    .B(_07352_),
    .Y(_07635_));
 NAND2x1_ASAP7_75t_R _30110_ (.A(_07622_),
    .B(_07635_),
    .Y(_07636_));
 NAND2x1_ASAP7_75t_R _30111_ (.A(_07194_),
    .B(_07449_),
    .Y(_07637_));
 NOR2x1_ASAP7_75t_R _30112_ (.A(_07279_),
    .B(_07372_),
    .Y(_07638_));
 OAI21x1_ASAP7_75t_R _30113_ (.A1(_07637_),
    .A2(_07638_),
    .B(net5989),
    .Y(_07639_));
 AO21x1_ASAP7_75t_R _30114_ (.A1(net5575),
    .A2(net6004),
    .B(_07194_),
    .Y(_07640_));
 NOR2x1_ASAP7_75t_R _30115_ (.A(net5335),
    .B(_07595_),
    .Y(_07641_));
 NOR2x1_ASAP7_75t_R _30116_ (.A(_07640_),
    .B(_07641_),
    .Y(_07642_));
 OAI21x1_ASAP7_75t_R _30117_ (.A1(_07639_),
    .A2(_07642_),
    .B(net5985),
    .Y(_07643_));
 AND2x2_ASAP7_75t_R _30118_ (.A(_07358_),
    .B(net6003),
    .Y(_07644_));
 NAND2x1_ASAP7_75t_R _30119_ (.A(_07194_),
    .B(_07566_),
    .Y(_07645_));
 AO21x1_ASAP7_75t_R _30120_ (.A1(_07644_),
    .A2(net5333),
    .B(_07645_),
    .Y(_07646_));
 NOR2x1_ASAP7_75t_R _30121_ (.A(_07378_),
    .B(_07227_),
    .Y(_07647_));
 NAND2x1_ASAP7_75t_R _30122_ (.A(net6008),
    .B(_07262_),
    .Y(_07648_));
 NOR2x1_ASAP7_75t_R _30123_ (.A(_07648_),
    .B(_07383_),
    .Y(_07649_));
 OAI21x1_ASAP7_75t_R _30124_ (.A1(_07647_),
    .A2(_07649_),
    .B(net5986),
    .Y(_07650_));
 AOI21x1_ASAP7_75t_R _30125_ (.A1(_07646_),
    .A2(_07650_),
    .B(net5990),
    .Y(_07651_));
 NOR2x1_ASAP7_75t_R _30126_ (.A(_07643_),
    .B(_07651_),
    .Y(_07652_));
 AO21x1_ASAP7_75t_R _30127_ (.A1(_07296_),
    .A2(net5269),
    .B(net5999),
    .Y(_07653_));
 OAI21x1_ASAP7_75t_R _30128_ (.A1(net5582),
    .A2(net5328),
    .B(net4811),
    .Y(_07654_));
 AOI21x1_ASAP7_75t_R _30129_ (.A1(_07653_),
    .A2(_07654_),
    .B(net5989),
    .Y(_07655_));
 OAI21x1_ASAP7_75t_R _30130_ (.A1(net5077),
    .A2(net5335),
    .B(net5999),
    .Y(_07656_));
 AO21x1_ASAP7_75t_R _30131_ (.A1(_07423_),
    .A2(_07429_),
    .B(net5999),
    .Y(_07657_));
 AOI21x1_ASAP7_75t_R _30132_ (.A1(_07656_),
    .A2(_07657_),
    .B(net5997),
    .Y(_07658_));
 OAI21x1_ASAP7_75t_R _30133_ (.A1(_07655_),
    .A2(_07658_),
    .B(net5987),
    .Y(_07659_));
 NAND2x1_ASAP7_75t_R _30134_ (.A(_07404_),
    .B(net5328),
    .Y(_07660_));
 AOI21x1_ASAP7_75t_R _30135_ (.A1(_07600_),
    .A2(_07660_),
    .B(net5989),
    .Y(_07661_));
 NAND2x1_ASAP7_75t_R _30136_ (.A(net5581),
    .B(net5583),
    .Y(_07662_));
 AO21x1_ASAP7_75t_R _30137_ (.A1(_07662_),
    .A2(net4817),
    .B(net6003),
    .Y(_07663_));
 AOI21x1_ASAP7_75t_R _30138_ (.A1(_07274_),
    .A2(_07663_),
    .B(net5996),
    .Y(_07664_));
 OAI21x1_ASAP7_75t_R _30139_ (.A1(_07661_),
    .A2(_07664_),
    .B(net5993),
    .Y(_07665_));
 AOI21x1_ASAP7_75t_R _30140_ (.A1(_07659_),
    .A2(_07665_),
    .B(net5985),
    .Y(_07666_));
 OAI21x1_ASAP7_75t_R _30141_ (.A1(_07652_),
    .A2(_07666_),
    .B(net5573),
    .Y(_07667_));
 NAND2x1_ASAP7_75t_R _30142_ (.A(_07636_),
    .B(_07667_),
    .Y(_00157_));
 AOI21x1_ASAP7_75t_R _30143_ (.A1(_07301_),
    .A2(_07587_),
    .B(net5989),
    .Y(_07668_));
 OAI21x1_ASAP7_75t_R _30144_ (.A1(_07668_),
    .A2(_07436_),
    .B(net5993),
    .Y(_07669_));
 OA21x2_ASAP7_75t_R _30145_ (.A1(_07372_),
    .A2(net4813),
    .B(_07400_),
    .Y(_07670_));
 AND2x2_ASAP7_75t_R _30146_ (.A(net6004),
    .B(_01398_),
    .Y(_07671_));
 AOI21x1_ASAP7_75t_R _30147_ (.A1(_07200_),
    .A2(net4811),
    .B(_07671_),
    .Y(_07672_));
 AOI21x1_ASAP7_75t_R _30148_ (.A1(net5989),
    .A2(_07672_),
    .B(_07194_),
    .Y(_07673_));
 OAI21x1_ASAP7_75t_R _30149_ (.A1(net5989),
    .A2(_07670_),
    .B(_07673_),
    .Y(_07674_));
 NAND2x1_ASAP7_75t_R _30150_ (.A(_07674_),
    .B(_07669_),
    .Y(_07675_));
 OAI21x1_ASAP7_75t_R _30151_ (.A1(net5574),
    .A2(_07675_),
    .B(net5984),
    .Y(_07676_));
 OA21x2_ASAP7_75t_R _30152_ (.A1(net5586),
    .A2(net6005),
    .B(_07541_),
    .Y(_07677_));
 AOI21x1_ASAP7_75t_R _30153_ (.A1(net5989),
    .A2(_07677_),
    .B(net5993),
    .Y(_07678_));
 AOI21x1_ASAP7_75t_R _30154_ (.A1(net6005),
    .A2(_07541_),
    .B(net5989),
    .Y(_07679_));
 OAI21x1_ASAP7_75t_R _30155_ (.A1(net5329),
    .A2(net4482),
    .B(_07679_),
    .Y(_07680_));
 NAND2x1_ASAP7_75t_R _30156_ (.A(net4816),
    .B(_07662_),
    .Y(_07681_));
 NOR2x1_ASAP7_75t_R _30157_ (.A(net6006),
    .B(_07267_),
    .Y(_07682_));
 AOI211x1_ASAP7_75t_R _30158_ (.A1(_07681_),
    .A2(net6006),
    .B(_07682_),
    .C(net5996),
    .Y(_07683_));
 NAND2x1_ASAP7_75t_R _30159_ (.A(net5996),
    .B(_07393_),
    .Y(_07684_));
 OAI21x1_ASAP7_75t_R _30160_ (.A1(_07684_),
    .A2(_07222_),
    .B(net5992),
    .Y(_07685_));
 NOR2x1_ASAP7_75t_R _30161_ (.A(_07683_),
    .B(_07685_),
    .Y(_07686_));
 AOI211x1_ASAP7_75t_R _30162_ (.A1(_07678_),
    .A2(_07680_),
    .B(_07686_),
    .C(net5985),
    .Y(_07687_));
 NAND2x1_ASAP7_75t_R _30163_ (.A(_07404_),
    .B(_07576_),
    .Y(_07688_));
 OA21x2_ASAP7_75t_R _30164_ (.A1(_07296_),
    .A2(net5999),
    .B(net5989),
    .Y(_07689_));
 NAND2x1_ASAP7_75t_R _30165_ (.A(_07205_),
    .B(_07458_),
    .Y(_07690_));
 AND3x1_ASAP7_75t_R _30166_ (.A(_07688_),
    .B(_07689_),
    .C(_07690_),
    .Y(_07691_));
 NOR2x1_ASAP7_75t_R _30167_ (.A(_07219_),
    .B(_07548_),
    .Y(_07692_));
 OAI21x1_ASAP7_75t_R _30168_ (.A1(net5073),
    .A2(_07508_),
    .B(_07506_),
    .Y(_07693_));
 OAI21x1_ASAP7_75t_R _30169_ (.A1(_07692_),
    .A2(_07693_),
    .B(_07194_),
    .Y(_07694_));
 NAND2x1_ASAP7_75t_R _30170_ (.A(net5328),
    .B(_07463_),
    .Y(_07695_));
 AO21x1_ASAP7_75t_R _30171_ (.A1(_01397_),
    .A2(_01401_),
    .B(net6004),
    .Y(_07696_));
 NAND3x1_ASAP7_75t_R _30172_ (.A(_07695_),
    .B(net5989),
    .C(_07696_),
    .Y(_07697_));
 OAI21x1_ASAP7_75t_R _30173_ (.A1(net6009),
    .A2(_07412_),
    .B(_07441_),
    .Y(_07698_));
 AOI21x1_ASAP7_75t_R _30174_ (.A1(_07506_),
    .A2(_07698_),
    .B(_07194_),
    .Y(_07699_));
 AOI21x1_ASAP7_75t_R _30175_ (.A1(_07697_),
    .A2(_07699_),
    .B(net5985),
    .Y(_07700_));
 OAI21x1_ASAP7_75t_R _30176_ (.A1(_07691_),
    .A2(_07694_),
    .B(_07700_),
    .Y(_07701_));
 AOI21x1_ASAP7_75t_R _30177_ (.A1(_07500_),
    .A2(_07311_),
    .B(_07179_),
    .Y(_07702_));
 OAI21x1_ASAP7_75t_R _30178_ (.A1(_07289_),
    .A2(_07559_),
    .B(_07702_),
    .Y(_07703_));
 OAI21x1_ASAP7_75t_R _30179_ (.A1(net5575),
    .A2(_07219_),
    .B(net6007),
    .Y(_07704_));
 OA21x2_ASAP7_75t_R _30180_ (.A1(_07262_),
    .A2(net6009),
    .B(_07179_),
    .Y(_07705_));
 AOI21x1_ASAP7_75t_R _30181_ (.A1(_07704_),
    .A2(_07705_),
    .B(net5986),
    .Y(_07706_));
 AOI21x1_ASAP7_75t_R _30182_ (.A1(_07703_),
    .A2(_07706_),
    .B(net5574),
    .Y(_07707_));
 INVx1_ASAP7_75t_R _30183_ (.A(_07515_),
    .Y(_07708_));
 AOI21x1_ASAP7_75t_R _30184_ (.A1(_07469_),
    .A2(_07202_),
    .B(_07708_),
    .Y(_07709_));
 AOI21x1_ASAP7_75t_R _30185_ (.A1(_07358_),
    .A2(_07439_),
    .B(net5994),
    .Y(_07710_));
 INVx1_ASAP7_75t_R _30186_ (.A(net5333),
    .Y(_07711_));
 OAI21x1_ASAP7_75t_R _30187_ (.A1(_07217_),
    .A2(_07711_),
    .B(net6009),
    .Y(_07712_));
 AOI21x1_ASAP7_75t_R _30188_ (.A1(_07710_),
    .A2(_07712_),
    .B(net5992),
    .Y(_07713_));
 OAI21x1_ASAP7_75t_R _30189_ (.A1(net5990),
    .A2(_07709_),
    .B(_07713_),
    .Y(_07714_));
 AOI21x1_ASAP7_75t_R _30190_ (.A1(_07707_),
    .A2(_07714_),
    .B(net5984),
    .Y(_07715_));
 NAND2x1_ASAP7_75t_R _30191_ (.A(_07701_),
    .B(_07715_),
    .Y(_07716_));
 OAI21x1_ASAP7_75t_R _30192_ (.A1(_07687_),
    .A2(_07676_),
    .B(_07716_),
    .Y(_00158_));
 AND3x1_ASAP7_75t_R _30193_ (.A(_07460_),
    .B(_07267_),
    .C(net6006),
    .Y(_07717_));
 AO21x1_ASAP7_75t_R _30194_ (.A1(_07226_),
    .A2(net5331),
    .B(net5988),
    .Y(_07718_));
 NAND2x1_ASAP7_75t_R _30195_ (.A(net6002),
    .B(net4726),
    .Y(_07719_));
 OAI21x1_ASAP7_75t_R _30196_ (.A1(_01401_),
    .A2(net5998),
    .B(net5988),
    .Y(_07720_));
 NOR2x1_ASAP7_75t_R _30197_ (.A(_07720_),
    .B(_07451_),
    .Y(_07721_));
 AOI21x1_ASAP7_75t_R _30198_ (.A1(_07719_),
    .A2(_07721_),
    .B(_07234_),
    .Y(_07722_));
 OA21x2_ASAP7_75t_R _30199_ (.A1(_07717_),
    .A2(_07718_),
    .B(_07722_),
    .Y(_07723_));
 AO21x1_ASAP7_75t_R _30200_ (.A1(_07540_),
    .A2(net5586),
    .B(net6005),
    .Y(_07724_));
 NAND2x1_ASAP7_75t_R _30201_ (.A(_07724_),
    .B(_07606_),
    .Y(_07725_));
 AOI21x1_ASAP7_75t_R _30202_ (.A1(_01394_),
    .A2(net6005),
    .B(net5997),
    .Y(_07726_));
 AOI21x1_ASAP7_75t_R _30203_ (.A1(_07726_),
    .A2(_07318_),
    .B(net5993),
    .Y(_07727_));
 AO21x1_ASAP7_75t_R _30204_ (.A1(_07725_),
    .A2(_07727_),
    .B(net5574),
    .Y(_07728_));
 NOR2x1_ASAP7_75t_R _30205_ (.A(_07723_),
    .B(_07728_),
    .Y(_07729_));
 OA21x2_ASAP7_75t_R _30206_ (.A1(net5575),
    .A2(net5584),
    .B(net5581),
    .Y(_07730_));
 OAI21x1_ASAP7_75t_R _30207_ (.A1(_07412_),
    .A2(_07730_),
    .B(net6002),
    .Y(_07731_));
 OA21x2_ASAP7_75t_R _30208_ (.A1(_07347_),
    .A2(_07256_),
    .B(net5988),
    .Y(_07732_));
 AOI21x1_ASAP7_75t_R _30209_ (.A1(_07731_),
    .A2(_07732_),
    .B(net5992),
    .Y(_07733_));
 AO21x1_ASAP7_75t_R _30210_ (.A1(_07576_),
    .A2(_07342_),
    .B(net5988),
    .Y(_07734_));
 OR2x2_ASAP7_75t_R _30211_ (.A(_07501_),
    .B(_07734_),
    .Y(_07735_));
 AND2x2_ASAP7_75t_R _30212_ (.A(_07733_),
    .B(_07735_),
    .Y(_07736_));
 INVx1_ASAP7_75t_R _30213_ (.A(_07393_),
    .Y(_07737_));
 OAI21x1_ASAP7_75t_R _30214_ (.A1(_07644_),
    .A2(_07737_),
    .B(_07315_),
    .Y(_07738_));
 NAND2x1_ASAP7_75t_R _30215_ (.A(net5990),
    .B(_07738_),
    .Y(_07739_));
 OA21x2_ASAP7_75t_R _30216_ (.A1(net5269),
    .A2(net6004),
    .B(net5997),
    .Y(_07740_));
 AOI21x1_ASAP7_75t_R _30217_ (.A1(_07740_),
    .A2(_07695_),
    .B(_07234_),
    .Y(_07741_));
 AO21x1_ASAP7_75t_R _30218_ (.A1(_07739_),
    .A2(_07741_),
    .B(net5985),
    .Y(_07742_));
 OAI21x1_ASAP7_75t_R _30219_ (.A1(_07736_),
    .A2(_07742_),
    .B(_07352_),
    .Y(_07743_));
 NOR2x1_ASAP7_75t_R _30220_ (.A(_07346_),
    .B(_07393_),
    .Y(_07744_));
 OA21x2_ASAP7_75t_R _30221_ (.A1(_07744_),
    .A2(_07614_),
    .B(net5995),
    .Y(_07745_));
 OAI21x1_ASAP7_75t_R _30222_ (.A1(_07711_),
    .A2(_07730_),
    .B(net6002),
    .Y(_07746_));
 AO21x1_ASAP7_75t_R _30223_ (.A1(_07746_),
    .A2(_07494_),
    .B(net5992),
    .Y(_07747_));
 OAI21x1_ASAP7_75t_R _30224_ (.A1(net5584),
    .A2(net5330),
    .B(_07439_),
    .Y(_07748_));
 AOI21x1_ASAP7_75t_R _30225_ (.A1(_07559_),
    .A2(_07748_),
    .B(net5990),
    .Y(_07749_));
 OA21x2_ASAP7_75t_R _30226_ (.A1(net4727),
    .A2(net6008),
    .B(net5988),
    .Y(_07750_));
 OA21x2_ASAP7_75t_R _30227_ (.A1(net6002),
    .A2(_07383_),
    .B(_07750_),
    .Y(_07751_));
 OAI21x1_ASAP7_75t_R _30228_ (.A1(_07749_),
    .A2(_07751_),
    .B(net5992),
    .Y(_07752_));
 OAI21x1_ASAP7_75t_R _30229_ (.A1(_07745_),
    .A2(_07747_),
    .B(_07752_),
    .Y(_07753_));
 AOI21x1_ASAP7_75t_R _30230_ (.A1(net6000),
    .A2(net4606),
    .B(_07194_),
    .Y(_07754_));
 AOI21x1_ASAP7_75t_R _30231_ (.A1(_07587_),
    .A2(_07754_),
    .B(net5997),
    .Y(_07755_));
 AOI21x1_ASAP7_75t_R _30232_ (.A1(net5325),
    .A2(net5324),
    .B(_07234_),
    .Y(_07756_));
 NAND2x1_ASAP7_75t_R _30233_ (.A(_07690_),
    .B(_07756_),
    .Y(_07757_));
 AOI21x1_ASAP7_75t_R _30234_ (.A1(_07755_),
    .A2(_07757_),
    .B(net5985),
    .Y(_07758_));
 OA21x2_ASAP7_75t_R _30235_ (.A1(_07730_),
    .A2(_07412_),
    .B(net6009),
    .Y(_07759_));
 AO21x1_ASAP7_75t_R _30236_ (.A1(net5575),
    .A2(net5580),
    .B(net5337),
    .Y(_07760_));
 AO21x1_ASAP7_75t_R _30237_ (.A1(_07760_),
    .A2(_07171_),
    .B(_07194_),
    .Y(_07761_));
 AOI21x1_ASAP7_75t_R _30238_ (.A1(_07396_),
    .A2(_07521_),
    .B(net5990),
    .Y(_07762_));
 OAI21x1_ASAP7_75t_R _30239_ (.A1(_07759_),
    .A2(_07761_),
    .B(_07762_),
    .Y(_07763_));
 AOI21x1_ASAP7_75t_R _30240_ (.A1(_07758_),
    .A2(_07763_),
    .B(_07352_),
    .Y(_07764_));
 OAI21x1_ASAP7_75t_R _30241_ (.A1(net5574),
    .A2(_07753_),
    .B(_07764_),
    .Y(_07765_));
 OAI21x1_ASAP7_75t_R _30242_ (.A1(_07729_),
    .A2(_07743_),
    .B(_07765_),
    .Y(_00159_));
 INVx1_ASAP7_75t_R _30243_ (.A(_00488_),
    .Y(net387));
 INVx1_ASAP7_75t_R _30244_ (.A(_00573_),
    .Y(net259));
 INVx1_ASAP7_75t_R _30245_ (.A(_00702_),
    .Y(net260));
 INVx1_ASAP7_75t_R _30246_ (.A(_00703_),
    .Y(net261));
 INVx1_ASAP7_75t_R _30247_ (.A(_00704_),
    .Y(net262));
 INVx1_ASAP7_75t_R _30248_ (.A(_00705_),
    .Y(net263));
 INVx1_ASAP7_75t_R _30249_ (.A(_00706_),
    .Y(net264));
 INVx1_ASAP7_75t_R _30250_ (.A(_00707_),
    .Y(net265));
 INVx1_ASAP7_75t_R _30251_ (.A(_00708_),
    .Y(net266));
 INVx1_ASAP7_75t_R _30252_ (.A(_00709_),
    .Y(net267));
 INVx1_ASAP7_75t_R _30253_ (.A(_00710_),
    .Y(net268));
 INVx1_ASAP7_75t_R _30254_ (.A(_00711_),
    .Y(net269));
 INVx1_ASAP7_75t_R _30255_ (.A(_00712_),
    .Y(net270));
 INVx1_ASAP7_75t_R _30256_ (.A(_00713_),
    .Y(net271));
 INVx1_ASAP7_75t_R _30257_ (.A(_00714_),
    .Y(net272));
 INVx1_ASAP7_75t_R _30258_ (.A(_00715_),
    .Y(net273));
 INVx1_ASAP7_75t_R _30259_ (.A(_00716_),
    .Y(net274));
 INVx1_ASAP7_75t_R _30260_ (.A(_00717_),
    .Y(net275));
 INVx1_ASAP7_75t_R _30261_ (.A(_00718_),
    .Y(net276));
 INVx1_ASAP7_75t_R _30262_ (.A(_00719_),
    .Y(net277));
 INVx1_ASAP7_75t_R _30263_ (.A(_00720_),
    .Y(net278));
 INVx1_ASAP7_75t_R _30264_ (.A(_00721_),
    .Y(net279));
 INVx1_ASAP7_75t_R _30265_ (.A(_00722_),
    .Y(net280));
 INVx1_ASAP7_75t_R _30266_ (.A(_00723_),
    .Y(net281));
 INVx1_ASAP7_75t_R _30267_ (.A(_00724_),
    .Y(net282));
 INVx1_ASAP7_75t_R _30268_ (.A(_00725_),
    .Y(net283));
 INVx1_ASAP7_75t_R _30269_ (.A(_00726_),
    .Y(net284));
 INVx1_ASAP7_75t_R _30270_ (.A(_00727_),
    .Y(net285));
 INVx1_ASAP7_75t_R _30271_ (.A(_00728_),
    .Y(net286));
 INVx1_ASAP7_75t_R _30272_ (.A(_00729_),
    .Y(net287));
 INVx1_ASAP7_75t_R _30273_ (.A(_00730_),
    .Y(net288));
 INVx1_ASAP7_75t_R _30274_ (.A(_00731_),
    .Y(net289));
 INVx1_ASAP7_75t_R _30275_ (.A(_00732_),
    .Y(net290));
 INVx1_ASAP7_75t_R _30276_ (.A(_00733_),
    .Y(net291));
 INVx1_ASAP7_75t_R _30277_ (.A(_00734_),
    .Y(net292));
 INVx1_ASAP7_75t_R _30278_ (.A(_00735_),
    .Y(net293));
 INVx1_ASAP7_75t_R _30279_ (.A(_00736_),
    .Y(net294));
 INVx1_ASAP7_75t_R _30280_ (.A(_00737_),
    .Y(net295));
 INVx1_ASAP7_75t_R _30281_ (.A(_00738_),
    .Y(net296));
 INVx1_ASAP7_75t_R _30282_ (.A(_00739_),
    .Y(net297));
 INVx1_ASAP7_75t_R _30283_ (.A(_00740_),
    .Y(net298));
 INVx1_ASAP7_75t_R _30284_ (.A(_00741_),
    .Y(net299));
 INVx1_ASAP7_75t_R _30285_ (.A(_00742_),
    .Y(net300));
 INVx1_ASAP7_75t_R _30286_ (.A(_00743_),
    .Y(net301));
 INVx1_ASAP7_75t_R _30287_ (.A(_00744_),
    .Y(net302));
 INVx1_ASAP7_75t_R _30288_ (.A(_00745_),
    .Y(net303));
 INVx1_ASAP7_75t_R _30289_ (.A(_00746_),
    .Y(net304));
 INVx1_ASAP7_75t_R _30290_ (.A(_00747_),
    .Y(net305));
 INVx1_ASAP7_75t_R _30291_ (.A(_00748_),
    .Y(net306));
 INVx1_ASAP7_75t_R _30292_ (.A(_00749_),
    .Y(net307));
 INVx1_ASAP7_75t_R _30293_ (.A(_00750_),
    .Y(net308));
 INVx1_ASAP7_75t_R _30294_ (.A(_00751_),
    .Y(net309));
 INVx1_ASAP7_75t_R _30295_ (.A(_00752_),
    .Y(net310));
 INVx1_ASAP7_75t_R _30296_ (.A(_00753_),
    .Y(net311));
 INVx1_ASAP7_75t_R _30297_ (.A(_00754_),
    .Y(net312));
 INVx1_ASAP7_75t_R _30298_ (.A(_00755_),
    .Y(net313));
 INVx1_ASAP7_75t_R _30299_ (.A(_00756_),
    .Y(net314));
 INVx1_ASAP7_75t_R _30300_ (.A(_00757_),
    .Y(net315));
 INVx1_ASAP7_75t_R _30301_ (.A(_00758_),
    .Y(net316));
 INVx1_ASAP7_75t_R _30302_ (.A(_00759_),
    .Y(net317));
 INVx1_ASAP7_75t_R _30303_ (.A(_00760_),
    .Y(net318));
 INVx1_ASAP7_75t_R _30304_ (.A(_00761_),
    .Y(net319));
 INVx1_ASAP7_75t_R _30305_ (.A(_00762_),
    .Y(net320));
 INVx1_ASAP7_75t_R _30306_ (.A(_00763_),
    .Y(net321));
 INVx1_ASAP7_75t_R _30307_ (.A(_00764_),
    .Y(net322));
 INVx1_ASAP7_75t_R _30308_ (.A(_00765_),
    .Y(net323));
 INVx1_ASAP7_75t_R _30309_ (.A(_00766_),
    .Y(net324));
 INVx1_ASAP7_75t_R _30310_ (.A(_00767_),
    .Y(net325));
 INVx1_ASAP7_75t_R _30311_ (.A(_00768_),
    .Y(net326));
 INVx1_ASAP7_75t_R _30312_ (.A(_00769_),
    .Y(net327));
 INVx1_ASAP7_75t_R _30313_ (.A(_00770_),
    .Y(net328));
 INVx1_ASAP7_75t_R _30314_ (.A(_00771_),
    .Y(net329));
 INVx1_ASAP7_75t_R _30315_ (.A(_00772_),
    .Y(net330));
 INVx1_ASAP7_75t_R _30316_ (.A(_00773_),
    .Y(net331));
 INVx1_ASAP7_75t_R _30317_ (.A(_00774_),
    .Y(net332));
 INVx1_ASAP7_75t_R _30318_ (.A(_00775_),
    .Y(net333));
 INVx1_ASAP7_75t_R _30319_ (.A(_00776_),
    .Y(net334));
 INVx1_ASAP7_75t_R _30320_ (.A(_00777_),
    .Y(net335));
 INVx1_ASAP7_75t_R _30321_ (.A(_00778_),
    .Y(net336));
 INVx1_ASAP7_75t_R _30322_ (.A(_00779_),
    .Y(net337));
 INVx1_ASAP7_75t_R _30323_ (.A(_00780_),
    .Y(net338));
 INVx1_ASAP7_75t_R _30324_ (.A(_00781_),
    .Y(net339));
 INVx1_ASAP7_75t_R _30325_ (.A(_00782_),
    .Y(net340));
 INVx1_ASAP7_75t_R _30326_ (.A(_00783_),
    .Y(net341));
 INVx1_ASAP7_75t_R _30327_ (.A(_00784_),
    .Y(net342));
 INVx1_ASAP7_75t_R _30328_ (.A(_00785_),
    .Y(net343));
 INVx1_ASAP7_75t_R _30329_ (.A(_00786_),
    .Y(net344));
 INVx1_ASAP7_75t_R _30330_ (.A(_00787_),
    .Y(net345));
 INVx1_ASAP7_75t_R _30331_ (.A(_00788_),
    .Y(net346));
 INVx1_ASAP7_75t_R _30332_ (.A(_00789_),
    .Y(net347));
 INVx1_ASAP7_75t_R _30333_ (.A(_00790_),
    .Y(net348));
 INVx1_ASAP7_75t_R _30334_ (.A(_00791_),
    .Y(net349));
 INVx1_ASAP7_75t_R _30335_ (.A(_00792_),
    .Y(net350));
 INVx1_ASAP7_75t_R _30336_ (.A(_00793_),
    .Y(net351));
 INVx1_ASAP7_75t_R _30337_ (.A(_00794_),
    .Y(net352));
 INVx1_ASAP7_75t_R _30338_ (.A(_00795_),
    .Y(net353));
 INVx1_ASAP7_75t_R _30339_ (.A(_00796_),
    .Y(net354));
 INVx1_ASAP7_75t_R _30340_ (.A(_00797_),
    .Y(net355));
 INVx1_ASAP7_75t_R _30341_ (.A(_00798_),
    .Y(net356));
 INVx1_ASAP7_75t_R _30342_ (.A(_00799_),
    .Y(net357));
 INVx1_ASAP7_75t_R _30343_ (.A(_00800_),
    .Y(net358));
 INVx1_ASAP7_75t_R _30344_ (.A(_00801_),
    .Y(net359));
 INVx1_ASAP7_75t_R _30345_ (.A(_00802_),
    .Y(net360));
 INVx1_ASAP7_75t_R _30346_ (.A(_00803_),
    .Y(net361));
 INVx1_ASAP7_75t_R _30347_ (.A(_00804_),
    .Y(net362));
 INVx1_ASAP7_75t_R _30348_ (.A(_00805_),
    .Y(net363));
 INVx1_ASAP7_75t_R _30349_ (.A(_00806_),
    .Y(net364));
 INVx1_ASAP7_75t_R _30350_ (.A(_00807_),
    .Y(net365));
 INVx1_ASAP7_75t_R _30351_ (.A(_00808_),
    .Y(net366));
 INVx1_ASAP7_75t_R _30352_ (.A(_00809_),
    .Y(net367));
 INVx1_ASAP7_75t_R _30353_ (.A(_00810_),
    .Y(net368));
 INVx1_ASAP7_75t_R _30354_ (.A(_00811_),
    .Y(net369));
 INVx1_ASAP7_75t_R _30355_ (.A(_00812_),
    .Y(net370));
 INVx1_ASAP7_75t_R _30356_ (.A(_00813_),
    .Y(net371));
 INVx1_ASAP7_75t_R _30357_ (.A(_00814_),
    .Y(net372));
 INVx1_ASAP7_75t_R _30358_ (.A(_00815_),
    .Y(net373));
 INVx1_ASAP7_75t_R _30359_ (.A(_00816_),
    .Y(net374));
 INVx1_ASAP7_75t_R _30360_ (.A(_00817_),
    .Y(net375));
 INVx1_ASAP7_75t_R _30361_ (.A(_00818_),
    .Y(net376));
 INVx1_ASAP7_75t_R _30362_ (.A(_00819_),
    .Y(net377));
 INVx1_ASAP7_75t_R _30363_ (.A(_00820_),
    .Y(net378));
 INVx1_ASAP7_75t_R _30364_ (.A(_00821_),
    .Y(net379));
 INVx1_ASAP7_75t_R _30365_ (.A(_00822_),
    .Y(net380));
 INVx1_ASAP7_75t_R _30366_ (.A(_00823_),
    .Y(net381));
 INVx1_ASAP7_75t_R _30367_ (.A(_00824_),
    .Y(net382));
 INVx1_ASAP7_75t_R _30368_ (.A(_00825_),
    .Y(net383));
 INVx1_ASAP7_75t_R _30369_ (.A(_00826_),
    .Y(net384));
 INVx1_ASAP7_75t_R _30370_ (.A(_00827_),
    .Y(net385));
 INVx1_ASAP7_75t_R _30371_ (.A(_00828_),
    .Y(net386));
 NOR2x1_ASAP7_75t_R _30372_ (.A(net6684),
    .B(_00409_),
    .Y(_07766_));
 AO21x1_ASAP7_75t_R _30373_ (.A1(net6684),
    .A2(net131),
    .B(_07766_),
    .Y(_01409_));
 NOR2x1_ASAP7_75t_R _30374_ (.A(net6681),
    .B(_00568_),
    .Y(_07767_));
 AO21x1_ASAP7_75t_R _30375_ (.A1(net6681),
    .A2(net132),
    .B(_07767_),
    .Y(_01410_));
 NOR2x1_ASAP7_75t_R _30376_ (.A(net6681),
    .B(_00567_),
    .Y(_07768_));
 AO21x1_ASAP7_75t_R _30377_ (.A1(net6681),
    .A2(net133),
    .B(_07768_),
    .Y(_01411_));
 NOR2x1_ASAP7_75t_R _30378_ (.A(net6681),
    .B(_00566_),
    .Y(_07769_));
 AO21x1_ASAP7_75t_R _30379_ (.A1(net6681),
    .A2(net134),
    .B(_07769_),
    .Y(_01412_));
 NOR2x1_ASAP7_75t_R _30380_ (.A(net6680),
    .B(_00565_),
    .Y(_07770_));
 AO21x1_ASAP7_75t_R _30381_ (.A1(net6680),
    .A2(net135),
    .B(_07770_),
    .Y(_01413_));
 NOR2x1_ASAP7_75t_R _30382_ (.A(net6681),
    .B(_00469_),
    .Y(_07771_));
 AO21x1_ASAP7_75t_R _30383_ (.A1(net6681),
    .A2(net136),
    .B(_07771_),
    .Y(_01414_));
 NOR2x1_ASAP7_75t_R _30384_ (.A(net6682),
    .B(_00468_),
    .Y(_07772_));
 AO21x1_ASAP7_75t_R _30385_ (.A1(net6682),
    .A2(net137),
    .B(_07772_),
    .Y(_01415_));
 NOR2x1_ASAP7_75t_R _30387_ (.A(net6682),
    .B(_00470_),
    .Y(_07774_));
 AO21x1_ASAP7_75t_R _30388_ (.A1(net6682),
    .A2(net138),
    .B(_07774_),
    .Y(_01416_));
 NOR2x1_ASAP7_75t_R _30389_ (.A(net6681),
    .B(_00564_),
    .Y(_07775_));
 AO21x1_ASAP7_75t_R _30390_ (.A1(net6681),
    .A2(net139),
    .B(_07775_),
    .Y(_01417_));
 NOR2x1_ASAP7_75t_R _30392_ (.A(net6680),
    .B(_00563_),
    .Y(_07777_));
 AO21x1_ASAP7_75t_R _30393_ (.A1(net6680),
    .A2(net140),
    .B(_07777_),
    .Y(_01418_));
 NOR2x1_ASAP7_75t_R _30394_ (.A(net6680),
    .B(_00562_),
    .Y(_07778_));
 AO21x1_ASAP7_75t_R _30395_ (.A1(net6680),
    .A2(net141),
    .B(_07778_),
    .Y(_01419_));
 NOR2x1_ASAP7_75t_R _30396_ (.A(net6686),
    .B(_00479_),
    .Y(_07779_));
 AO21x1_ASAP7_75t_R _30397_ (.A1(net6686),
    .A2(net142),
    .B(_07779_),
    .Y(_01420_));
 NOR2x1_ASAP7_75t_R _30398_ (.A(net6680),
    .B(_00561_),
    .Y(_07780_));
 AO21x1_ASAP7_75t_R _30399_ (.A1(net6680),
    .A2(net143),
    .B(_07780_),
    .Y(_01421_));
 NOR2x1_ASAP7_75t_R _30400_ (.A(net6680),
    .B(_00560_),
    .Y(_07781_));
 AO21x1_ASAP7_75t_R _30401_ (.A1(net6680),
    .A2(net144),
    .B(_07781_),
    .Y(_01422_));
 NOR2x1_ASAP7_75t_R _30402_ (.A(net6684),
    .B(_00457_),
    .Y(_07782_));
 AO21x1_ASAP7_75t_R _30403_ (.A1(net6684),
    .A2(net145),
    .B(_07782_),
    .Y(_01423_));
 NOR2x1_ASAP7_75t_R _30404_ (.A(net6683),
    .B(_00456_),
    .Y(_07783_));
 AO21x1_ASAP7_75t_R _30405_ (.A1(net6683),
    .A2(net146),
    .B(_07783_),
    .Y(_01424_));
 NOR2x1_ASAP7_75t_R _30406_ (.A(net6684),
    .B(_00458_),
    .Y(_07784_));
 AO21x1_ASAP7_75t_R _30407_ (.A1(net6684),
    .A2(net147),
    .B(_07784_),
    .Y(_01425_));
 NOR2x1_ASAP7_75t_R _30409_ (.A(net6684),
    .B(_00559_),
    .Y(_07786_));
 AO21x1_ASAP7_75t_R _30410_ (.A1(net6684),
    .A2(net148),
    .B(_07786_),
    .Y(_01426_));
 NOR2x1_ASAP7_75t_R _30411_ (.A(net6682),
    .B(_00558_),
    .Y(_07787_));
 AO21x1_ASAP7_75t_R _30412_ (.A1(net6682),
    .A2(net149),
    .B(_07787_),
    .Y(_01427_));
 NOR2x1_ASAP7_75t_R _30415_ (.A(net6681),
    .B(_00557_),
    .Y(_07790_));
 AO21x1_ASAP7_75t_R _30416_ (.A1(net6681),
    .A2(net150),
    .B(_07790_),
    .Y(_01428_));
 NOR2x1_ASAP7_75t_R _30417_ (.A(net6681),
    .B(_00556_),
    .Y(_07791_));
 AO21x1_ASAP7_75t_R _30418_ (.A1(net6681),
    .A2(net151),
    .B(_07791_),
    .Y(_01429_));
 NOR2x1_ASAP7_75t_R _30419_ (.A(net6683),
    .B(_00555_),
    .Y(_07792_));
 AO21x1_ASAP7_75t_R _30420_ (.A1(net6683),
    .A2(net152),
    .B(_07792_),
    .Y(_01430_));
 NOR2x1_ASAP7_75t_R _30421_ (.A(net6689),
    .B(_00554_),
    .Y(_07793_));
 AO21x1_ASAP7_75t_R _30422_ (.A1(net6689),
    .A2(net153),
    .B(_07793_),
    .Y(_01431_));
 NOR2x1_ASAP7_75t_R _30423_ (.A(net6681),
    .B(_00445_),
    .Y(_07794_));
 AO21x1_ASAP7_75t_R _30424_ (.A1(net6681),
    .A2(net154),
    .B(_07794_),
    .Y(_01432_));
 NOR2x1_ASAP7_75t_R _30425_ (.A(net6681),
    .B(_00444_),
    .Y(_07795_));
 AO21x1_ASAP7_75t_R _30426_ (.A1(net6681),
    .A2(net155),
    .B(_07795_),
    .Y(_01433_));
 NOR2x1_ASAP7_75t_R _30427_ (.A(net6681),
    .B(_00446_),
    .Y(_07796_));
 AO21x1_ASAP7_75t_R _30428_ (.A1(net6681),
    .A2(net156),
    .B(_07796_),
    .Y(_01434_));
 NOR2x1_ASAP7_75t_R _30429_ (.A(net6681),
    .B(_00553_),
    .Y(_07797_));
 AO21x1_ASAP7_75t_R _30430_ (.A1(net6681),
    .A2(net157),
    .B(_07797_),
    .Y(_01435_));
 NOR2x1_ASAP7_75t_R _30432_ (.A(net6682),
    .B(_00552_),
    .Y(_07799_));
 AO21x1_ASAP7_75t_R _30433_ (.A1(net6682),
    .A2(net158),
    .B(_07799_),
    .Y(_01436_));
 NOR2x1_ASAP7_75t_R _30434_ (.A(net6681),
    .B(_00551_),
    .Y(_07800_));
 AO21x1_ASAP7_75t_R _30435_ (.A1(net6681),
    .A2(net159),
    .B(_07800_),
    .Y(_01437_));
 NOR2x1_ASAP7_75t_R _30437_ (.A(net6681),
    .B(_00550_),
    .Y(_07802_));
 AO21x1_ASAP7_75t_R _30438_ (.A1(net6681),
    .A2(net160),
    .B(_07802_),
    .Y(_01438_));
 NOR2x1_ASAP7_75t_R _30439_ (.A(net6681),
    .B(_00549_),
    .Y(_07803_));
 AO21x1_ASAP7_75t_R _30440_ (.A1(net6681),
    .A2(net161),
    .B(_07803_),
    .Y(_01439_));
 NOR2x1_ASAP7_75t_R _30441_ (.A(net6684),
    .B(_00548_),
    .Y(_07804_));
 AO21x1_ASAP7_75t_R _30442_ (.A1(net6684),
    .A2(net162),
    .B(_07804_),
    .Y(_01440_));
 NOR2x1_ASAP7_75t_R _30443_ (.A(net6684),
    .B(_00547_),
    .Y(_07805_));
 AO21x1_ASAP7_75t_R _30444_ (.A1(net6684),
    .A2(net163),
    .B(_07805_),
    .Y(_01441_));
 NOR2x1_ASAP7_75t_R _30445_ (.A(net6684),
    .B(_00546_),
    .Y(_07806_));
 AO21x1_ASAP7_75t_R _30446_ (.A1(net6684),
    .A2(net164),
    .B(_07806_),
    .Y(_01442_));
 NOR2x1_ASAP7_75t_R _30447_ (.A(net6684),
    .B(_00545_),
    .Y(_07807_));
 AO21x1_ASAP7_75t_R _30448_ (.A1(net6684),
    .A2(net165),
    .B(_07807_),
    .Y(_01443_));
 NOR2x1_ASAP7_75t_R _30449_ (.A(net6689),
    .B(_00466_),
    .Y(_07808_));
 AO21x1_ASAP7_75t_R _30450_ (.A1(net6689),
    .A2(net166),
    .B(_07808_),
    .Y(_01444_));
 NOR2x1_ASAP7_75t_R _30451_ (.A(net6689),
    .B(_00465_),
    .Y(_07809_));
 AO21x1_ASAP7_75t_R _30452_ (.A1(net6689),
    .A2(net167),
    .B(_07809_),
    .Y(_01445_));
 NOR2x1_ASAP7_75t_R _30454_ (.A(net6689),
    .B(_00467_),
    .Y(_07811_));
 AO21x1_ASAP7_75t_R _30455_ (.A1(net6689),
    .A2(net168),
    .B(_07811_),
    .Y(_01446_));
 NOR2x1_ASAP7_75t_R _30456_ (.A(net6689),
    .B(_00544_),
    .Y(_07812_));
 AO21x1_ASAP7_75t_R _30457_ (.A1(net6689),
    .A2(net169),
    .B(_07812_),
    .Y(_01447_));
 NOR2x1_ASAP7_75t_R _30459_ (.A(net6684),
    .B(_00408_),
    .Y(_07814_));
 AO21x1_ASAP7_75t_R _30460_ (.A1(net6684),
    .A2(net170),
    .B(_07814_),
    .Y(_01448_));
 NOR2x1_ASAP7_75t_R _30461_ (.A(net6689),
    .B(_00543_),
    .Y(_07815_));
 AO21x1_ASAP7_75t_R _30462_ (.A1(net6689),
    .A2(net171),
    .B(_07815_),
    .Y(_01449_));
 NOR2x1_ASAP7_75t_R _30463_ (.A(net6689),
    .B(_00542_),
    .Y(_07816_));
 AO21x1_ASAP7_75t_R _30464_ (.A1(net6689),
    .A2(net172),
    .B(_07816_),
    .Y(_01450_));
 NOR2x1_ASAP7_75t_R _30465_ (.A(net6689),
    .B(_00541_),
    .Y(_07817_));
 AO21x1_ASAP7_75t_R _30466_ (.A1(net6689),
    .A2(net173),
    .B(_07817_),
    .Y(_01451_));
 NOR2x1_ASAP7_75t_R _30467_ (.A(net6689),
    .B(_00540_),
    .Y(_07818_));
 AO21x1_ASAP7_75t_R _30468_ (.A1(net6689),
    .A2(net174),
    .B(_07818_),
    .Y(_01452_));
 NOR2x1_ASAP7_75t_R _30469_ (.A(net6689),
    .B(_00454_),
    .Y(_07819_));
 AO21x1_ASAP7_75t_R _30470_ (.A1(net6689),
    .A2(net175),
    .B(_07819_),
    .Y(_01453_));
 NOR2x1_ASAP7_75t_R _30471_ (.A(net6689),
    .B(_00453_),
    .Y(_07820_));
 AO21x1_ASAP7_75t_R _30472_ (.A1(net6689),
    .A2(net176),
    .B(_07820_),
    .Y(_01454_));
 NOR2x1_ASAP7_75t_R _30473_ (.A(net6689),
    .B(_00455_),
    .Y(_07821_));
 AO21x1_ASAP7_75t_R _30474_ (.A1(net6689),
    .A2(net177),
    .B(_07821_),
    .Y(_01455_));
 NOR2x1_ASAP7_75t_R _30476_ (.A(net6689),
    .B(_00539_),
    .Y(_07823_));
 AO21x1_ASAP7_75t_R _30477_ (.A1(net6689),
    .A2(net178),
    .B(_07823_),
    .Y(_01456_));
 NOR2x1_ASAP7_75t_R _30478_ (.A(net6689),
    .B(_00538_),
    .Y(_07824_));
 AO21x1_ASAP7_75t_R _30479_ (.A1(net6689),
    .A2(net179),
    .B(_07824_),
    .Y(_01457_));
 NOR2x1_ASAP7_75t_R _30481_ (.A(net6689),
    .B(_00537_),
    .Y(_07826_));
 AO21x1_ASAP7_75t_R _30482_ (.A1(net6689),
    .A2(net180),
    .B(_07826_),
    .Y(_01458_));
 NOR2x1_ASAP7_75t_R _30483_ (.A(net6680),
    .B(_00410_),
    .Y(_07827_));
 AO21x1_ASAP7_75t_R _30484_ (.A1(net6680),
    .A2(net181),
    .B(_07827_),
    .Y(_01459_));
 NOR2x1_ASAP7_75t_R _30485_ (.A(net6684),
    .B(_00536_),
    .Y(_07828_));
 AO21x1_ASAP7_75t_R _30486_ (.A1(net6684),
    .A2(net182),
    .B(_07828_),
    .Y(_01460_));
 NOR2x1_ASAP7_75t_R _30487_ (.A(net6689),
    .B(_00535_),
    .Y(_07829_));
 AO21x1_ASAP7_75t_R _30488_ (.A1(net6689),
    .A2(net183),
    .B(_07829_),
    .Y(_01461_));
 NOR2x1_ASAP7_75t_R _30489_ (.A(net6683),
    .B(_00406_),
    .Y(_07830_));
 AO21x1_ASAP7_75t_R _30490_ (.A1(net6683),
    .A2(net184),
    .B(_07830_),
    .Y(_01462_));
 NOR2x1_ASAP7_75t_R _30491_ (.A(net6680),
    .B(_00405_),
    .Y(_07831_));
 AO21x1_ASAP7_75t_R _30492_ (.A1(net6680),
    .A2(net185),
    .B(_07831_),
    .Y(_01463_));
 NOR2x1_ASAP7_75t_R _30493_ (.A(net6680),
    .B(_00407_),
    .Y(_07832_));
 AO21x1_ASAP7_75t_R _30494_ (.A1(net6680),
    .A2(net186),
    .B(_07832_),
    .Y(_01464_));
 NOR2x1_ASAP7_75t_R _30495_ (.A(net6686),
    .B(_00534_),
    .Y(_07833_));
 AO21x1_ASAP7_75t_R _30496_ (.A1(net6686),
    .A2(net187),
    .B(_07833_),
    .Y(_01465_));
 NOR2x1_ASAP7_75t_R _30498_ (.A(net6684),
    .B(_00533_),
    .Y(_07835_));
 AO21x1_ASAP7_75t_R _30499_ (.A1(net6684),
    .A2(net188),
    .B(_07835_),
    .Y(_01466_));
 NOR2x1_ASAP7_75t_R _30500_ (.A(net6684),
    .B(_00532_),
    .Y(_07836_));
 AO21x1_ASAP7_75t_R _30501_ (.A1(net6684),
    .A2(net189),
    .B(_07836_),
    .Y(_01467_));
 NOR2x1_ASAP7_75t_R _30503_ (.A(net6680),
    .B(_00531_),
    .Y(_07838_));
 AO21x1_ASAP7_75t_R _30504_ (.A1(net6680),
    .A2(net190),
    .B(_07838_),
    .Y(_01468_));
 NOR2x1_ASAP7_75t_R _30505_ (.A(net6684),
    .B(_00530_),
    .Y(_07839_));
 AO21x1_ASAP7_75t_R _30506_ (.A1(net6684),
    .A2(net191),
    .B(_07839_),
    .Y(_01469_));
 NOR2x1_ASAP7_75t_R _30507_ (.A(net6689),
    .B(_00529_),
    .Y(_07840_));
 AO21x1_ASAP7_75t_R _30508_ (.A1(net6689),
    .A2(net192),
    .B(_07840_),
    .Y(_01470_));
 NOR2x1_ASAP7_75t_R _30509_ (.A(net6680),
    .B(_00475_),
    .Y(_07841_));
 AO21x1_ASAP7_75t_R _30510_ (.A1(net6680),
    .A2(net193),
    .B(_07841_),
    .Y(_01471_));
 NOR2x1_ASAP7_75t_R _30511_ (.A(net6680),
    .B(_00474_),
    .Y(_07842_));
 AO21x1_ASAP7_75t_R _30512_ (.A1(net6680),
    .A2(net194),
    .B(_07842_),
    .Y(_01472_));
 NOR2x1_ASAP7_75t_R _30513_ (.A(net6680),
    .B(_00476_),
    .Y(_07843_));
 AO21x1_ASAP7_75t_R _30514_ (.A1(net6680),
    .A2(net195),
    .B(_07843_),
    .Y(_01473_));
 NOR2x1_ASAP7_75t_R _30515_ (.A(net6680),
    .B(_00528_),
    .Y(_07844_));
 AO21x1_ASAP7_75t_R _30516_ (.A1(net6680),
    .A2(net196),
    .B(_07844_),
    .Y(_01474_));
 NOR2x1_ASAP7_75t_R _30517_ (.A(net6680),
    .B(_00527_),
    .Y(_07845_));
 AO21x1_ASAP7_75t_R _30518_ (.A1(net6680),
    .A2(net197),
    .B(_07845_),
    .Y(_01475_));
 NOR2x1_ASAP7_75t_R _30520_ (.A(net6680),
    .B(_00526_),
    .Y(_07847_));
 AO21x1_ASAP7_75t_R _30521_ (.A1(net6680),
    .A2(net198),
    .B(_07847_),
    .Y(_01476_));
 NOR2x1_ASAP7_75t_R _30522_ (.A(net6680),
    .B(_00525_),
    .Y(_07848_));
 AO21x1_ASAP7_75t_R _30523_ (.A1(net6680),
    .A2(net199),
    .B(_07848_),
    .Y(_01477_));
 NOR2x1_ASAP7_75t_R _30525_ (.A(net6680),
    .B(_00524_),
    .Y(_07850_));
 AO21x1_ASAP7_75t_R _30526_ (.A1(net6680),
    .A2(net200),
    .B(_07850_),
    .Y(_01478_));
 NOR2x1_ASAP7_75t_R _30527_ (.A(net6681),
    .B(_00463_),
    .Y(_07851_));
 AO21x1_ASAP7_75t_R _30528_ (.A1(net6681),
    .A2(net201),
    .B(_07851_),
    .Y(_01479_));
 NOR2x1_ASAP7_75t_R _30529_ (.A(net6680),
    .B(_00462_),
    .Y(_07852_));
 AO21x1_ASAP7_75t_R _30530_ (.A1(net6680),
    .A2(net202),
    .B(_07852_),
    .Y(_01480_));
 NOR2x1_ASAP7_75t_R _30531_ (.A(net6680),
    .B(_00523_),
    .Y(_07853_));
 AO21x1_ASAP7_75t_R _30532_ (.A1(net6680),
    .A2(net203),
    .B(_07853_),
    .Y(_01481_));
 NOR2x1_ASAP7_75t_R _30533_ (.A(net6689),
    .B(_00464_),
    .Y(_07854_));
 AO21x1_ASAP7_75t_R _30534_ (.A1(net6689),
    .A2(net204),
    .B(_07854_),
    .Y(_01482_));
 NOR2x1_ASAP7_75t_R _30535_ (.A(net6681),
    .B(_00522_),
    .Y(_07855_));
 AO21x1_ASAP7_75t_R _30536_ (.A1(net6681),
    .A2(net205),
    .B(_07855_),
    .Y(_01483_));
 NOR2x1_ASAP7_75t_R _30537_ (.A(net6682),
    .B(_00521_),
    .Y(_07856_));
 AO21x1_ASAP7_75t_R _30538_ (.A1(net6682),
    .A2(net206),
    .B(_07856_),
    .Y(_01484_));
 NOR2x1_ASAP7_75t_R _30539_ (.A(net6682),
    .B(_00520_),
    .Y(_07857_));
 AO21x1_ASAP7_75t_R _30540_ (.A1(net6682),
    .A2(net207),
    .B(_07857_),
    .Y(_01485_));
 NOR2x1_ASAP7_75t_R _30542_ (.A(net6680),
    .B(_00519_),
    .Y(_07859_));
 AO21x1_ASAP7_75t_R _30543_ (.A1(net6680),
    .A2(net208),
    .B(_07859_),
    .Y(_01486_));
 NOR2x1_ASAP7_75t_R _30544_ (.A(net6682),
    .B(_00518_),
    .Y(_07860_));
 AO21x1_ASAP7_75t_R _30545_ (.A1(net6683),
    .A2(net209),
    .B(_07860_),
    .Y(_01487_));
 NOR2x1_ASAP7_75t_R _30547_ (.A(net6680),
    .B(_00451_),
    .Y(_07862_));
 AO21x1_ASAP7_75t_R _30548_ (.A1(net6680),
    .A2(net210),
    .B(_07862_),
    .Y(_01488_));
 NOR2x1_ASAP7_75t_R _30549_ (.A(net6680),
    .B(_00450_),
    .Y(_07863_));
 AO21x1_ASAP7_75t_R _30550_ (.A1(net6680),
    .A2(net211),
    .B(_07863_),
    .Y(_01489_));
 NOR2x1_ASAP7_75t_R _30551_ (.A(net6683),
    .B(_00452_),
    .Y(_07864_));
 AO21x1_ASAP7_75t_R _30552_ (.A1(net6683),
    .A2(net212),
    .B(_07864_),
    .Y(_01490_));
 NOR2x1_ASAP7_75t_R _30553_ (.A(net6680),
    .B(_00517_),
    .Y(_07865_));
 AO21x1_ASAP7_75t_R _30554_ (.A1(net6680),
    .A2(net213),
    .B(_07865_),
    .Y(_01491_));
 NOR2x1_ASAP7_75t_R _30555_ (.A(net6686),
    .B(_00516_),
    .Y(_07866_));
 AO21x1_ASAP7_75t_R _30556_ (.A1(net6686),
    .A2(net214),
    .B(_07866_),
    .Y(_01492_));
 NOR2x1_ASAP7_75t_R _30557_ (.A(net6680),
    .B(_00515_),
    .Y(_07867_));
 AO21x1_ASAP7_75t_R _30558_ (.A1(net6680),
    .A2(net215),
    .B(_07867_),
    .Y(_01493_));
 NOR2x1_ASAP7_75t_R _30559_ (.A(net6680),
    .B(_00514_),
    .Y(_07868_));
 AO21x1_ASAP7_75t_R _30560_ (.A1(net6680),
    .A2(net216),
    .B(_07868_),
    .Y(_01494_));
 NOR2x1_ASAP7_75t_R _30561_ (.A(net6680),
    .B(_00513_),
    .Y(_07869_));
 AO21x1_ASAP7_75t_R _30562_ (.A1(net6680),
    .A2(net217),
    .B(_07869_),
    .Y(_01495_));
 NOR2x1_ASAP7_75t_R _30564_ (.A(net6683),
    .B(_00512_),
    .Y(_07871_));
 AO21x1_ASAP7_75t_R _30565_ (.A1(net6683),
    .A2(net218),
    .B(_07871_),
    .Y(_01496_));
 NOR2x1_ASAP7_75t_R _30566_ (.A(net6682),
    .B(_00484_),
    .Y(_07872_));
 AO21x1_ASAP7_75t_R _30567_ (.A1(net6682),
    .A2(net219),
    .B(_07872_),
    .Y(_01497_));
 NOR2x1_ASAP7_75t_R _30569_ (.A(net6682),
    .B(_00483_),
    .Y(_07874_));
 AO21x1_ASAP7_75t_R _30570_ (.A1(net6682),
    .A2(net220),
    .B(_07874_),
    .Y(_01498_));
 NOR2x1_ASAP7_75t_R _30571_ (.A(net6681),
    .B(_00485_),
    .Y(_07875_));
 AO21x1_ASAP7_75t_R _30572_ (.A1(net6681),
    .A2(net221),
    .B(_07875_),
    .Y(_01499_));
 NOR2x1_ASAP7_75t_R _30573_ (.A(net6681),
    .B(_00511_),
    .Y(_07876_));
 AO21x1_ASAP7_75t_R _30574_ (.A1(net6681),
    .A2(net222),
    .B(_07876_),
    .Y(_01500_));
 NOR2x1_ASAP7_75t_R _30575_ (.A(net6681),
    .B(_00510_),
    .Y(_07877_));
 AO21x1_ASAP7_75t_R _30576_ (.A1(net6681),
    .A2(net223),
    .B(_07877_),
    .Y(_01501_));
 NOR2x1_ASAP7_75t_R _30577_ (.A(net6681),
    .B(_00509_),
    .Y(_07878_));
 AO21x1_ASAP7_75t_R _30578_ (.A1(net6681),
    .A2(net224),
    .B(_07878_),
    .Y(_01502_));
 NOR2x1_ASAP7_75t_R _30579_ (.A(net6681),
    .B(_00508_),
    .Y(_07879_));
 AO21x1_ASAP7_75t_R _30580_ (.A1(net6681),
    .A2(net225),
    .B(_07879_),
    .Y(_01503_));
 NOR2x1_ASAP7_75t_R _30581_ (.A(net6681),
    .B(_00507_),
    .Y(_07880_));
 AO21x1_ASAP7_75t_R _30582_ (.A1(net6681),
    .A2(net226),
    .B(_07880_),
    .Y(_01504_));
 NOR2x1_ASAP7_75t_R _30583_ (.A(net6681),
    .B(_00506_),
    .Y(_07881_));
 AO21x1_ASAP7_75t_R _30584_ (.A1(net6681),
    .A2(net227),
    .B(_07881_),
    .Y(_01505_));
 NOR2x1_ASAP7_75t_R _30586_ (.A(net6682),
    .B(_00472_),
    .Y(_07883_));
 AO21x1_ASAP7_75t_R _30587_ (.A1(net6682),
    .A2(net228),
    .B(_07883_),
    .Y(_01506_));
 NOR2x1_ASAP7_75t_R _30588_ (.A(net6682),
    .B(_00471_),
    .Y(_07884_));
 AO21x1_ASAP7_75t_R _30589_ (.A1(net6682),
    .A2(net229),
    .B(_07884_),
    .Y(_01507_));
 NOR2x1_ASAP7_75t_R _30591_ (.A(net6681),
    .B(_00473_),
    .Y(_07886_));
 AO21x1_ASAP7_75t_R _30592_ (.A1(net6681),
    .A2(net230),
    .B(_07886_),
    .Y(_01508_));
 NOR2x1_ASAP7_75t_R _30593_ (.A(net6681),
    .B(_00505_),
    .Y(_07887_));
 AO21x1_ASAP7_75t_R _30594_ (.A1(net6681),
    .A2(net231),
    .B(_07887_),
    .Y(_01509_));
 NOR2x1_ASAP7_75t_R _30595_ (.A(net6681),
    .B(_00504_),
    .Y(_07888_));
 AO21x1_ASAP7_75t_R _30596_ (.A1(net6681),
    .A2(net232),
    .B(_07888_),
    .Y(_01510_));
 NOR2x1_ASAP7_75t_R _30597_ (.A(net6681),
    .B(_00503_),
    .Y(_07889_));
 AO21x1_ASAP7_75t_R _30598_ (.A1(net6681),
    .A2(net233),
    .B(_07889_),
    .Y(_01511_));
 NOR2x1_ASAP7_75t_R _30599_ (.A(net6681),
    .B(_00502_),
    .Y(_07890_));
 AO21x1_ASAP7_75t_R _30600_ (.A1(net6681),
    .A2(net234),
    .B(_07890_),
    .Y(_01512_));
 NOR2x1_ASAP7_75t_R _30601_ (.A(net6681),
    .B(_00501_),
    .Y(_07891_));
 AO21x1_ASAP7_75t_R _30602_ (.A1(net6681),
    .A2(net235),
    .B(_07891_),
    .Y(_01513_));
 NOR2x1_ASAP7_75t_R _30603_ (.A(net6681),
    .B(_00500_),
    .Y(_07892_));
 AO21x1_ASAP7_75t_R _30604_ (.A1(net6681),
    .A2(net236),
    .B(_07892_),
    .Y(_01514_));
 NOR2x1_ASAP7_75t_R _30605_ (.A(net6681),
    .B(_00460_),
    .Y(_07893_));
 AO21x1_ASAP7_75t_R _30606_ (.A1(net6681),
    .A2(net237),
    .B(_07893_),
    .Y(_01515_));
 NOR2x1_ASAP7_75t_R _30608_ (.A(net6681),
    .B(_00459_),
    .Y(_07895_));
 AO21x1_ASAP7_75t_R _30609_ (.A1(net6681),
    .A2(net238),
    .B(_07895_),
    .Y(_01516_));
 NOR2x1_ASAP7_75t_R _30610_ (.A(net6681),
    .B(_00461_),
    .Y(_07896_));
 AO21x1_ASAP7_75t_R _30611_ (.A1(net6681),
    .A2(net239),
    .B(_07896_),
    .Y(_01517_));
 NOR2x1_ASAP7_75t_R _30613_ (.A(net6681),
    .B(_00499_),
    .Y(_07898_));
 AO21x1_ASAP7_75t_R _30614_ (.A1(net6681),
    .A2(net240),
    .B(_07898_),
    .Y(_01518_));
 NOR2x1_ASAP7_75t_R _30615_ (.A(net6681),
    .B(_00498_),
    .Y(_07899_));
 AO21x1_ASAP7_75t_R _30616_ (.A1(net6681),
    .A2(net241),
    .B(_07899_),
    .Y(_01519_));
 NOR2x1_ASAP7_75t_R _30617_ (.A(net6681),
    .B(_00497_),
    .Y(_07900_));
 AO21x1_ASAP7_75t_R _30618_ (.A1(net6681),
    .A2(net242),
    .B(_07900_),
    .Y(_01520_));
 NOR2x1_ASAP7_75t_R _30619_ (.A(net6681),
    .B(_00496_),
    .Y(_07901_));
 AO21x1_ASAP7_75t_R _30620_ (.A1(net6681),
    .A2(net243),
    .B(_07901_),
    .Y(_01521_));
 NOR2x1_ASAP7_75t_R _30621_ (.A(net6681),
    .B(_00495_),
    .Y(_07902_));
 AO21x1_ASAP7_75t_R _30622_ (.A1(net6681),
    .A2(net244),
    .B(_07902_),
    .Y(_01522_));
 NOR2x1_ASAP7_75t_R _30623_ (.A(net6681),
    .B(_00448_),
    .Y(_07903_));
 AO21x1_ASAP7_75t_R _30624_ (.A1(net6681),
    .A2(net245),
    .B(_07903_),
    .Y(_01523_));
 NOR2x1_ASAP7_75t_R _30625_ (.A(net6681),
    .B(_00447_),
    .Y(_07904_));
 AO21x1_ASAP7_75t_R _30626_ (.A1(net6681),
    .A2(net246),
    .B(_07904_),
    .Y(_01524_));
 NOR2x1_ASAP7_75t_R _30627_ (.A(net6682),
    .B(_00478_),
    .Y(_07905_));
 AO21x1_ASAP7_75t_R _30628_ (.A1(net6682),
    .A2(net247),
    .B(_07905_),
    .Y(_01525_));
 NOR2x1_ASAP7_75t_R _30630_ (.A(net6681),
    .B(_00449_),
    .Y(_07907_));
 AO21x1_ASAP7_75t_R _30631_ (.A1(net6681),
    .A2(net248),
    .B(_07907_),
    .Y(_01526_));
 NOR2x1_ASAP7_75t_R _30632_ (.A(net6681),
    .B(_00494_),
    .Y(_07908_));
 AO21x1_ASAP7_75t_R _30633_ (.A1(net6681),
    .A2(net249),
    .B(_07908_),
    .Y(_01527_));
 NOR2x1_ASAP7_75t_R _30634_ (.A(net6681),
    .B(_00493_),
    .Y(_07909_));
 AO21x1_ASAP7_75t_R _30635_ (.A1(net6681),
    .A2(net250),
    .B(_07909_),
    .Y(_01528_));
 NOR2x1_ASAP7_75t_R _30636_ (.A(net6681),
    .B(_00492_),
    .Y(_07910_));
 AO21x1_ASAP7_75t_R _30637_ (.A1(net6681),
    .A2(net251),
    .B(_07910_),
    .Y(_01529_));
 NOR2x1_ASAP7_75t_R _30638_ (.A(net6681),
    .B(_00491_),
    .Y(_07911_));
 AO21x1_ASAP7_75t_R _30639_ (.A1(net6681),
    .A2(net252),
    .B(_07911_),
    .Y(_01530_));
 NOR2x1_ASAP7_75t_R _30640_ (.A(net6681),
    .B(_00490_),
    .Y(_07912_));
 AO21x1_ASAP7_75t_R _30641_ (.A1(net6681),
    .A2(net253),
    .B(_07912_),
    .Y(_01531_));
 NOR2x1_ASAP7_75t_R _30642_ (.A(net6681),
    .B(_00481_),
    .Y(_07913_));
 AO21x1_ASAP7_75t_R _30643_ (.A1(net6681),
    .A2(net254),
    .B(_07913_),
    .Y(_01532_));
 NOR2x1_ASAP7_75t_R _30644_ (.A(net6681),
    .B(_00480_),
    .Y(_07914_));
 AO21x1_ASAP7_75t_R _30645_ (.A1(net6681),
    .A2(net255),
    .B(_07914_),
    .Y(_01533_));
 NOR2x1_ASAP7_75t_R _30646_ (.A(net6681),
    .B(_00482_),
    .Y(_07915_));
 AO21x1_ASAP7_75t_R _30647_ (.A1(net6681),
    .A2(net256),
    .B(_07915_),
    .Y(_01534_));
 NOR2x1_ASAP7_75t_R _30648_ (.A(net6681),
    .B(_00489_),
    .Y(_07916_));
 AO21x1_ASAP7_75t_R _30649_ (.A1(net6681),
    .A2(net257),
    .B(_07916_),
    .Y(_01535_));
 NOR2x1_ASAP7_75t_R _30650_ (.A(net6690),
    .B(_00477_),
    .Y(_07917_));
 AO21x1_ASAP7_75t_R _30651_ (.A1(net6690),
    .A2(net258),
    .B(_07917_),
    .Y(_01536_));
 AND3x1_ASAP7_75t_R _30652_ (.A(_00570_),
    .B(_00571_),
    .C(_00572_),
    .Y(_07918_));
 AOI21x1_ASAP7_75t_R _30653_ (.A1(_00571_),
    .A2(_00572_),
    .B(_00570_),
    .Y(_07919_));
 INVx1_ASAP7_75t_R _30654_ (.A(net130),
    .Y(_07920_));
 AOI21x1_ASAP7_75t_R _30655_ (.A1(_00411_),
    .A2(_07918_),
    .B(_07920_),
    .Y(_07921_));
 OA211x2_ASAP7_75t_R _30656_ (.A1(_07918_),
    .A2(_07919_),
    .B(_07921_),
    .C(net6679),
    .Y(_01407_));
 XNOR2x2_ASAP7_75t_R _30657_ (.A(_00487_),
    .B(_00971_),
    .Y(_07922_));
 INVx1_ASAP7_75t_R _30658_ (.A(_07922_),
    .Y(_07923_));
 OAI21x1_ASAP7_75t_R _30659_ (.A1(_00970_),
    .A2(_07923_),
    .B(net6678),
    .Y(_01537_));
 OR3x1_ASAP7_75t_R _30660_ (.A(_00487_),
    .B(_00965_),
    .C(\u0.r0.rcnt_next[0] ),
    .Y(_07924_));
 XOR2x2_ASAP7_75t_R _30661_ (.A(_07924_),
    .B(_00829_),
    .Y(_07925_));
 OR3x1_ASAP7_75t_R _30662_ (.A(_07925_),
    .B(_00966_),
    .C(_07923_),
    .Y(_07926_));
 INVx1_ASAP7_75t_R _30663_ (.A(_07925_),
    .Y(_07927_));
 INVx1_ASAP7_75t_R _30664_ (.A(_00967_),
    .Y(_07928_));
 OR3x1_ASAP7_75t_R _30665_ (.A(_07927_),
    .B(_07928_),
    .C(_07923_),
    .Y(_07929_));
 AOI21x1_ASAP7_75t_R _30666_ (.A1(_07926_),
    .A2(_07929_),
    .B(net6688),
    .Y(_01538_));
 OR3x1_ASAP7_75t_R _30667_ (.A(_07925_),
    .B(_00969_),
    .C(_07923_),
    .Y(_07930_));
 OR3x1_ASAP7_75t_R _30668_ (.A(_07927_),
    .B(_00966_),
    .C(_07923_),
    .Y(_07931_));
 AOI21x1_ASAP7_75t_R _30669_ (.A1(_07930_),
    .A2(_07931_),
    .B(net6688),
    .Y(_01539_));
 OR3x1_ASAP7_75t_R _30670_ (.A(_07925_),
    .B(_00968_),
    .C(_07923_),
    .Y(_07932_));
 OR3x1_ASAP7_75t_R _30671_ (.A(_07927_),
    .B(_00970_),
    .C(_07923_),
    .Y(_07933_));
 AOI21x1_ASAP7_75t_R _30672_ (.A1(_07932_),
    .A2(_07933_),
    .B(net6688),
    .Y(_01540_));
 OR3x1_ASAP7_75t_R _30673_ (.A(_07925_),
    .B(_00970_),
    .C(_07922_),
    .Y(_07934_));
 AOI21x1_ASAP7_75t_R _30674_ (.A1(_07934_),
    .A2(_07929_),
    .B(net6688),
    .Y(_01541_));
 OR3x1_ASAP7_75t_R _30675_ (.A(_07925_),
    .B(_00966_),
    .C(_07922_),
    .Y(_07935_));
 AOI21x1_ASAP7_75t_R _30676_ (.A1(_07935_),
    .A2(_07931_),
    .B(net6688),
    .Y(_01542_));
 INVx1_ASAP7_75t_R _30677_ (.A(_00969_),
    .Y(_07936_));
 NOR2x1_ASAP7_75t_R _30678_ (.A(net6688),
    .B(_07922_),
    .Y(_01547_));
 AND3x1_ASAP7_75t_R _30679_ (.A(_07927_),
    .B(_07936_),
    .C(_01547_),
    .Y(_01543_));
 INVx1_ASAP7_75t_R _30680_ (.A(_00968_),
    .Y(_07937_));
 AND3x1_ASAP7_75t_R _30681_ (.A(_07927_),
    .B(_07937_),
    .C(_01547_),
    .Y(_01544_));
 NOR2x1_ASAP7_75t_R _30682_ (.A(net6688),
    .B(\u0.r0.rcnt[0] ),
    .Y(_01545_));
 NOR2x1_ASAP7_75t_R _30683_ (.A(net6688),
    .B(_00967_),
    .Y(_01546_));
 NOR2x1_ASAP7_75t_R _30684_ (.A(net6688),
    .B(_07927_),
    .Y(_01548_));
 AO22x1_ASAP7_75t_R _30685_ (.A1(net6689),
    .A2(net130),
    .B1(_07921_),
    .B2(_00572_),
    .Y(_01405_));
 OA21x2_ASAP7_75t_R _30686_ (.A1(_00571_),
    .A2(_00572_),
    .B(net6679),
    .Y(_07938_));
 NAND2x1_ASAP7_75t_R _30687_ (.A(_00571_),
    .B(_00572_),
    .Y(_07939_));
 AO21x1_ASAP7_75t_R _30688_ (.A1(_00411_),
    .A2(_00570_),
    .B(_07939_),
    .Y(_07940_));
 AOI21x1_ASAP7_75t_R _30689_ (.A1(_07938_),
    .A2(_07940_),
    .B(_07920_),
    .Y(_01406_));
 NOR2x1_ASAP7_75t_R _30690_ (.A(_00411_),
    .B(_07918_),
    .Y(_07941_));
 OA21x2_ASAP7_75t_R _30691_ (.A1(_07941_),
    .A2(net6689),
    .B(net130),
    .Y(_01408_));
 HAxp5_ASAP7_75t_R _30692_ (.A(\u0.r0.rcnt_next[0] ),
    .B(_00965_),
    .CON(_00966_),
    .SN(_00967_));
 HAxp5_ASAP7_75t_R _30693_ (.A(\u0.r0.rcnt_next[0] ),
    .B(\u0.r0.rcnt[1] ),
    .CON(_00968_),
    .SN(_15602_));
 HAxp5_ASAP7_75t_R _30694_ (.A(\u0.r0.rcnt[0] ),
    .B(_00965_),
    .CON(_00969_),
    .SN(_15603_));
 HAxp5_ASAP7_75t_R _30695_ (.A(\u0.r0.rcnt[0] ),
    .B(\u0.r0.rcnt[1] ),
    .CON(_00970_),
    .SN(_15604_));
 HAxp5_ASAP7_75t_R _30696_ (.A(\u0.r0.rcnt[0] ),
    .B(\u0.r0.rcnt[1] ),
    .CON(_00971_),
    .SN(_15605_));
 HAxp5_ASAP7_75t_R _30697_ (.A(_00973_),
    .B(_00972_),
    .CON(_00974_),
    .SN(_00975_));
 HAxp5_ASAP7_75t_R _30698_ (.A(_00972_),
    .B(net5981),
    .CON(_00976_),
    .SN(_15606_));
 HAxp5_ASAP7_75t_R _30699_ (.A(net5982),
    .B(net6340),
    .CON(_00978_),
    .SN(_15607_));
 HAxp5_ASAP7_75t_R _30700_ (.A(_00972_),
    .B(net6340),
    .CON(_00979_),
    .SN(_15608_));
 HAxp5_ASAP7_75t_R _30701_ (.A(net6337),
    .B(net5981),
    .CON(_00981_),
    .SN(_15609_));
 HAxp5_ASAP7_75t_R _30702_ (.A(net6337),
    .B(net5981),
    .CON(_00982_),
    .SN(_15610_));
 HAxp5_ASAP7_75t_R _30703_ (.A(net6337),
    .B(net6340),
    .CON(_00983_),
    .SN(_15611_));
 HAxp5_ASAP7_75t_R _30704_ (.A(net6337),
    .B(net6340),
    .CON(_00984_),
    .SN(_15612_));
 HAxp5_ASAP7_75t_R _30705_ (.A(net5982),
    .B(net6371),
    .CON(_00986_),
    .SN(_00987_));
 HAxp5_ASAP7_75t_R _30706_ (.A(net5982),
    .B(net6372),
    .CON(_00988_),
    .SN(_15613_));
 HAxp5_ASAP7_75t_R _30707_ (.A(net5982),
    .B(net6339),
    .CON(_00990_),
    .SN(_15614_));
 HAxp5_ASAP7_75t_R _30708_ (.A(net5983),
    .B(net6338),
    .CON(_00991_),
    .SN(_15615_));
 HAxp5_ASAP7_75t_R _30709_ (.A(net6337),
    .B(net6373),
    .CON(_00992_),
    .SN(_15616_));
 HAxp5_ASAP7_75t_R _30710_ (.A(net6337),
    .B(net6369),
    .CON(_00993_),
    .SN(_15617_));
 HAxp5_ASAP7_75t_R _30711_ (.A(net6337),
    .B(net6338),
    .CON(_00994_),
    .SN(_15618_));
 HAxp5_ASAP7_75t_R _30712_ (.A(_08950_),
    .B(_00995_),
    .CON(_00997_),
    .SN(_00998_));
 HAxp5_ASAP7_75t_R _30713_ (.A(net5931),
    .B(net6310),
    .CON(_00999_),
    .SN(_15619_));
 HAxp5_ASAP7_75t_R _30714_ (.A(net5931),
    .B(_01000_),
    .CON(_01001_),
    .SN(_15620_));
 HAxp5_ASAP7_75t_R _30715_ (.A(net5931),
    .B(_01000_),
    .CON(_01002_),
    .SN(_15621_));
 HAxp5_ASAP7_75t_R _30716_ (.A(net6309),
    .B(net6311),
    .CON(_01004_),
    .SN(_15622_));
 HAxp5_ASAP7_75t_R _30717_ (.A(net6309),
    .B(net6311),
    .CON(_01005_),
    .SN(_15623_));
 HAxp5_ASAP7_75t_R _30718_ (.A(net6309),
    .B(_01000_),
    .CON(_01006_),
    .SN(_15624_));
 HAxp5_ASAP7_75t_R _30719_ (.A(net6309),
    .B(_01000_),
    .CON(_01007_),
    .SN(_15625_));
 HAxp5_ASAP7_75t_R _30720_ (.A(net5931),
    .B(net6308),
    .CON(_01009_),
    .SN(_01010_));
 HAxp5_ASAP7_75t_R _30721_ (.A(net5931),
    .B(net6308),
    .CON(_01011_),
    .SN(_15626_));
 HAxp5_ASAP7_75t_R _30722_ (.A(net5931),
    .B(net5950),
    .CON(_01013_),
    .SN(_15627_));
 HAxp5_ASAP7_75t_R _30723_ (.A(net5931),
    .B(_08962_),
    .CON(_01014_),
    .SN(_15628_));
 HAxp5_ASAP7_75t_R _30724_ (.A(net6309),
    .B(net6308),
    .CON(_01015_),
    .SN(_15629_));
 HAxp5_ASAP7_75t_R _30725_ (.A(net6309),
    .B(net6308),
    .CON(_01016_),
    .SN(_15630_));
 HAxp5_ASAP7_75t_R _30726_ (.A(_09567_),
    .B(_08916_),
    .CON(_01019_),
    .SN(_01020_));
 HAxp5_ASAP7_75t_R _30727_ (.A(net6323),
    .B(net6296),
    .CON(_01021_),
    .SN(_15631_));
 HAxp5_ASAP7_75t_R _30728_ (.A(net6323),
    .B(_08911_),
    .CON(_01023_),
    .SN(_15632_));
 HAxp5_ASAP7_75t_R _30729_ (.A(net6323),
    .B(_08911_),
    .CON(_01024_),
    .SN(_15633_));
 HAxp5_ASAP7_75t_R _30730_ (.A(_01025_),
    .B(net6296),
    .CON(_01026_),
    .SN(_15634_));
 HAxp5_ASAP7_75t_R _30731_ (.A(_01025_),
    .B(net6296),
    .CON(_01027_),
    .SN(_15635_));
 HAxp5_ASAP7_75t_R _30732_ (.A(_01025_),
    .B(_08911_),
    .CON(_01028_),
    .SN(_15636_));
 HAxp5_ASAP7_75t_R _30733_ (.A(net5966),
    .B(_08911_),
    .CON(_01029_),
    .SN(_15637_));
 HAxp5_ASAP7_75t_R _30734_ (.A(net6323),
    .B(net6322),
    .CON(_01031_),
    .SN(_01032_));
 HAxp5_ASAP7_75t_R _30735_ (.A(net6323),
    .B(net6321),
    .CON(_01033_),
    .SN(_15638_));
 HAxp5_ASAP7_75t_R _30736_ (.A(net6323),
    .B(net5963),
    .CON(_01035_),
    .SN(_15639_));
 HAxp5_ASAP7_75t_R _30737_ (.A(net6323),
    .B(_08923_),
    .CON(_01036_),
    .SN(_15640_));
 HAxp5_ASAP7_75t_R _30738_ (.A(net5965),
    .B(net6322),
    .CON(_01037_),
    .SN(_15641_));
 HAxp5_ASAP7_75t_R _30739_ (.A(net5965),
    .B(net6322),
    .CON(_01038_),
    .SN(_15642_));
 HAxp5_ASAP7_75t_R _30740_ (.A(_10111_),
    .B(_08997_),
    .CON(_01041_),
    .SN(_01042_));
 HAxp5_ASAP7_75t_R _30741_ (.A(net6299),
    .B(net6287),
    .CON(_01043_),
    .SN(_15643_));
 HAxp5_ASAP7_75t_R _30742_ (.A(net6300),
    .B(_08992_),
    .CON(_01045_),
    .SN(_15644_));
 HAxp5_ASAP7_75t_R _30743_ (.A(net6300),
    .B(_08992_),
    .CON(_01046_),
    .SN(_15645_));
 HAxp5_ASAP7_75t_R _30744_ (.A(_01047_),
    .B(net6287),
    .CON(_01048_),
    .SN(_15646_));
 HAxp5_ASAP7_75t_R _30745_ (.A(_01047_),
    .B(net6287),
    .CON(_01049_),
    .SN(_15647_));
 HAxp5_ASAP7_75t_R _30746_ (.A(_01047_),
    .B(_08992_),
    .CON(_01050_),
    .SN(_15648_));
 HAxp5_ASAP7_75t_R _30747_ (.A(_01047_),
    .B(_08992_),
    .CON(_01051_),
    .SN(_15649_));
 HAxp5_ASAP7_75t_R _30748_ (.A(net6289),
    .B(net6299),
    .CON(_01053_),
    .SN(_01054_));
 HAxp5_ASAP7_75t_R _30749_ (.A(net6289),
    .B(net6299),
    .CON(_01055_),
    .SN(_15650_));
 HAxp5_ASAP7_75t_R _30750_ (.A(net5939),
    .B(net6300),
    .CON(_01057_),
    .SN(_15651_));
 HAxp5_ASAP7_75t_R _30751_ (.A(net5939),
    .B(net6299),
    .CON(_01058_),
    .SN(_15652_));
 HAxp5_ASAP7_75t_R _30752_ (.A(net5938),
    .B(net5940),
    .CON(_01059_),
    .SN(_15653_));
 HAxp5_ASAP7_75t_R _30753_ (.A(net5938),
    .B(net5940),
    .CON(_01060_),
    .SN(_15654_));
 HAxp5_ASAP7_75t_R _30754_ (.A(_10835_),
    .B(_10736_),
    .CON(_01063_),
    .SN(_01064_));
 HAxp5_ASAP7_75t_R _30755_ (.A(net5901),
    .B(net5894),
    .CON(_01065_),
    .SN(_15655_));
 HAxp5_ASAP7_75t_R _30756_ (.A(_10695_),
    .B(net5901),
    .CON(_01067_),
    .SN(_15656_));
 HAxp5_ASAP7_75t_R _30757_ (.A(_10715_),
    .B(net5894),
    .CON(_01069_),
    .SN(_15657_));
 HAxp5_ASAP7_75t_R _30758_ (.A(_10715_),
    .B(net5894),
    .CON(_01070_),
    .SN(_15658_));
 HAxp5_ASAP7_75t_R _30759_ (.A(net5907),
    .B(net5910),
    .CON(_01071_),
    .SN(_15659_));
 HAxp5_ASAP7_75t_R _30760_ (.A(_10715_),
    .B(_10695_),
    .CON(_01072_),
    .SN(_15660_));
 HAxp5_ASAP7_75t_R _30761_ (.A(net5899),
    .B(net5893),
    .CON(_01074_),
    .SN(_01075_));
 HAxp5_ASAP7_75t_R _30762_ (.A(net5899),
    .B(net5909),
    .CON(_01076_),
    .SN(_15661_));
 HAxp5_ASAP7_75t_R _30763_ (.A(net5899),
    .B(net5909),
    .CON(_01077_),
    .SN(_15662_));
 HAxp5_ASAP7_75t_R _30764_ (.A(net5905),
    .B(net5894),
    .CON(_01079_),
    .SN(_15663_));
 HAxp5_ASAP7_75t_R _30765_ (.A(net5905),
    .B(net5893),
    .CON(_01080_),
    .SN(_15664_));
 HAxp5_ASAP7_75t_R _30766_ (.A(net5905),
    .B(net5909),
    .CON(_01081_),
    .SN(_15665_));
 HAxp5_ASAP7_75t_R _30767_ (.A(_11553_),
    .B(_11446_),
    .CON(_01084_),
    .SN(_01085_));
 HAxp5_ASAP7_75t_R _30768_ (.A(net5882),
    .B(net5878),
    .CON(_01086_),
    .SN(_15666_));
 HAxp5_ASAP7_75t_R _30769_ (.A(net5882),
    .B(_11409_),
    .CON(_01088_),
    .SN(_15667_));
 HAxp5_ASAP7_75t_R _30770_ (.A(_11426_),
    .B(net5878),
    .CON(_01090_),
    .SN(_15668_));
 HAxp5_ASAP7_75t_R _30771_ (.A(_11426_),
    .B(net5878),
    .CON(_01091_),
    .SN(_15669_));
 HAxp5_ASAP7_75t_R _30772_ (.A(net5887),
    .B(net5891),
    .CON(_01092_),
    .SN(_15670_));
 HAxp5_ASAP7_75t_R _30773_ (.A(_11426_),
    .B(net5890),
    .CON(_01093_),
    .SN(_15671_));
 HAxp5_ASAP7_75t_R _30774_ (.A(net5524),
    .B(net5877),
    .CON(_01095_),
    .SN(_01096_));
 HAxp5_ASAP7_75t_R _30775_ (.A(net5524),
    .B(net5891),
    .CON(_01097_),
    .SN(_15672_));
 HAxp5_ASAP7_75t_R _30776_ (.A(net5524),
    .B(net5889),
    .CON(_01098_),
    .SN(_15673_));
 HAxp5_ASAP7_75t_R _30777_ (.A(_11443_),
    .B(net5877),
    .CON(_01100_),
    .SN(_15674_));
 HAxp5_ASAP7_75t_R _30778_ (.A(_11443_),
    .B(net5877),
    .CON(_01101_),
    .SN(_15675_));
 HAxp5_ASAP7_75t_R _30779_ (.A(net5883),
    .B(net5891),
    .CON(_01102_),
    .SN(_15676_));
 HAxp5_ASAP7_75t_R _30780_ (.A(_01104_),
    .B(_12178_),
    .CON(_01105_),
    .SN(_01106_));
 HAxp5_ASAP7_75t_R _30781_ (.A(net5870),
    .B(net5508),
    .CON(_01107_),
    .SN(_15677_));
 HAxp5_ASAP7_75t_R _30782_ (.A(net5870),
    .B(net5874),
    .CON(_01109_),
    .SN(_15678_));
 HAxp5_ASAP7_75t_R _30783_ (.A(_01110_),
    .B(net5508),
    .CON(_01111_),
    .SN(_15679_));
 HAxp5_ASAP7_75t_R _30784_ (.A(_01110_),
    .B(net5508),
    .CON(_01112_),
    .SN(_15680_));
 HAxp5_ASAP7_75t_R _30785_ (.A(net5873),
    .B(net5874),
    .CON(_01113_),
    .SN(_15681_));
 HAxp5_ASAP7_75t_R _30786_ (.A(_01110_),
    .B(net5874),
    .CON(_01114_),
    .SN(_15682_));
 HAxp5_ASAP7_75t_R _30787_ (.A(net5868),
    .B(net5507),
    .CON(_01116_),
    .SN(_01117_));
 HAxp5_ASAP7_75t_R _30788_ (.A(net5868),
    .B(net5874),
    .CON(_01118_),
    .SN(_15683_));
 HAxp5_ASAP7_75t_R _30789_ (.A(net5868),
    .B(net5874),
    .CON(_01119_),
    .SN(_15684_));
 HAxp5_ASAP7_75t_R _30790_ (.A(net5518),
    .B(net5507),
    .CON(_01121_),
    .SN(_15685_));
 HAxp5_ASAP7_75t_R _30791_ (.A(net5518),
    .B(net5507),
    .CON(_01122_),
    .SN(_15686_));
 HAxp5_ASAP7_75t_R _30792_ (.A(net5518),
    .B(net5874),
    .CON(_01123_),
    .SN(_15687_));
 HAxp5_ASAP7_75t_R _30793_ (.A(_01125_),
    .B(_12870_),
    .CON(_01126_),
    .SN(_01127_));
 HAxp5_ASAP7_75t_R _30794_ (.A(net5859),
    .B(net5496),
    .CON(_01128_),
    .SN(_15688_));
 HAxp5_ASAP7_75t_R _30795_ (.A(net5859),
    .B(net5864),
    .CON(_01130_),
    .SN(_15689_));
 HAxp5_ASAP7_75t_R _30796_ (.A(_12849_),
    .B(net5496),
    .CON(_01132_),
    .SN(_15690_));
 HAxp5_ASAP7_75t_R _30797_ (.A(_12849_),
    .B(net5496),
    .CON(_01133_),
    .SN(_15691_));
 HAxp5_ASAP7_75t_R _30798_ (.A(net5863),
    .B(net5864),
    .CON(_01134_),
    .SN(_15692_));
 HAxp5_ASAP7_75t_R _30799_ (.A(net5864),
    .B(_12849_),
    .CON(_01135_),
    .SN(_15693_));
 HAxp5_ASAP7_75t_R _30800_ (.A(net5857),
    .B(net5496),
    .CON(_01137_),
    .SN(_01138_));
 HAxp5_ASAP7_75t_R _30801_ (.A(net5857),
    .B(net5864),
    .CON(_01139_),
    .SN(_15694_));
 HAxp5_ASAP7_75t_R _30802_ (.A(net5857),
    .B(net5864),
    .CON(_01140_),
    .SN(_15695_));
 HAxp5_ASAP7_75t_R _30803_ (.A(net5861),
    .B(net5496),
    .CON(_01142_),
    .SN(_15696_));
 HAxp5_ASAP7_75t_R _30804_ (.A(net5862),
    .B(net5496),
    .CON(_01143_),
    .SN(_15697_));
 HAxp5_ASAP7_75t_R _30805_ (.A(net5860),
    .B(net5864),
    .CON(_01144_),
    .SN(_15698_));
 HAxp5_ASAP7_75t_R _30806_ (.A(_13634_),
    .B(_13576_),
    .CON(_01147_),
    .SN(_01148_));
 HAxp5_ASAP7_75t_R _30807_ (.A(net5483),
    .B(net6193),
    .CON(_01149_),
    .SN(_15699_));
 HAxp5_ASAP7_75t_R _30808_ (.A(net5484),
    .B(_13533_),
    .CON(_01151_),
    .SN(_15700_));
 HAxp5_ASAP7_75t_R _30809_ (.A(_01152_),
    .B(net6193),
    .CON(_01153_),
    .SN(_15701_));
 HAxp5_ASAP7_75t_R _30810_ (.A(_01152_),
    .B(net6193),
    .CON(_01154_),
    .SN(_15702_));
 HAxp5_ASAP7_75t_R _30811_ (.A(net5846),
    .B(net6197),
    .CON(_01155_),
    .SN(_15703_));
 HAxp5_ASAP7_75t_R _30812_ (.A(_01152_),
    .B(net6198),
    .CON(_01156_),
    .SN(_15704_));
 HAxp5_ASAP7_75t_R _30813_ (.A(net5482),
    .B(net6193),
    .CON(_01158_),
    .SN(_01159_));
 HAxp5_ASAP7_75t_R _30814_ (.A(net5482),
    .B(net6197),
    .CON(_01160_),
    .SN(_15705_));
 HAxp5_ASAP7_75t_R _30815_ (.A(net5480),
    .B(net6197),
    .CON(_01161_),
    .SN(_15706_));
 HAxp5_ASAP7_75t_R _30816_ (.A(net5487),
    .B(net6193),
    .CON(_01163_),
    .SN(_15707_));
 HAxp5_ASAP7_75t_R _30817_ (.A(net5487),
    .B(net6193),
    .CON(_01164_),
    .SN(_15708_));
 HAxp5_ASAP7_75t_R _30818_ (.A(net5487),
    .B(net6197),
    .CON(_01165_),
    .SN(_15709_));
 HAxp5_ASAP7_75t_R _30819_ (.A(_14272_),
    .B(_14263_),
    .CON(_01168_),
    .SN(_01169_));
 HAxp5_ASAP7_75t_R _30820_ (.A(net5817),
    .B(net6185),
    .CON(_01170_),
    .SN(_15710_));
 HAxp5_ASAP7_75t_R _30821_ (.A(net5817),
    .B(_14224_),
    .CON(_01172_),
    .SN(_15711_));
 HAxp5_ASAP7_75t_R _30822_ (.A(_14242_),
    .B(net6185),
    .CON(_01174_),
    .SN(_15712_));
 HAxp5_ASAP7_75t_R _30823_ (.A(_14242_),
    .B(net6185),
    .CON(_01175_),
    .SN(_15713_));
 HAxp5_ASAP7_75t_R _30824_ (.A(net5822),
    .B(net6191),
    .CON(_01176_),
    .SN(_15714_));
 HAxp5_ASAP7_75t_R _30825_ (.A(_14242_),
    .B(_14224_),
    .CON(_01177_),
    .SN(_15715_));
 HAxp5_ASAP7_75t_R _30826_ (.A(_14266_),
    .B(net6184),
    .CON(_01179_),
    .SN(_01180_));
 HAxp5_ASAP7_75t_R _30827_ (.A(net5814),
    .B(net6191),
    .CON(_01181_),
    .SN(_15716_));
 HAxp5_ASAP7_75t_R _30828_ (.A(net5815),
    .B(net6190),
    .CON(_01182_),
    .SN(_15717_));
 HAxp5_ASAP7_75t_R _30829_ (.A(net5818),
    .B(net6185),
    .CON(_01184_),
    .SN(_15718_));
 HAxp5_ASAP7_75t_R _30830_ (.A(net5821),
    .B(net6184),
    .CON(_01185_),
    .SN(_15719_));
 HAxp5_ASAP7_75t_R _30831_ (.A(net5818),
    .B(net6191),
    .CON(_01186_),
    .SN(_15720_));
 HAxp5_ASAP7_75t_R _30832_ (.A(_15161_),
    .B(_14971_),
    .CON(_01189_),
    .SN(_01190_));
 HAxp5_ASAP7_75t_R _30833_ (.A(net5778),
    .B(net6172),
    .CON(_01191_),
    .SN(_15721_));
 HAxp5_ASAP7_75t_R _30834_ (.A(net5778),
    .B(_14927_),
    .CON(_01193_),
    .SN(_15722_));
 HAxp5_ASAP7_75t_R _30835_ (.A(_01194_),
    .B(net6172),
    .CON(_01195_),
    .SN(_15723_));
 HAxp5_ASAP7_75t_R _30836_ (.A(_01194_),
    .B(net6172),
    .CON(_01196_),
    .SN(_15724_));
 HAxp5_ASAP7_75t_R _30837_ (.A(net5452),
    .B(net6179),
    .CON(_01197_),
    .SN(_15725_));
 HAxp5_ASAP7_75t_R _30838_ (.A(_01194_),
    .B(_14927_),
    .CON(_01198_),
    .SN(_15726_));
 HAxp5_ASAP7_75t_R _30839_ (.A(net5444),
    .B(net6172),
    .CON(_01200_),
    .SN(_01201_));
 HAxp5_ASAP7_75t_R _30840_ (.A(net5444),
    .B(net6178),
    .CON(_01202_),
    .SN(_15727_));
 HAxp5_ASAP7_75t_R _30841_ (.A(net5444),
    .B(net6178),
    .CON(_01203_),
    .SN(_15728_));
 HAxp5_ASAP7_75t_R _30842_ (.A(net5449),
    .B(net6172),
    .CON(_01205_),
    .SN(_15729_));
 HAxp5_ASAP7_75t_R _30843_ (.A(net5448),
    .B(net6172),
    .CON(_01206_),
    .SN(_15730_));
 HAxp5_ASAP7_75t_R _30844_ (.A(net5448),
    .B(net6178),
    .CON(_01207_),
    .SN(_15731_));
 HAxp5_ASAP7_75t_R _30845_ (.A(_01674_),
    .B(_01636_),
    .CON(_01210_),
    .SN(_01211_));
 HAxp5_ASAP7_75t_R _30846_ (.A(net5742),
    .B(net5724),
    .CON(_01212_),
    .SN(_15732_));
 HAxp5_ASAP7_75t_R _30847_ (.A(_01599_),
    .B(net5742),
    .CON(_01214_),
    .SN(_15733_));
 HAxp5_ASAP7_75t_R _30848_ (.A(_01215_),
    .B(net5724),
    .CON(_01216_),
    .SN(_15734_));
 HAxp5_ASAP7_75t_R _30849_ (.A(_01215_),
    .B(net5724),
    .CON(_01217_),
    .SN(_15735_));
 HAxp5_ASAP7_75t_R _30850_ (.A(net5744),
    .B(net5745),
    .CON(_01218_),
    .SN(_15736_));
 HAxp5_ASAP7_75t_R _30851_ (.A(_01215_),
    .B(_01599_),
    .CON(_01219_),
    .SN(_15737_));
 HAxp5_ASAP7_75t_R _30852_ (.A(net5430),
    .B(net5724),
    .CON(_01221_),
    .SN(_01222_));
 HAxp5_ASAP7_75t_R _30853_ (.A(net5431),
    .B(net5747),
    .CON(_01223_),
    .SN(_15738_));
 HAxp5_ASAP7_75t_R _30854_ (.A(net5431),
    .B(net5747),
    .CON(_01224_),
    .SN(_15739_));
 HAxp5_ASAP7_75t_R _30855_ (.A(net5437),
    .B(net5724),
    .CON(_01226_),
    .SN(_15740_));
 HAxp5_ASAP7_75t_R _30856_ (.A(net5434),
    .B(net5724),
    .CON(_01227_),
    .SN(_15741_));
 HAxp5_ASAP7_75t_R _30857_ (.A(net5435),
    .B(net5747),
    .CON(_01228_),
    .SN(_15742_));
 HAxp5_ASAP7_75t_R _30858_ (.A(_01230_),
    .B(_02387_),
    .CON(_01231_),
    .SN(_01232_));
 HAxp5_ASAP7_75t_R _30859_ (.A(net5114),
    .B(net5711),
    .CON(_01233_),
    .SN(_15743_));
 HAxp5_ASAP7_75t_R _30860_ (.A(net5114),
    .B(_02297_),
    .CON(_01235_),
    .SN(_15744_));
 HAxp5_ASAP7_75t_R _30861_ (.A(_02297_),
    .B(net5114),
    .CON(_01236_),
    .SN(_15745_));
 HAxp5_ASAP7_75t_R _30862_ (.A(net5415),
    .B(net5711),
    .CON(_01238_),
    .SN(_15746_));
 HAxp5_ASAP7_75t_R _30863_ (.A(_01237_),
    .B(net5711),
    .CON(_01239_),
    .SN(_15747_));
 HAxp5_ASAP7_75t_R _30864_ (.A(_01237_),
    .B(_02297_),
    .CON(_01240_),
    .SN(_15748_));
 HAxp5_ASAP7_75t_R _30865_ (.A(_01237_),
    .B(_02297_),
    .CON(_01241_),
    .SN(_15749_));
 HAxp5_ASAP7_75t_R _30866_ (.A(net5412),
    .B(net5711),
    .CON(_01243_),
    .SN(_01244_));
 HAxp5_ASAP7_75t_R _30867_ (.A(net5412),
    .B(net5714),
    .CON(_01245_),
    .SN(_15750_));
 HAxp5_ASAP7_75t_R _30868_ (.A(net5412),
    .B(net5714),
    .CON(_01246_),
    .SN(_15751_));
 HAxp5_ASAP7_75t_R _30869_ (.A(net5413),
    .B(net5711),
    .CON(_01248_),
    .SN(_15752_));
 HAxp5_ASAP7_75t_R _30870_ (.A(net5413),
    .B(net5711),
    .CON(_01249_),
    .SN(_15753_));
 HAxp5_ASAP7_75t_R _30871_ (.A(_02336_),
    .B(net5714),
    .CON(_01250_),
    .SN(_15754_));
 HAxp5_ASAP7_75t_R _30872_ (.A(net5413),
    .B(net5714),
    .CON(_01251_),
    .SN(_15755_));
 HAxp5_ASAP7_75t_R _30873_ (.A(_01253_),
    .B(_03032_),
    .CON(_01254_),
    .SN(_01255_));
 HAxp5_ASAP7_75t_R _30874_ (.A(net5691),
    .B(net5395),
    .CON(_01256_),
    .SN(_15756_));
 HAxp5_ASAP7_75t_R _30875_ (.A(net5690),
    .B(net5403),
    .CON(_01258_),
    .SN(_15757_));
 HAxp5_ASAP7_75t_R _30876_ (.A(net5691),
    .B(_03011_),
    .CON(_01259_),
    .SN(_15758_));
 HAxp5_ASAP7_75t_R _30877_ (.A(net5695),
    .B(net5395),
    .CON(_01261_),
    .SN(_15759_));
 HAxp5_ASAP7_75t_R _30878_ (.A(_01260_),
    .B(net5395),
    .CON(_01262_),
    .SN(_15760_));
 HAxp5_ASAP7_75t_R _30879_ (.A(net5693),
    .B(net5403),
    .CON(_01263_),
    .SN(_15761_));
 HAxp5_ASAP7_75t_R _30880_ (.A(net5695),
    .B(net5403),
    .CON(_01264_),
    .SN(_15762_));
 HAxp5_ASAP7_75t_R _30881_ (.A(net5691),
    .B(net5396),
    .CON(_01266_),
    .SN(_01267_));
 HAxp5_ASAP7_75t_R _30882_ (.A(net5690),
    .B(net5400),
    .CON(_01269_),
    .SN(_15763_));
 HAxp5_ASAP7_75t_R _30883_ (.A(net5691),
    .B(net5399),
    .CON(_01270_),
    .SN(_15764_));
 HAxp5_ASAP7_75t_R _30884_ (.A(net5693),
    .B(net5396),
    .CON(_01271_),
    .SN(_15765_));
 HAxp5_ASAP7_75t_R _30885_ (.A(net5694),
    .B(net5398),
    .CON(_01272_),
    .SN(_15766_));
 HAxp5_ASAP7_75t_R _30886_ (.A(net5693),
    .B(net5399),
    .CON(_01273_),
    .SN(_15767_));
 HAxp5_ASAP7_75t_R _30887_ (.A(net5693),
    .B(net5399),
    .CON(_01274_),
    .SN(_15768_));
 HAxp5_ASAP7_75t_R _30888_ (.A(_03796_),
    .B(_01275_),
    .CON(_01277_),
    .SN(_01278_));
 HAxp5_ASAP7_75t_R _30889_ (.A(net5675),
    .B(net5384),
    .CON(_01279_),
    .SN(_15769_));
 HAxp5_ASAP7_75t_R _30890_ (.A(net5675),
    .B(_01280_),
    .CON(_01281_),
    .SN(_15770_));
 HAxp5_ASAP7_75t_R _30891_ (.A(net5675),
    .B(_01280_),
    .CON(_01282_),
    .SN(_15771_));
 HAxp5_ASAP7_75t_R _30892_ (.A(net5678),
    .B(net5384),
    .CON(_01284_),
    .SN(_15772_));
 HAxp5_ASAP7_75t_R _30893_ (.A(_01283_),
    .B(net5385),
    .CON(_01285_),
    .SN(_15773_));
 HAxp5_ASAP7_75t_R _30894_ (.A(net5678),
    .B(_01280_),
    .CON(_01286_),
    .SN(_15774_));
 HAxp5_ASAP7_75t_R _30895_ (.A(net5678),
    .B(_01280_),
    .CON(_01287_),
    .SN(_15775_));
 HAxp5_ASAP7_75t_R _30896_ (.A(net5675),
    .B(net5387),
    .CON(_01289_),
    .SN(_01290_));
 HAxp5_ASAP7_75t_R _30897_ (.A(net5675),
    .B(net5388),
    .CON(_01292_),
    .SN(_15776_));
 HAxp5_ASAP7_75t_R _30898_ (.A(net5675),
    .B(net5388),
    .CON(_01293_),
    .SN(_15777_));
 HAxp5_ASAP7_75t_R _30899_ (.A(net5677),
    .B(net5387),
    .CON(_01294_),
    .SN(_15778_));
 HAxp5_ASAP7_75t_R _30900_ (.A(net5677),
    .B(net5386),
    .CON(_01295_),
    .SN(_15779_));
 HAxp5_ASAP7_75t_R _30901_ (.A(net5677),
    .B(net5388),
    .CON(_01296_),
    .SN(_15780_));
 HAxp5_ASAP7_75t_R _30902_ (.A(net5677),
    .B(net5388),
    .CON(_01297_),
    .SN(_15781_));
 HAxp5_ASAP7_75t_R _30903_ (.A(_04500_),
    .B(_04431_),
    .CON(_01300_),
    .SN(_01301_));
 HAxp5_ASAP7_75t_R _30904_ (.A(net5663),
    .B(net5379),
    .CON(_01302_),
    .SN(_15782_));
 HAxp5_ASAP7_75t_R _30905_ (.A(net5663),
    .B(net5383),
    .CON(_01304_),
    .SN(_15783_));
 HAxp5_ASAP7_75t_R _30906_ (.A(net5663),
    .B(_01303_),
    .CON(_01305_),
    .SN(_15784_));
 HAxp5_ASAP7_75t_R _30907_ (.A(_01306_),
    .B(net5379),
    .CON(_01307_),
    .SN(_15785_));
 HAxp5_ASAP7_75t_R _30908_ (.A(_01306_),
    .B(net5379),
    .CON(_01308_),
    .SN(_15786_));
 HAxp5_ASAP7_75t_R _30909_ (.A(_01306_),
    .B(_01303_),
    .CON(_01309_),
    .SN(_15787_));
 HAxp5_ASAP7_75t_R _30910_ (.A(net5665),
    .B(_01303_),
    .CON(_01310_),
    .SN(_15788_));
 HAxp5_ASAP7_75t_R _30911_ (.A(net5663),
    .B(net5102),
    .CON(_01312_),
    .SN(_01313_));
 HAxp5_ASAP7_75t_R _30912_ (.A(net5663),
    .B(net5104),
    .CON(_01315_),
    .SN(_15789_));
 HAxp5_ASAP7_75t_R _30913_ (.A(net5663),
    .B(net5104),
    .CON(_01316_),
    .SN(_15790_));
 HAxp5_ASAP7_75t_R _30914_ (.A(net5666),
    .B(_04434_),
    .CON(_01317_),
    .SN(_15791_));
 HAxp5_ASAP7_75t_R _30915_ (.A(net5666),
    .B(net5102),
    .CON(_01318_),
    .SN(_15792_));
 HAxp5_ASAP7_75t_R _30916_ (.A(net5666),
    .B(net5103),
    .CON(_01319_),
    .SN(_15793_));
 HAxp5_ASAP7_75t_R _30917_ (.A(net5666),
    .B(net5103),
    .CON(_01320_),
    .SN(_15794_));
 HAxp5_ASAP7_75t_R _30918_ (.A(_05123_),
    .B(_01321_),
    .CON(_01323_),
    .SN(_01324_));
 HAxp5_ASAP7_75t_R _30919_ (.A(net5374),
    .B(net5096),
    .CON(_01325_),
    .SN(_15795_));
 HAxp5_ASAP7_75t_R _30920_ (.A(net5374),
    .B(net5098),
    .CON(_01327_),
    .SN(_15796_));
 HAxp5_ASAP7_75t_R _30921_ (.A(net5374),
    .B(_05103_),
    .CON(_01328_),
    .SN(_15797_));
 HAxp5_ASAP7_75t_R _30922_ (.A(net5096),
    .B(net5642),
    .CON(_01330_),
    .SN(_15798_));
 HAxp5_ASAP7_75t_R _30923_ (.A(net5641),
    .B(net5097),
    .CON(_01331_),
    .SN(_15799_));
 HAxp5_ASAP7_75t_R _30924_ (.A(net5642),
    .B(_05103_),
    .CON(_01332_),
    .SN(_15800_));
 HAxp5_ASAP7_75t_R _30925_ (.A(net5373),
    .B(net5636),
    .CON(_01334_),
    .SN(_01335_));
 HAxp5_ASAP7_75t_R _30926_ (.A(net5374),
    .B(net5639),
    .CON(_01337_),
    .SN(_15801_));
 HAxp5_ASAP7_75t_R _30927_ (.A(net5373),
    .B(net5638),
    .CON(_01338_),
    .SN(_15802_));
 HAxp5_ASAP7_75t_R _30928_ (.A(net5641),
    .B(net5637),
    .CON(_01339_),
    .SN(_15803_));
 HAxp5_ASAP7_75t_R _30929_ (.A(net5640),
    .B(net5636),
    .CON(_01340_),
    .SN(_15804_));
 HAxp5_ASAP7_75t_R _30930_ (.A(net5641),
    .B(net5638),
    .CON(_01341_),
    .SN(_15805_));
 HAxp5_ASAP7_75t_R _30931_ (.A(_05800_),
    .B(_05845_),
    .CON(_01344_),
    .SN(_01345_));
 HAxp5_ASAP7_75t_R _30932_ (.A(net5608),
    .B(net5619),
    .CON(_01346_),
    .SN(_15806_));
 HAxp5_ASAP7_75t_R _30933_ (.A(net5608),
    .B(_05777_),
    .CON(_01348_),
    .SN(_15807_));
 HAxp5_ASAP7_75t_R _30934_ (.A(net5608),
    .B(_05777_),
    .CON(_01349_),
    .SN(_15808_));
 HAxp5_ASAP7_75t_R _30935_ (.A(_05766_),
    .B(net5619),
    .CON(_01351_),
    .SN(_15809_));
 HAxp5_ASAP7_75t_R _30936_ (.A(net5628),
    .B(net5625),
    .CON(_01352_),
    .SN(_15810_));
 HAxp5_ASAP7_75t_R _30937_ (.A(net5629),
    .B(_05777_),
    .CON(_01353_),
    .SN(_15811_));
 HAxp5_ASAP7_75t_R _30938_ (.A(net5608),
    .B(net5616),
    .CON(_01355_),
    .SN(_01356_));
 HAxp5_ASAP7_75t_R _30939_ (.A(net5607),
    .B(net5623),
    .CON(_01358_),
    .SN(_15812_));
 HAxp5_ASAP7_75t_R _30940_ (.A(net5608),
    .B(net5623),
    .CON(_01359_),
    .SN(_15813_));
 HAxp5_ASAP7_75t_R _30941_ (.A(net5630),
    .B(net5616),
    .CON(_01360_),
    .SN(_15814_));
 HAxp5_ASAP7_75t_R _30942_ (.A(net5627),
    .B(net5616),
    .CON(_01361_),
    .SN(_15815_));
 HAxp5_ASAP7_75t_R _30943_ (.A(net5630),
    .B(net5620),
    .CON(_01362_),
    .SN(_15816_));
 HAxp5_ASAP7_75t_R _30944_ (.A(_06492_),
    .B(_06582_),
    .CON(_01365_),
    .SN(_01366_));
 HAxp5_ASAP7_75t_R _30945_ (.A(net5590),
    .B(net5081),
    .CON(_01367_),
    .SN(_15817_));
 HAxp5_ASAP7_75t_R _30946_ (.A(net5590),
    .B(_06472_),
    .CON(_01369_),
    .SN(_15818_));
 HAxp5_ASAP7_75t_R _30947_ (.A(net5590),
    .B(_06472_),
    .CON(_01370_),
    .SN(_15819_));
 HAxp5_ASAP7_75t_R _30948_ (.A(_06457_),
    .B(net5081),
    .CON(_01372_),
    .SN(_15820_));
 HAxp5_ASAP7_75t_R _30949_ (.A(net5603),
    .B(net5083),
    .CON(_01373_),
    .SN(_15821_));
 HAxp5_ASAP7_75t_R _30950_ (.A(_06457_),
    .B(_06472_),
    .CON(_01374_),
    .SN(_15822_));
 HAxp5_ASAP7_75t_R _30951_ (.A(net5590),
    .B(net5595),
    .CON(_01376_),
    .SN(_01377_));
 HAxp5_ASAP7_75t_R _30952_ (.A(net5590),
    .B(net5600),
    .CON(_01379_),
    .SN(_15823_));
 HAxp5_ASAP7_75t_R _30953_ (.A(net5590),
    .B(net5600),
    .CON(_01380_),
    .SN(_15824_));
 HAxp5_ASAP7_75t_R _30954_ (.A(net5602),
    .B(net5595),
    .CON(_01381_),
    .SN(_15825_));
 HAxp5_ASAP7_75t_R _30955_ (.A(net5602),
    .B(net5596),
    .CON(_01382_),
    .SN(_15826_));
 HAxp5_ASAP7_75t_R _30956_ (.A(net5602),
    .B(net5600),
    .CON(_01383_),
    .SN(_15827_));
 HAxp5_ASAP7_75t_R _30957_ (.A(_07136_),
    .B(_01384_),
    .CON(_01386_),
    .SN(_01387_));
 HAxp5_ASAP7_75t_R _30958_ (.A(net5575),
    .B(net5585),
    .CON(_01388_),
    .SN(_15828_));
 HAxp5_ASAP7_75t_R _30959_ (.A(net5575),
    .B(_01389_),
    .CON(_01390_),
    .SN(_15829_));
 HAxp5_ASAP7_75t_R _30960_ (.A(net5575),
    .B(_01389_),
    .CON(_01391_),
    .SN(_15830_));
 HAxp5_ASAP7_75t_R _30961_ (.A(_07123_),
    .B(net5585),
    .CON(_01393_),
    .SN(_15831_));
 HAxp5_ASAP7_75t_R _30962_ (.A(net5586),
    .B(net5337),
    .CON(_01394_),
    .SN(_15832_));
 HAxp5_ASAP7_75t_R _30963_ (.A(_07123_),
    .B(_01389_),
    .CON(_01395_),
    .SN(_15833_));
 HAxp5_ASAP7_75t_R _30964_ (.A(net5575),
    .B(net5576),
    .CON(_01397_),
    .SN(_01398_));
 HAxp5_ASAP7_75t_R _30965_ (.A(net5575),
    .B(net5581),
    .CON(_01400_),
    .SN(_15834_));
 HAxp5_ASAP7_75t_R _30966_ (.A(net5575),
    .B(net5582),
    .CON(_01401_),
    .SN(_15835_));
 HAxp5_ASAP7_75t_R _30967_ (.A(net5586),
    .B(net5576),
    .CON(_01402_),
    .SN(_15836_));
 HAxp5_ASAP7_75t_R _30968_ (.A(net5586),
    .B(net5576),
    .CON(_01403_),
    .SN(_15837_));
 HAxp5_ASAP7_75t_R _30969_ (.A(net5586),
    .B(net5582),
    .CON(_01404_),
    .SN(_15838_));
 BUFx16f_ASAP7_75t_R clkbuf_0_clk (.A(clk),
    .Y(clknet_0_clk));
 BUFx24_ASAP7_75t_R clkbuf_2_0_0_clk (.A(clknet_0_clk),
    .Y(clknet_2_0_0_clk));
 BUFx24_ASAP7_75t_R clkbuf_2_1_0_clk (.A(clknet_0_clk),
    .Y(clknet_2_1_0_clk));
 BUFx24_ASAP7_75t_R clkbuf_2_2_0_clk (.A(clknet_0_clk),
    .Y(clknet_2_2_0_clk));
 BUFx24_ASAP7_75t_R clkbuf_2_3_0_clk (.A(clknet_0_clk),
    .Y(clknet_2_3_0_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_0_clk (.A(clknet_2_0_0_clk),
    .Y(clknet_leaf_0_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_10_clk (.A(clknet_2_1_0_clk),
    .Y(clknet_leaf_10_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_11_clk (.A(clknet_2_3_0_clk),
    .Y(clknet_leaf_11_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_12_clk (.A(clknet_2_3_0_clk),
    .Y(clknet_leaf_12_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_13_clk (.A(clknet_2_3_0_clk),
    .Y(clknet_leaf_13_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_14_clk (.A(clknet_2_3_0_clk),
    .Y(clknet_leaf_14_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_15_clk (.A(clknet_2_3_0_clk),
    .Y(clknet_leaf_15_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_16_clk (.A(clknet_2_3_0_clk),
    .Y(clknet_leaf_16_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_17_clk (.A(clknet_2_3_0_clk),
    .Y(clknet_leaf_17_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_18_clk (.A(clknet_2_3_0_clk),
    .Y(clknet_leaf_18_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_19_clk (.A(clknet_2_3_0_clk),
    .Y(clknet_leaf_19_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_1_clk (.A(clknet_2_0_0_clk),
    .Y(clknet_leaf_1_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_20_clk (.A(clknet_2_2_0_clk),
    .Y(clknet_leaf_20_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_21_clk (.A(clknet_2_2_0_clk),
    .Y(clknet_leaf_21_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_22_clk (.A(clknet_2_2_0_clk),
    .Y(clknet_leaf_22_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_23_clk (.A(clknet_2_2_0_clk),
    .Y(clknet_leaf_23_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_24_clk (.A(clknet_2_2_0_clk),
    .Y(clknet_leaf_24_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_25_clk (.A(clknet_2_2_0_clk),
    .Y(clknet_leaf_25_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_26_clk (.A(clknet_2_2_0_clk),
    .Y(clknet_leaf_26_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_27_clk (.A(clknet_2_2_0_clk),
    .Y(clknet_leaf_27_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_28_clk (.A(clknet_2_2_0_clk),
    .Y(clknet_leaf_28_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_29_clk (.A(clknet_2_0_0_clk),
    .Y(clknet_leaf_29_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_2_clk (.A(clknet_2_1_0_clk),
    .Y(clknet_leaf_2_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_30_clk (.A(clknet_2_0_0_clk),
    .Y(clknet_leaf_30_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_31_clk (.A(clknet_2_0_0_clk),
    .Y(clknet_leaf_31_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_32_clk (.A(clknet_2_0_0_clk),
    .Y(clknet_leaf_32_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_33_clk (.A(clknet_2_0_0_clk),
    .Y(clknet_leaf_33_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_34_clk (.A(clknet_2_0_0_clk),
    .Y(clknet_leaf_34_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_3_clk (.A(clknet_2_1_0_clk),
    .Y(clknet_leaf_3_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_4_clk (.A(clknet_2_1_0_clk),
    .Y(clknet_leaf_4_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_5_clk (.A(clknet_2_1_0_clk),
    .Y(clknet_leaf_5_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_6_clk (.A(clknet_2_1_0_clk),
    .Y(clknet_leaf_6_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_7_clk (.A(clknet_2_1_0_clk),
    .Y(clknet_leaf_7_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_8_clk (.A(clknet_2_1_0_clk),
    .Y(clknet_leaf_8_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_9_clk (.A(clknet_2_1_0_clk),
    .Y(clknet_leaf_9_clk));
 BUFx24_ASAP7_75t_R clkload0 (.A(clknet_2_0_0_clk));
 CKINVDCx6p67_ASAP7_75t_R clkload1 (.A(clknet_leaf_0_clk));
 BUFx24_ASAP7_75t_R clkload10 (.A(clknet_leaf_5_clk));
 BUFx2_ASAP7_75t_R clkload11 (.A(clknet_leaf_6_clk));
 CKINVDCx8_ASAP7_75t_R clkload12 (.A(clknet_leaf_7_clk));
 INVx6_ASAP7_75t_R clkload13 (.A(clknet_leaf_8_clk));
 CKINVDCx5p33_ASAP7_75t_R clkload14 (.A(clknet_leaf_9_clk));
 CKINVDCx6p67_ASAP7_75t_R clkload15 (.A(clknet_leaf_10_clk));
 BUFx24_ASAP7_75t_R clkload16 (.A(clknet_leaf_20_clk));
 INVx5_ASAP7_75t_R clkload17 (.A(clknet_leaf_21_clk));
 INVx6_ASAP7_75t_R clkload18 (.A(clknet_leaf_22_clk));
 BUFx24_ASAP7_75t_R clkload19 (.A(clknet_leaf_23_clk));
 INVx3_ASAP7_75t_R clkload2 (.A(clknet_leaf_1_clk));
 CKINVDCx9p33_ASAP7_75t_R clkload20 (.A(clknet_leaf_25_clk));
 CKINVDCx9p33_ASAP7_75t_R clkload21 (.A(clknet_leaf_26_clk));
 CKINVDCx5p33_ASAP7_75t_R clkload22 (.A(clknet_leaf_27_clk));
 CKINVDCx8_ASAP7_75t_R clkload23 (.A(clknet_leaf_28_clk));
 BUFx24_ASAP7_75t_R clkload24 (.A(clknet_leaf_11_clk));
 CKINVDCx5p33_ASAP7_75t_R clkload25 (.A(clknet_leaf_12_clk));
 BUFx12_ASAP7_75t_R clkload26 (.A(clknet_leaf_13_clk));
 BUFx12_ASAP7_75t_R clkload27 (.A(clknet_leaf_14_clk));
 INVx8_ASAP7_75t_R clkload28 (.A(clknet_leaf_15_clk));
 INVx5_ASAP7_75t_R clkload29 (.A(clknet_leaf_17_clk));
 BUFx24_ASAP7_75t_R clkload3 (.A(clknet_leaf_29_clk));
 CKINVDCx5p33_ASAP7_75t_R clkload30 (.A(clknet_leaf_18_clk));
 INVx5_ASAP7_75t_R clkload31 (.A(clknet_leaf_19_clk));
 INVx6_ASAP7_75t_R clkload4 (.A(clknet_leaf_30_clk));
 INVx6_ASAP7_75t_R clkload5 (.A(clknet_leaf_32_clk));
 INVx3_ASAP7_75t_R clkload6 (.A(clknet_leaf_33_clk));
 CKINVDCx10_ASAP7_75t_R clkload7 (.A(clknet_leaf_34_clk));
 CKINVDCx6p67_ASAP7_75t_R clkload8 (.A(clknet_leaf_2_clk));
 BUFx4f_ASAP7_75t_R clkload9 (.A(clknet_leaf_4_clk));
 DFFHQNx1_ASAP7_75t_R \dcnt[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .D(_01405_),
    .QN(_00572_));
 DFFHQNx1_ASAP7_75t_R \dcnt[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .D(_01406_),
    .QN(_00571_));
 DFFHQNx1_ASAP7_75t_R \dcnt[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_32_clk),
    .D(_01407_),
    .QN(_00570_));
 DFFHQNx1_ASAP7_75t_R \dcnt[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .D(_01408_),
    .QN(_00411_));
 DFFHQNx1_ASAP7_75t_R \done$_DFF_P_  (.CLK(clknet_leaf_32_clk),
    .D(_00160_),
    .QN(_00573_));
 BUFx2_ASAP7_75t_R input1 (.A(key[0]),
    .Y(net1));
 BUFx2_ASAP7_75t_R input10 (.A(key[108]),
    .Y(net10));
 BUFx2_ASAP7_75t_R input100 (.A(key[74]),
    .Y(net100));
 BUFx2_ASAP7_75t_R input101 (.A(key[75]),
    .Y(net101));
 BUFx2_ASAP7_75t_R input102 (.A(key[76]),
    .Y(net102));
 BUFx2_ASAP7_75t_R input103 (.A(key[77]),
    .Y(net103));
 BUFx2_ASAP7_75t_R input104 (.A(key[78]),
    .Y(net104));
 BUFx2_ASAP7_75t_R input105 (.A(key[79]),
    .Y(net105));
 BUFx2_ASAP7_75t_R input106 (.A(key[7]),
    .Y(net106));
 BUFx2_ASAP7_75t_R input107 (.A(key[80]),
    .Y(net107));
 BUFx2_ASAP7_75t_R input108 (.A(key[81]),
    .Y(net108));
 BUFx2_ASAP7_75t_R input109 (.A(key[82]),
    .Y(net109));
 BUFx2_ASAP7_75t_R input11 (.A(key[109]),
    .Y(net11));
 BUFx2_ASAP7_75t_R input110 (.A(key[83]),
    .Y(net110));
 BUFx2_ASAP7_75t_R input111 (.A(key[84]),
    .Y(net111));
 BUFx2_ASAP7_75t_R input112 (.A(key[85]),
    .Y(net112));
 BUFx2_ASAP7_75t_R input113 (.A(key[86]),
    .Y(net113));
 BUFx2_ASAP7_75t_R input114 (.A(key[87]),
    .Y(net114));
 BUFx2_ASAP7_75t_R input115 (.A(key[88]),
    .Y(net115));
 BUFx2_ASAP7_75t_R input116 (.A(key[89]),
    .Y(net116));
 BUFx2_ASAP7_75t_R input117 (.A(key[8]),
    .Y(net117));
 BUFx2_ASAP7_75t_R input118 (.A(key[90]),
    .Y(net118));
 BUFx2_ASAP7_75t_R input119 (.A(key[91]),
    .Y(net119));
 BUFx2_ASAP7_75t_R input12 (.A(key[10]),
    .Y(net12));
 BUFx2_ASAP7_75t_R input120 (.A(key[92]),
    .Y(net120));
 BUFx2_ASAP7_75t_R input121 (.A(key[93]),
    .Y(net121));
 BUFx2_ASAP7_75t_R input122 (.A(key[94]),
    .Y(net122));
 BUFx2_ASAP7_75t_R input123 (.A(key[95]),
    .Y(net123));
 BUFx2_ASAP7_75t_R input124 (.A(key[96]),
    .Y(net124));
 BUFx2_ASAP7_75t_R input125 (.A(key[97]),
    .Y(net125));
 BUFx2_ASAP7_75t_R input126 (.A(key[98]),
    .Y(net126));
 BUFx2_ASAP7_75t_R input127 (.A(key[99]),
    .Y(net127));
 BUFx2_ASAP7_75t_R input128 (.A(key[9]),
    .Y(net128));
 BUFx8_ASAP7_75t_R input129 (.A(ld),
    .Y(net129));
 BUFx2_ASAP7_75t_R input13 (.A(key[110]),
    .Y(net13));
 BUFx2_ASAP7_75t_R input130 (.A(rst),
    .Y(net130));
 BUFx2_ASAP7_75t_R input131 (.A(text_in[0]),
    .Y(net131));
 BUFx2_ASAP7_75t_R input132 (.A(text_in[100]),
    .Y(net132));
 BUFx2_ASAP7_75t_R input133 (.A(text_in[101]),
    .Y(net133));
 BUFx2_ASAP7_75t_R input134 (.A(text_in[102]),
    .Y(net134));
 BUFx2_ASAP7_75t_R input135 (.A(text_in[103]),
    .Y(net135));
 BUFx2_ASAP7_75t_R input136 (.A(text_in[104]),
    .Y(net136));
 BUFx2_ASAP7_75t_R input137 (.A(text_in[105]),
    .Y(net137));
 BUFx2_ASAP7_75t_R input138 (.A(text_in[106]),
    .Y(net138));
 BUFx2_ASAP7_75t_R input139 (.A(text_in[107]),
    .Y(net139));
 BUFx2_ASAP7_75t_R input14 (.A(key[111]),
    .Y(net14));
 BUFx2_ASAP7_75t_R input140 (.A(text_in[108]),
    .Y(net140));
 BUFx2_ASAP7_75t_R input141 (.A(text_in[109]),
    .Y(net141));
 BUFx2_ASAP7_75t_R input142 (.A(text_in[10]),
    .Y(net142));
 BUFx2_ASAP7_75t_R input143 (.A(text_in[110]),
    .Y(net143));
 BUFx2_ASAP7_75t_R input144 (.A(text_in[111]),
    .Y(net144));
 BUFx2_ASAP7_75t_R input145 (.A(text_in[112]),
    .Y(net145));
 BUFx2_ASAP7_75t_R input146 (.A(text_in[113]),
    .Y(net146));
 BUFx2_ASAP7_75t_R input147 (.A(text_in[114]),
    .Y(net147));
 BUFx2_ASAP7_75t_R input148 (.A(text_in[115]),
    .Y(net148));
 BUFx2_ASAP7_75t_R input149 (.A(text_in[116]),
    .Y(net149));
 BUFx2_ASAP7_75t_R input15 (.A(key[112]),
    .Y(net15));
 BUFx2_ASAP7_75t_R input150 (.A(text_in[117]),
    .Y(net150));
 BUFx2_ASAP7_75t_R input151 (.A(text_in[118]),
    .Y(net151));
 BUFx2_ASAP7_75t_R input152 (.A(text_in[119]),
    .Y(net152));
 BUFx2_ASAP7_75t_R input153 (.A(text_in[11]),
    .Y(net153));
 BUFx2_ASAP7_75t_R input154 (.A(text_in[120]),
    .Y(net154));
 BUFx2_ASAP7_75t_R input155 (.A(text_in[121]),
    .Y(net155));
 BUFx2_ASAP7_75t_R input156 (.A(text_in[122]),
    .Y(net156));
 BUFx2_ASAP7_75t_R input157 (.A(text_in[123]),
    .Y(net157));
 BUFx2_ASAP7_75t_R input158 (.A(text_in[124]),
    .Y(net158));
 BUFx2_ASAP7_75t_R input159 (.A(text_in[125]),
    .Y(net159));
 BUFx2_ASAP7_75t_R input16 (.A(key[113]),
    .Y(net16));
 BUFx2_ASAP7_75t_R input160 (.A(text_in[126]),
    .Y(net160));
 BUFx2_ASAP7_75t_R input161 (.A(text_in[127]),
    .Y(net161));
 BUFx2_ASAP7_75t_R input162 (.A(text_in[12]),
    .Y(net162));
 BUFx2_ASAP7_75t_R input163 (.A(text_in[13]),
    .Y(net163));
 BUFx2_ASAP7_75t_R input164 (.A(text_in[14]),
    .Y(net164));
 BUFx2_ASAP7_75t_R input165 (.A(text_in[15]),
    .Y(net165));
 BUFx2_ASAP7_75t_R input166 (.A(text_in[16]),
    .Y(net166));
 BUFx2_ASAP7_75t_R input167 (.A(text_in[17]),
    .Y(net167));
 BUFx2_ASAP7_75t_R input168 (.A(text_in[18]),
    .Y(net168));
 BUFx2_ASAP7_75t_R input169 (.A(text_in[19]),
    .Y(net169));
 BUFx2_ASAP7_75t_R input17 (.A(key[114]),
    .Y(net17));
 BUFx2_ASAP7_75t_R input170 (.A(text_in[1]),
    .Y(net170));
 BUFx2_ASAP7_75t_R input171 (.A(text_in[20]),
    .Y(net171));
 BUFx2_ASAP7_75t_R input172 (.A(text_in[21]),
    .Y(net172));
 BUFx2_ASAP7_75t_R input173 (.A(text_in[22]),
    .Y(net173));
 BUFx2_ASAP7_75t_R input174 (.A(text_in[23]),
    .Y(net174));
 BUFx2_ASAP7_75t_R input175 (.A(text_in[24]),
    .Y(net175));
 BUFx2_ASAP7_75t_R input176 (.A(text_in[25]),
    .Y(net176));
 BUFx2_ASAP7_75t_R input177 (.A(text_in[26]),
    .Y(net177));
 BUFx2_ASAP7_75t_R input178 (.A(text_in[27]),
    .Y(net178));
 BUFx2_ASAP7_75t_R input179 (.A(text_in[28]),
    .Y(net179));
 BUFx2_ASAP7_75t_R input18 (.A(key[115]),
    .Y(net18));
 BUFx2_ASAP7_75t_R input180 (.A(text_in[29]),
    .Y(net180));
 BUFx2_ASAP7_75t_R input181 (.A(text_in[2]),
    .Y(net181));
 BUFx2_ASAP7_75t_R input182 (.A(text_in[30]),
    .Y(net182));
 BUFx2_ASAP7_75t_R input183 (.A(text_in[31]),
    .Y(net183));
 BUFx2_ASAP7_75t_R input184 (.A(text_in[32]),
    .Y(net184));
 BUFx2_ASAP7_75t_R input185 (.A(text_in[33]),
    .Y(net185));
 BUFx2_ASAP7_75t_R input186 (.A(text_in[34]),
    .Y(net186));
 BUFx2_ASAP7_75t_R input187 (.A(text_in[35]),
    .Y(net187));
 BUFx2_ASAP7_75t_R input188 (.A(text_in[36]),
    .Y(net188));
 BUFx2_ASAP7_75t_R input189 (.A(text_in[37]),
    .Y(net189));
 BUFx2_ASAP7_75t_R input19 (.A(key[116]),
    .Y(net19));
 BUFx2_ASAP7_75t_R input190 (.A(text_in[38]),
    .Y(net190));
 BUFx2_ASAP7_75t_R input191 (.A(text_in[39]),
    .Y(net191));
 BUFx2_ASAP7_75t_R input192 (.A(text_in[3]),
    .Y(net192));
 BUFx2_ASAP7_75t_R input193 (.A(text_in[40]),
    .Y(net193));
 BUFx2_ASAP7_75t_R input194 (.A(text_in[41]),
    .Y(net194));
 BUFx2_ASAP7_75t_R input195 (.A(text_in[42]),
    .Y(net195));
 BUFx2_ASAP7_75t_R input196 (.A(text_in[43]),
    .Y(net196));
 BUFx2_ASAP7_75t_R input197 (.A(text_in[44]),
    .Y(net197));
 BUFx2_ASAP7_75t_R input198 (.A(text_in[45]),
    .Y(net198));
 BUFx2_ASAP7_75t_R input199 (.A(text_in[46]),
    .Y(net199));
 BUFx2_ASAP7_75t_R input2 (.A(key[100]),
    .Y(net2));
 BUFx2_ASAP7_75t_R input20 (.A(key[117]),
    .Y(net20));
 BUFx2_ASAP7_75t_R input200 (.A(text_in[47]),
    .Y(net200));
 BUFx2_ASAP7_75t_R input201 (.A(text_in[48]),
    .Y(net201));
 BUFx2_ASAP7_75t_R input202 (.A(text_in[49]),
    .Y(net202));
 BUFx2_ASAP7_75t_R input203 (.A(text_in[4]),
    .Y(net203));
 BUFx2_ASAP7_75t_R input204 (.A(text_in[50]),
    .Y(net204));
 BUFx2_ASAP7_75t_R input205 (.A(text_in[51]),
    .Y(net205));
 BUFx2_ASAP7_75t_R input206 (.A(text_in[52]),
    .Y(net206));
 BUFx2_ASAP7_75t_R input207 (.A(text_in[53]),
    .Y(net207));
 BUFx2_ASAP7_75t_R input208 (.A(text_in[54]),
    .Y(net208));
 BUFx2_ASAP7_75t_R input209 (.A(text_in[55]),
    .Y(net209));
 BUFx2_ASAP7_75t_R input21 (.A(key[118]),
    .Y(net21));
 BUFx2_ASAP7_75t_R input210 (.A(text_in[56]),
    .Y(net210));
 BUFx2_ASAP7_75t_R input211 (.A(text_in[57]),
    .Y(net211));
 BUFx2_ASAP7_75t_R input212 (.A(text_in[58]),
    .Y(net212));
 BUFx2_ASAP7_75t_R input213 (.A(text_in[59]),
    .Y(net213));
 BUFx2_ASAP7_75t_R input214 (.A(text_in[5]),
    .Y(net214));
 BUFx2_ASAP7_75t_R input215 (.A(text_in[60]),
    .Y(net215));
 BUFx2_ASAP7_75t_R input216 (.A(text_in[61]),
    .Y(net216));
 BUFx2_ASAP7_75t_R input217 (.A(text_in[62]),
    .Y(net217));
 BUFx2_ASAP7_75t_R input218 (.A(text_in[63]),
    .Y(net218));
 BUFx2_ASAP7_75t_R input219 (.A(text_in[64]),
    .Y(net219));
 BUFx2_ASAP7_75t_R input22 (.A(key[119]),
    .Y(net22));
 BUFx2_ASAP7_75t_R input220 (.A(text_in[65]),
    .Y(net220));
 BUFx2_ASAP7_75t_R input221 (.A(text_in[66]),
    .Y(net221));
 BUFx2_ASAP7_75t_R input222 (.A(text_in[67]),
    .Y(net222));
 BUFx2_ASAP7_75t_R input223 (.A(text_in[68]),
    .Y(net223));
 BUFx2_ASAP7_75t_R input224 (.A(text_in[69]),
    .Y(net224));
 BUFx2_ASAP7_75t_R input225 (.A(text_in[6]),
    .Y(net225));
 BUFx2_ASAP7_75t_R input226 (.A(text_in[70]),
    .Y(net226));
 BUFx2_ASAP7_75t_R input227 (.A(text_in[71]),
    .Y(net227));
 BUFx2_ASAP7_75t_R input228 (.A(text_in[72]),
    .Y(net228));
 BUFx2_ASAP7_75t_R input229 (.A(text_in[73]),
    .Y(net229));
 BUFx2_ASAP7_75t_R input23 (.A(key[11]),
    .Y(net23));
 BUFx2_ASAP7_75t_R input230 (.A(text_in[74]),
    .Y(net230));
 BUFx2_ASAP7_75t_R input231 (.A(text_in[75]),
    .Y(net231));
 BUFx2_ASAP7_75t_R input232 (.A(text_in[76]),
    .Y(net232));
 BUFx2_ASAP7_75t_R input233 (.A(text_in[77]),
    .Y(net233));
 BUFx2_ASAP7_75t_R input234 (.A(text_in[78]),
    .Y(net234));
 BUFx2_ASAP7_75t_R input235 (.A(text_in[79]),
    .Y(net235));
 BUFx2_ASAP7_75t_R input236 (.A(text_in[7]),
    .Y(net236));
 BUFx2_ASAP7_75t_R input237 (.A(text_in[80]),
    .Y(net237));
 BUFx2_ASAP7_75t_R input238 (.A(text_in[81]),
    .Y(net238));
 BUFx2_ASAP7_75t_R input239 (.A(text_in[82]),
    .Y(net239));
 BUFx2_ASAP7_75t_R input24 (.A(key[120]),
    .Y(net24));
 BUFx2_ASAP7_75t_R input240 (.A(text_in[83]),
    .Y(net240));
 BUFx2_ASAP7_75t_R input241 (.A(text_in[84]),
    .Y(net241));
 BUFx2_ASAP7_75t_R input242 (.A(text_in[85]),
    .Y(net242));
 BUFx2_ASAP7_75t_R input243 (.A(text_in[86]),
    .Y(net243));
 BUFx2_ASAP7_75t_R input244 (.A(text_in[87]),
    .Y(net244));
 BUFx2_ASAP7_75t_R input245 (.A(text_in[88]),
    .Y(net245));
 BUFx2_ASAP7_75t_R input246 (.A(text_in[89]),
    .Y(net246));
 BUFx2_ASAP7_75t_R input247 (.A(text_in[8]),
    .Y(net247));
 BUFx2_ASAP7_75t_R input248 (.A(text_in[90]),
    .Y(net248));
 BUFx2_ASAP7_75t_R input249 (.A(text_in[91]),
    .Y(net249));
 BUFx2_ASAP7_75t_R input25 (.A(key[121]),
    .Y(net25));
 BUFx2_ASAP7_75t_R input250 (.A(text_in[92]),
    .Y(net250));
 BUFx2_ASAP7_75t_R input251 (.A(text_in[93]),
    .Y(net251));
 BUFx2_ASAP7_75t_R input252 (.A(text_in[94]),
    .Y(net252));
 BUFx2_ASAP7_75t_R input253 (.A(text_in[95]),
    .Y(net253));
 BUFx2_ASAP7_75t_R input254 (.A(text_in[96]),
    .Y(net254));
 BUFx2_ASAP7_75t_R input255 (.A(text_in[97]),
    .Y(net255));
 BUFx2_ASAP7_75t_R input256 (.A(text_in[98]),
    .Y(net256));
 BUFx2_ASAP7_75t_R input257 (.A(text_in[99]),
    .Y(net257));
 BUFx2_ASAP7_75t_R input258 (.A(text_in[9]),
    .Y(net258));
 BUFx2_ASAP7_75t_R input26 (.A(key[122]),
    .Y(net26));
 BUFx2_ASAP7_75t_R input27 (.A(key[123]),
    .Y(net27));
 BUFx2_ASAP7_75t_R input28 (.A(key[124]),
    .Y(net28));
 BUFx2_ASAP7_75t_R input29 (.A(key[125]),
    .Y(net29));
 BUFx2_ASAP7_75t_R input3 (.A(key[101]),
    .Y(net3));
 BUFx2_ASAP7_75t_R input30 (.A(key[126]),
    .Y(net30));
 BUFx2_ASAP7_75t_R input31 (.A(key[127]),
    .Y(net31));
 BUFx2_ASAP7_75t_R input32 (.A(key[12]),
    .Y(net32));
 BUFx2_ASAP7_75t_R input33 (.A(key[13]),
    .Y(net33));
 BUFx2_ASAP7_75t_R input34 (.A(key[14]),
    .Y(net34));
 BUFx2_ASAP7_75t_R input35 (.A(key[15]),
    .Y(net35));
 BUFx2_ASAP7_75t_R input36 (.A(key[16]),
    .Y(net36));
 BUFx2_ASAP7_75t_R input37 (.A(key[17]),
    .Y(net37));
 BUFx2_ASAP7_75t_R input38 (.A(key[18]),
    .Y(net38));
 BUFx2_ASAP7_75t_R input39 (.A(key[19]),
    .Y(net39));
 BUFx2_ASAP7_75t_R input4 (.A(key[102]),
    .Y(net4));
 BUFx2_ASAP7_75t_R input40 (.A(key[1]),
    .Y(net40));
 BUFx2_ASAP7_75t_R input41 (.A(key[20]),
    .Y(net41));
 BUFx2_ASAP7_75t_R input42 (.A(key[21]),
    .Y(net42));
 BUFx2_ASAP7_75t_R input43 (.A(key[22]),
    .Y(net43));
 BUFx2_ASAP7_75t_R input44 (.A(key[23]),
    .Y(net44));
 BUFx2_ASAP7_75t_R input45 (.A(key[24]),
    .Y(net45));
 BUFx2_ASAP7_75t_R input46 (.A(key[25]),
    .Y(net46));
 BUFx2_ASAP7_75t_R input47 (.A(key[26]),
    .Y(net47));
 BUFx2_ASAP7_75t_R input48 (.A(key[27]),
    .Y(net48));
 BUFx2_ASAP7_75t_R input49 (.A(key[28]),
    .Y(net49));
 BUFx2_ASAP7_75t_R input5 (.A(key[103]),
    .Y(net5));
 BUFx2_ASAP7_75t_R input50 (.A(key[29]),
    .Y(net50));
 BUFx2_ASAP7_75t_R input51 (.A(key[2]),
    .Y(net51));
 BUFx2_ASAP7_75t_R input52 (.A(key[30]),
    .Y(net52));
 BUFx2_ASAP7_75t_R input53 (.A(key[31]),
    .Y(net53));
 BUFx2_ASAP7_75t_R input54 (.A(key[32]),
    .Y(net54));
 BUFx2_ASAP7_75t_R input55 (.A(key[33]),
    .Y(net55));
 BUFx2_ASAP7_75t_R input56 (.A(key[34]),
    .Y(net56));
 BUFx2_ASAP7_75t_R input57 (.A(key[35]),
    .Y(net57));
 BUFx2_ASAP7_75t_R input58 (.A(key[36]),
    .Y(net58));
 BUFx2_ASAP7_75t_R input59 (.A(key[37]),
    .Y(net59));
 BUFx2_ASAP7_75t_R input6 (.A(key[104]),
    .Y(net6));
 BUFx2_ASAP7_75t_R input60 (.A(key[38]),
    .Y(net60));
 BUFx2_ASAP7_75t_R input61 (.A(key[39]),
    .Y(net61));
 BUFx2_ASAP7_75t_R input62 (.A(key[3]),
    .Y(net62));
 BUFx2_ASAP7_75t_R input63 (.A(key[40]),
    .Y(net63));
 BUFx2_ASAP7_75t_R input64 (.A(key[41]),
    .Y(net64));
 BUFx2_ASAP7_75t_R input65 (.A(key[42]),
    .Y(net65));
 BUFx2_ASAP7_75t_R input66 (.A(key[43]),
    .Y(net66));
 BUFx2_ASAP7_75t_R input67 (.A(key[44]),
    .Y(net67));
 BUFx2_ASAP7_75t_R input68 (.A(key[45]),
    .Y(net68));
 BUFx2_ASAP7_75t_R input69 (.A(key[46]),
    .Y(net69));
 BUFx2_ASAP7_75t_R input7 (.A(key[105]),
    .Y(net7));
 BUFx2_ASAP7_75t_R input70 (.A(key[47]),
    .Y(net70));
 BUFx2_ASAP7_75t_R input71 (.A(key[48]),
    .Y(net71));
 BUFx2_ASAP7_75t_R input72 (.A(key[49]),
    .Y(net72));
 BUFx2_ASAP7_75t_R input73 (.A(key[4]),
    .Y(net73));
 BUFx2_ASAP7_75t_R input74 (.A(key[50]),
    .Y(net74));
 BUFx2_ASAP7_75t_R input75 (.A(key[51]),
    .Y(net75));
 BUFx2_ASAP7_75t_R input76 (.A(key[52]),
    .Y(net76));
 BUFx2_ASAP7_75t_R input77 (.A(key[53]),
    .Y(net77));
 BUFx2_ASAP7_75t_R input78 (.A(key[54]),
    .Y(net78));
 BUFx2_ASAP7_75t_R input79 (.A(key[55]),
    .Y(net79));
 BUFx2_ASAP7_75t_R input8 (.A(key[106]),
    .Y(net8));
 BUFx2_ASAP7_75t_R input80 (.A(key[56]),
    .Y(net80));
 BUFx2_ASAP7_75t_R input81 (.A(key[57]),
    .Y(net81));
 BUFx2_ASAP7_75t_R input82 (.A(key[58]),
    .Y(net82));
 BUFx2_ASAP7_75t_R input83 (.A(key[59]),
    .Y(net83));
 BUFx2_ASAP7_75t_R input84 (.A(key[5]),
    .Y(net84));
 BUFx2_ASAP7_75t_R input85 (.A(key[60]),
    .Y(net85));
 BUFx2_ASAP7_75t_R input86 (.A(key[61]),
    .Y(net86));
 BUFx2_ASAP7_75t_R input87 (.A(key[62]),
    .Y(net87));
 BUFx2_ASAP7_75t_R input88 (.A(key[63]),
    .Y(net88));
 BUFx2_ASAP7_75t_R input89 (.A(key[64]),
    .Y(net89));
 BUFx2_ASAP7_75t_R input9 (.A(key[107]),
    .Y(net9));
 BUFx2_ASAP7_75t_R input90 (.A(key[65]),
    .Y(net90));
 BUFx2_ASAP7_75t_R input91 (.A(key[66]),
    .Y(net91));
 BUFx2_ASAP7_75t_R input92 (.A(key[67]),
    .Y(net92));
 BUFx2_ASAP7_75t_R input93 (.A(key[68]),
    .Y(net93));
 BUFx2_ASAP7_75t_R input94 (.A(key[69]),
    .Y(net94));
 BUFx2_ASAP7_75t_R input95 (.A(key[6]),
    .Y(net95));
 BUFx2_ASAP7_75t_R input96 (.A(key[70]),
    .Y(net96));
 BUFx2_ASAP7_75t_R input97 (.A(key[71]),
    .Y(net97));
 BUFx2_ASAP7_75t_R input98 (.A(key[72]),
    .Y(net98));
 BUFx2_ASAP7_75t_R input99 (.A(key[73]),
    .Y(net99));
 DFFHQNx3_ASAP7_75t_R \ld_r$_DFF_P_  (.CLK(clknet_leaf_19_clk),
    .D(net6683),
    .QN(_00574_));
 BUFx2_ASAP7_75t_R output259 (.A(net259),
    .Y(done));
 BUFx2_ASAP7_75t_R output260 (.A(net260),
    .Y(text_out[0]));
 BUFx2_ASAP7_75t_R output261 (.A(net261),
    .Y(text_out[100]));
 BUFx2_ASAP7_75t_R output262 (.A(net262),
    .Y(text_out[101]));
 BUFx2_ASAP7_75t_R output263 (.A(net263),
    .Y(text_out[102]));
 BUFx2_ASAP7_75t_R output264 (.A(net264),
    .Y(text_out[103]));
 BUFx2_ASAP7_75t_R output265 (.A(net265),
    .Y(text_out[104]));
 BUFx2_ASAP7_75t_R output266 (.A(net266),
    .Y(text_out[105]));
 BUFx2_ASAP7_75t_R output267 (.A(net267),
    .Y(text_out[106]));
 BUFx2_ASAP7_75t_R output268 (.A(net268),
    .Y(text_out[107]));
 BUFx2_ASAP7_75t_R output269 (.A(net269),
    .Y(text_out[108]));
 BUFx2_ASAP7_75t_R output270 (.A(net270),
    .Y(text_out[109]));
 BUFx2_ASAP7_75t_R output271 (.A(net271),
    .Y(text_out[10]));
 BUFx2_ASAP7_75t_R output272 (.A(net272),
    .Y(text_out[110]));
 BUFx2_ASAP7_75t_R output273 (.A(net273),
    .Y(text_out[111]));
 BUFx2_ASAP7_75t_R output274 (.A(net274),
    .Y(text_out[112]));
 BUFx2_ASAP7_75t_R output275 (.A(net275),
    .Y(text_out[113]));
 BUFx2_ASAP7_75t_R output276 (.A(net276),
    .Y(text_out[114]));
 BUFx2_ASAP7_75t_R output277 (.A(net277),
    .Y(text_out[115]));
 BUFx2_ASAP7_75t_R output278 (.A(net278),
    .Y(text_out[116]));
 BUFx2_ASAP7_75t_R output279 (.A(net279),
    .Y(text_out[117]));
 BUFx2_ASAP7_75t_R output280 (.A(net280),
    .Y(text_out[118]));
 BUFx2_ASAP7_75t_R output281 (.A(net281),
    .Y(text_out[119]));
 BUFx2_ASAP7_75t_R output282 (.A(net282),
    .Y(text_out[11]));
 BUFx2_ASAP7_75t_R output283 (.A(net283),
    .Y(text_out[120]));
 BUFx2_ASAP7_75t_R output284 (.A(net284),
    .Y(text_out[121]));
 BUFx2_ASAP7_75t_R output285 (.A(net285),
    .Y(text_out[122]));
 BUFx2_ASAP7_75t_R output286 (.A(net286),
    .Y(text_out[123]));
 BUFx2_ASAP7_75t_R output287 (.A(net287),
    .Y(text_out[124]));
 BUFx2_ASAP7_75t_R output288 (.A(net288),
    .Y(text_out[125]));
 BUFx2_ASAP7_75t_R output289 (.A(net289),
    .Y(text_out[126]));
 BUFx2_ASAP7_75t_R output290 (.A(net290),
    .Y(text_out[127]));
 BUFx2_ASAP7_75t_R output291 (.A(net291),
    .Y(text_out[12]));
 BUFx2_ASAP7_75t_R output292 (.A(net292),
    .Y(text_out[13]));
 BUFx2_ASAP7_75t_R output293 (.A(net293),
    .Y(text_out[14]));
 BUFx2_ASAP7_75t_R output294 (.A(net294),
    .Y(text_out[15]));
 BUFx2_ASAP7_75t_R output295 (.A(net295),
    .Y(text_out[16]));
 BUFx2_ASAP7_75t_R output296 (.A(net296),
    .Y(text_out[17]));
 BUFx2_ASAP7_75t_R output297 (.A(net297),
    .Y(text_out[18]));
 BUFx2_ASAP7_75t_R output298 (.A(net298),
    .Y(text_out[19]));
 BUFx2_ASAP7_75t_R output299 (.A(net299),
    .Y(text_out[1]));
 BUFx2_ASAP7_75t_R output300 (.A(net300),
    .Y(text_out[20]));
 BUFx2_ASAP7_75t_R output301 (.A(net301),
    .Y(text_out[21]));
 BUFx2_ASAP7_75t_R output302 (.A(net302),
    .Y(text_out[22]));
 BUFx2_ASAP7_75t_R output303 (.A(net303),
    .Y(text_out[23]));
 BUFx2_ASAP7_75t_R output304 (.A(net304),
    .Y(text_out[24]));
 BUFx2_ASAP7_75t_R output305 (.A(net305),
    .Y(text_out[25]));
 BUFx2_ASAP7_75t_R output306 (.A(net306),
    .Y(text_out[26]));
 BUFx2_ASAP7_75t_R output307 (.A(net307),
    .Y(text_out[27]));
 BUFx2_ASAP7_75t_R output308 (.A(net308),
    .Y(text_out[28]));
 BUFx2_ASAP7_75t_R output309 (.A(net309),
    .Y(text_out[29]));
 BUFx2_ASAP7_75t_R output310 (.A(net310),
    .Y(text_out[2]));
 BUFx2_ASAP7_75t_R output311 (.A(net311),
    .Y(text_out[30]));
 BUFx2_ASAP7_75t_R output312 (.A(net312),
    .Y(text_out[31]));
 BUFx2_ASAP7_75t_R output313 (.A(net313),
    .Y(text_out[32]));
 BUFx2_ASAP7_75t_R output314 (.A(net314),
    .Y(text_out[33]));
 BUFx2_ASAP7_75t_R output315 (.A(net315),
    .Y(text_out[34]));
 BUFx2_ASAP7_75t_R output316 (.A(net316),
    .Y(text_out[35]));
 BUFx2_ASAP7_75t_R output317 (.A(net317),
    .Y(text_out[36]));
 BUFx2_ASAP7_75t_R output318 (.A(net318),
    .Y(text_out[37]));
 BUFx2_ASAP7_75t_R output319 (.A(net319),
    .Y(text_out[38]));
 BUFx2_ASAP7_75t_R output320 (.A(net320),
    .Y(text_out[39]));
 BUFx2_ASAP7_75t_R output321 (.A(net321),
    .Y(text_out[3]));
 BUFx2_ASAP7_75t_R output322 (.A(net322),
    .Y(text_out[40]));
 BUFx2_ASAP7_75t_R output323 (.A(net323),
    .Y(text_out[41]));
 BUFx2_ASAP7_75t_R output324 (.A(net324),
    .Y(text_out[42]));
 BUFx2_ASAP7_75t_R output325 (.A(net325),
    .Y(text_out[43]));
 BUFx2_ASAP7_75t_R output326 (.A(net326),
    .Y(text_out[44]));
 BUFx2_ASAP7_75t_R output327 (.A(net327),
    .Y(text_out[45]));
 BUFx2_ASAP7_75t_R output328 (.A(net328),
    .Y(text_out[46]));
 BUFx2_ASAP7_75t_R output329 (.A(net329),
    .Y(text_out[47]));
 BUFx2_ASAP7_75t_R output330 (.A(net330),
    .Y(text_out[48]));
 BUFx2_ASAP7_75t_R output331 (.A(net331),
    .Y(text_out[49]));
 BUFx2_ASAP7_75t_R output332 (.A(net332),
    .Y(text_out[4]));
 BUFx2_ASAP7_75t_R output333 (.A(net333),
    .Y(text_out[50]));
 BUFx2_ASAP7_75t_R output334 (.A(net334),
    .Y(text_out[51]));
 BUFx2_ASAP7_75t_R output335 (.A(net335),
    .Y(text_out[52]));
 BUFx2_ASAP7_75t_R output336 (.A(net336),
    .Y(text_out[53]));
 BUFx2_ASAP7_75t_R output337 (.A(net337),
    .Y(text_out[54]));
 BUFx2_ASAP7_75t_R output338 (.A(net338),
    .Y(text_out[55]));
 BUFx2_ASAP7_75t_R output339 (.A(net339),
    .Y(text_out[56]));
 BUFx2_ASAP7_75t_R output340 (.A(net340),
    .Y(text_out[57]));
 BUFx2_ASAP7_75t_R output341 (.A(net341),
    .Y(text_out[58]));
 BUFx2_ASAP7_75t_R output342 (.A(net342),
    .Y(text_out[59]));
 BUFx2_ASAP7_75t_R output343 (.A(net343),
    .Y(text_out[5]));
 BUFx2_ASAP7_75t_R output344 (.A(net344),
    .Y(text_out[60]));
 BUFx2_ASAP7_75t_R output345 (.A(net345),
    .Y(text_out[61]));
 BUFx2_ASAP7_75t_R output346 (.A(net346),
    .Y(text_out[62]));
 BUFx2_ASAP7_75t_R output347 (.A(net347),
    .Y(text_out[63]));
 BUFx2_ASAP7_75t_R output348 (.A(net348),
    .Y(text_out[64]));
 BUFx2_ASAP7_75t_R output349 (.A(net349),
    .Y(text_out[65]));
 BUFx2_ASAP7_75t_R output350 (.A(net350),
    .Y(text_out[66]));
 BUFx2_ASAP7_75t_R output351 (.A(net351),
    .Y(text_out[67]));
 BUFx2_ASAP7_75t_R output352 (.A(net352),
    .Y(text_out[68]));
 BUFx2_ASAP7_75t_R output353 (.A(net353),
    .Y(text_out[69]));
 BUFx2_ASAP7_75t_R output354 (.A(net354),
    .Y(text_out[6]));
 BUFx2_ASAP7_75t_R output355 (.A(net355),
    .Y(text_out[70]));
 BUFx2_ASAP7_75t_R output356 (.A(net356),
    .Y(text_out[71]));
 BUFx2_ASAP7_75t_R output357 (.A(net357),
    .Y(text_out[72]));
 BUFx2_ASAP7_75t_R output358 (.A(net358),
    .Y(text_out[73]));
 BUFx2_ASAP7_75t_R output359 (.A(net359),
    .Y(text_out[74]));
 BUFx2_ASAP7_75t_R output360 (.A(net360),
    .Y(text_out[75]));
 BUFx2_ASAP7_75t_R output361 (.A(net361),
    .Y(text_out[76]));
 BUFx2_ASAP7_75t_R output362 (.A(net362),
    .Y(text_out[77]));
 BUFx2_ASAP7_75t_R output363 (.A(net363),
    .Y(text_out[78]));
 BUFx2_ASAP7_75t_R output364 (.A(net364),
    .Y(text_out[79]));
 BUFx2_ASAP7_75t_R output365 (.A(net365),
    .Y(text_out[7]));
 BUFx2_ASAP7_75t_R output366 (.A(net366),
    .Y(text_out[80]));
 BUFx2_ASAP7_75t_R output367 (.A(net367),
    .Y(text_out[81]));
 BUFx2_ASAP7_75t_R output368 (.A(net368),
    .Y(text_out[82]));
 BUFx2_ASAP7_75t_R output369 (.A(net369),
    .Y(text_out[83]));
 BUFx2_ASAP7_75t_R output370 (.A(net370),
    .Y(text_out[84]));
 BUFx2_ASAP7_75t_R output371 (.A(net371),
    .Y(text_out[85]));
 BUFx2_ASAP7_75t_R output372 (.A(net372),
    .Y(text_out[86]));
 BUFx2_ASAP7_75t_R output373 (.A(net373),
    .Y(text_out[87]));
 BUFx2_ASAP7_75t_R output374 (.A(net374),
    .Y(text_out[88]));
 BUFx2_ASAP7_75t_R output375 (.A(net375),
    .Y(text_out[89]));
 BUFx2_ASAP7_75t_R output376 (.A(net376),
    .Y(text_out[8]));
 BUFx2_ASAP7_75t_R output377 (.A(net377),
    .Y(text_out[90]));
 BUFx2_ASAP7_75t_R output378 (.A(net378),
    .Y(text_out[91]));
 BUFx2_ASAP7_75t_R output379 (.A(net379),
    .Y(text_out[92]));
 BUFx2_ASAP7_75t_R output380 (.A(net380),
    .Y(text_out[93]));
 BUFx2_ASAP7_75t_R output381 (.A(net381),
    .Y(text_out[94]));
 BUFx2_ASAP7_75t_R output382 (.A(net382),
    .Y(text_out[95]));
 BUFx2_ASAP7_75t_R output383 (.A(net383),
    .Y(text_out[96]));
 BUFx2_ASAP7_75t_R output384 (.A(net384),
    .Y(text_out[97]));
 BUFx2_ASAP7_75t_R output385 (.A(net385),
    .Y(text_out[98]));
 BUFx2_ASAP7_75t_R output386 (.A(net386),
    .Y(text_out[99]));
 BUFx2_ASAP7_75t_R output387 (.A(net387),
    .Y(text_out[9]));
 BUFx3_ASAP7_75t_R place4424 (.A(_06665_),
    .Y(net4424));
 BUFx3_ASAP7_75t_R place4425 (.A(_05362_),
    .Y(net4425));
 BUFx3_ASAP7_75t_R place4426 (.A(_02569_),
    .Y(net4426));
 BUFx3_ASAP7_75t_R place4427 (.A(_06883_),
    .Y(net4427));
 BUFx3_ASAP7_75t_R place4428 (.A(_06877_),
    .Y(net4428));
 BUFx3_ASAP7_75t_R place4429 (.A(_05339_),
    .Y(net4429));
 BUFx3_ASAP7_75t_R place4430 (.A(_05339_),
    .Y(net4430));
 BUFx3_ASAP7_75t_R place4431 (.A(_05339_),
    .Y(net4431));
 BUFx3_ASAP7_75t_R place4432 (.A(_03292_),
    .Y(net4432));
 BUFx3_ASAP7_75t_R place4433 (.A(_02514_),
    .Y(net4433));
 BUFx3_ASAP7_75t_R place4434 (.A(_13034_),
    .Y(net4434));
 BUFx3_ASAP7_75t_R place4435 (.A(_12630_),
    .Y(net4435));
 BUFx3_ASAP7_75t_R place4436 (.A(_06824_),
    .Y(net4436));
 BUFx3_ASAP7_75t_R place4437 (.A(_06742_),
    .Y(net4437));
 BUFx3_ASAP7_75t_R place4438 (.A(_05584_),
    .Y(net4438));
 BUFx3_ASAP7_75t_R place4439 (.A(_05224_),
    .Y(net4439));
 BUFx3_ASAP7_75t_R place4440 (.A(_04750_),
    .Y(net4440));
 BUFx3_ASAP7_75t_R place4441 (.A(_03914_),
    .Y(net4441));
 BUFx6f_ASAP7_75t_R place4442 (.A(_02581_),
    .Y(net4442));
 BUFx3_ASAP7_75t_R place4443 (.A(_02564_),
    .Y(net4443));
 BUFx3_ASAP7_75t_R place4444 (.A(_02522_),
    .Y(net4444));
 BUFx3_ASAP7_75t_R place4445 (.A(_02460_),
    .Y(net4445));
 BUFx6f_ASAP7_75t_R place4446 (.A(_02374_),
    .Y(net4446));
 BUFx3_ASAP7_75t_R place4447 (.A(_13806_),
    .Y(net4447));
 BUFx3_ASAP7_75t_R place4448 (.A(_13645_),
    .Y(net4448));
 BUFx3_ASAP7_75t_R place4449 (.A(_13642_),
    .Y(net4449));
 BUFx3_ASAP7_75t_R place4450 (.A(_07372_),
    .Y(net4450));
 BUFx6f_ASAP7_75t_R place4451 (.A(_06662_),
    .Y(net4451));
 BUFx3_ASAP7_75t_R place4452 (.A(_06662_),
    .Y(net4452));
 BUFx3_ASAP7_75t_R place4453 (.A(net4454),
    .Y(net4453));
 BUFx3_ASAP7_75t_R place4454 (.A(_06536_),
    .Y(net4454));
 BUFx3_ASAP7_75t_R place4455 (.A(_06038_),
    .Y(net4455));
 BUFx3_ASAP7_75t_R place4456 (.A(_05427_),
    .Y(net4456));
 BUFx3_ASAP7_75t_R place4457 (.A(_05359_),
    .Y(net4457));
 BUFx3_ASAP7_75t_R place4458 (.A(_05150_),
    .Y(net4458));
 BUFx3_ASAP7_75t_R place4459 (.A(_04516_),
    .Y(net4459));
 BUFx3_ASAP7_75t_R place4460 (.A(_04516_),
    .Y(net4460));
 BUFx3_ASAP7_75t_R place4461 (.A(_04479_),
    .Y(net4461));
 BUFx6f_ASAP7_75t_R place4462 (.A(_03734_),
    .Y(net4462));
 BUFx3_ASAP7_75t_R place4463 (.A(_03217_),
    .Y(net4463));
 BUFx3_ASAP7_75t_R place4464 (.A(_02513_),
    .Y(net4464));
 BUFx3_ASAP7_75t_R place4465 (.A(_02513_),
    .Y(net4465));
 BUFx3_ASAP7_75t_R place4466 (.A(_02479_),
    .Y(net4466));
 BUFx3_ASAP7_75t_R place4467 (.A(_02468_),
    .Y(net4467));
 BUFx3_ASAP7_75t_R place4468 (.A(_02382_),
    .Y(net4468));
 BUFx3_ASAP7_75t_R place4469 (.A(_14023_),
    .Y(net4469));
 BUFx3_ASAP7_75t_R place4470 (.A(_13937_),
    .Y(net4470));
 BUFx3_ASAP7_75t_R place4471 (.A(_13937_),
    .Y(net4471));
 BUFx3_ASAP7_75t_R place4472 (.A(_13711_),
    .Y(net4472));
 BUFx3_ASAP7_75t_R place4473 (.A(_13621_),
    .Y(net4473));
 BUFx3_ASAP7_75t_R place4474 (.A(_13621_),
    .Y(net4474));
 BUFx3_ASAP7_75t_R place4475 (.A(_13254_),
    .Y(net4475));
 BUFx6f_ASAP7_75t_R place4476 (.A(_13033_),
    .Y(net4476));
 BUFx3_ASAP7_75t_R place4477 (.A(_13033_),
    .Y(net4477));
 BUFx3_ASAP7_75t_R place4478 (.A(_12542_),
    .Y(net4478));
 BUFx6f_ASAP7_75t_R place4479 (.A(_12416_),
    .Y(net4479));
 BUFx3_ASAP7_75t_R place4480 (.A(_12416_),
    .Y(net4480));
 BUFx6f_ASAP7_75t_R place4481 (.A(_11597_),
    .Y(net4481));
 BUFx3_ASAP7_75t_R place4482 (.A(_07355_),
    .Y(net4482));
 BUFx3_ASAP7_75t_R place4483 (.A(_06944_),
    .Y(net4483));
 BUFx3_ASAP7_75t_R place4484 (.A(net4485),
    .Y(net4484));
 BUFx3_ASAP7_75t_R place4485 (.A(_06868_),
    .Y(net4485));
 BUFx3_ASAP7_75t_R place4486 (.A(_06804_),
    .Y(net4486));
 BUFx3_ASAP7_75t_R place4487 (.A(_06680_),
    .Y(net4487));
 BUFx3_ASAP7_75t_R place4488 (.A(_06670_),
    .Y(net4488));
 BUFx3_ASAP7_75t_R place4489 (.A(_06670_),
    .Y(net4489));
 BUFx3_ASAP7_75t_R place4490 (.A(_06670_),
    .Y(net4490));
 BUFx3_ASAP7_75t_R place4491 (.A(_06599_),
    .Y(net4491));
 BUFx3_ASAP7_75t_R place4492 (.A(_06515_),
    .Y(net4492));
 BUFx3_ASAP7_75t_R place4493 (.A(_05519_),
    .Y(net4493));
 BUFx3_ASAP7_75t_R place4494 (.A(_05451_),
    .Y(net4494));
 BUFx3_ASAP7_75t_R place4495 (.A(_05343_),
    .Y(net4495));
 BUFx3_ASAP7_75t_R place4496 (.A(_05243_),
    .Y(net4496));
 BUFx3_ASAP7_75t_R place4497 (.A(_05008_),
    .Y(net4497));
 BUFx3_ASAP7_75t_R place4498 (.A(_04944_),
    .Y(net4498));
 BUFx3_ASAP7_75t_R place4499 (.A(_04727_),
    .Y(net4499));
 BUFx3_ASAP7_75t_R place4500 (.A(_04595_),
    .Y(net4500));
 BUFx3_ASAP7_75t_R place4501 (.A(_04591_),
    .Y(net4501));
 BUFx6f_ASAP7_75t_R place4502 (.A(_03987_),
    .Y(net4502));
 BUFx3_ASAP7_75t_R place4503 (.A(_03987_),
    .Y(net4503));
 BUFx3_ASAP7_75t_R place4504 (.A(_03907_),
    .Y(net4504));
 BUFx3_ASAP7_75t_R place4505 (.A(_03804_),
    .Y(net4505));
 BUFx3_ASAP7_75t_R place4506 (.A(_03226_),
    .Y(net4506));
 BUFx3_ASAP7_75t_R place4507 (.A(_03177_),
    .Y(net4507));
 BUFx3_ASAP7_75t_R place4508 (.A(_02532_),
    .Y(net4508));
 BUFx3_ASAP7_75t_R place4509 (.A(_02507_),
    .Y(net4509));
 BUFx3_ASAP7_75t_R place4510 (.A(_02489_),
    .Y(net4510));
 BUFx3_ASAP7_75t_R place4511 (.A(_02489_),
    .Y(net4511));
 BUFx3_ASAP7_75t_R place4512 (.A(_02474_),
    .Y(net4512));
 BUFx3_ASAP7_75t_R place4513 (.A(_02459_),
    .Y(net4513));
 BUFx3_ASAP7_75t_R place4514 (.A(_02459_),
    .Y(net4514));
 BUFx3_ASAP7_75t_R place4515 (.A(_02373_),
    .Y(net4515));
 BUFx3_ASAP7_75t_R place4516 (.A(_02015_),
    .Y(net4516));
 BUFx3_ASAP7_75t_R place4517 (.A(_15369_),
    .Y(net4517));
 BUFx3_ASAP7_75t_R place4518 (.A(_15256_),
    .Y(net4518));
 BUFx3_ASAP7_75t_R place4519 (.A(_13930_),
    .Y(net4519));
 BUFx3_ASAP7_75t_R place4520 (.A(_13804_),
    .Y(net4520));
 BUFx3_ASAP7_75t_R place4521 (.A(_13644_),
    .Y(net4521));
 BUFx3_ASAP7_75t_R place4522 (.A(_13618_),
    .Y(net4522));
 BUFx3_ASAP7_75t_R place4523 (.A(_13260_),
    .Y(net4523));
 BUFx6f_ASAP7_75t_R place4524 (.A(_12905_),
    .Y(net4524));
 BUFx3_ASAP7_75t_R place4525 (.A(_12666_),
    .Y(net4525));
 BUFx3_ASAP7_75t_R place4526 (.A(_12554_),
    .Y(net4526));
 BUFx3_ASAP7_75t_R place4527 (.A(_11118_),
    .Y(net4527));
 BUFx3_ASAP7_75t_R place4528 (.A(_09954_),
    .Y(net4528));
 BUFx6f_ASAP7_75t_R place4529 (.A(_09846_),
    .Y(net4529));
 BUFx3_ASAP7_75t_R place4530 (.A(_09419_),
    .Y(net4530));
 BUFx3_ASAP7_75t_R place4531 (.A(_08119_),
    .Y(net4531));
 BUFx3_ASAP7_75t_R place4532 (.A(_08108_),
    .Y(net4532));
 BUFx3_ASAP7_75t_R place4533 (.A(_07273_),
    .Y(net4533));
 BUFx3_ASAP7_75t_R place4534 (.A(_07273_),
    .Y(net4534));
 BUFx3_ASAP7_75t_R place4535 (.A(_06654_),
    .Y(net4535));
 BUFx3_ASAP7_75t_R place4536 (.A(_06654_),
    .Y(net4536));
 BUFx3_ASAP7_75t_R place4537 (.A(_06532_),
    .Y(net4537));
 BUFx6f_ASAP7_75t_R place4538 (.A(_06520_),
    .Y(net4538));
 BUFx3_ASAP7_75t_R place4539 (.A(_06520_),
    .Y(net4539));
 BUFx3_ASAP7_75t_R place4540 (.A(_06100_),
    .Y(net4540));
 BUFx6f_ASAP7_75t_R place4541 (.A(_05915_),
    .Y(net4541));
 BUFx3_ASAP7_75t_R place4542 (.A(_05915_),
    .Y(net4542));
 BUFx3_ASAP7_75t_R place4543 (.A(_05281_),
    .Y(net4543));
 BUFx3_ASAP7_75t_R place4544 (.A(_05162_),
    .Y(net4544));
 BUFx3_ASAP7_75t_R place4545 (.A(_05162_),
    .Y(net4545));
 BUFx3_ASAP7_75t_R place4546 (.A(_05149_),
    .Y(net4546));
 BUFx3_ASAP7_75t_R place4547 (.A(_04806_),
    .Y(net4547));
 BUFx3_ASAP7_75t_R place4548 (.A(net4549),
    .Y(net4548));
 BUFx6f_ASAP7_75t_R place4549 (.A(_04616_),
    .Y(net4549));
 BUFx3_ASAP7_75t_R place4550 (.A(_04515_),
    .Y(net4550));
 BUFx3_ASAP7_75t_R place4551 (.A(_04478_),
    .Y(net4551));
 BUFx3_ASAP7_75t_R place4552 (.A(_04458_),
    .Y(net4552));
 BUFx3_ASAP7_75t_R place4553 (.A(_03854_),
    .Y(net4553));
 BUFx3_ASAP7_75t_R place4554 (.A(_03826_),
    .Y(net4554));
 BUFx3_ASAP7_75t_R place4555 (.A(_03733_),
    .Y(net4555));
 BUFx6f_ASAP7_75t_R place4556 (.A(_03249_),
    .Y(net4556));
 BUFx3_ASAP7_75t_R place4557 (.A(_03228_),
    .Y(net4557));
 BUFx6f_ASAP7_75t_R place4558 (.A(_03118_),
    .Y(net4558));
 BUFx3_ASAP7_75t_R place4559 (.A(net4561),
    .Y(net4559));
 BUFx3_ASAP7_75t_R place4560 (.A(net4561),
    .Y(net4560));
 BUFx3_ASAP7_75t_R place4561 (.A(_02478_),
    .Y(net4561));
 BUFx3_ASAP7_75t_R place4562 (.A(_02467_),
    .Y(net4562));
 BUFx3_ASAP7_75t_R place4563 (.A(net4565),
    .Y(net4563));
 BUFx3_ASAP7_75t_R place4564 (.A(net4565),
    .Y(net4564));
 BUFx6f_ASAP7_75t_R place4565 (.A(_02381_),
    .Y(net4565));
 BUFx3_ASAP7_75t_R place4566 (.A(_01817_),
    .Y(net4566));
 BUFx3_ASAP7_75t_R place4567 (.A(_01746_),
    .Y(net4567));
 BUFx3_ASAP7_75t_R place4568 (.A(_01723_),
    .Y(net4568));
 BUFx3_ASAP7_75t_R place4569 (.A(_15191_),
    .Y(net4569));
 BUFx6f_ASAP7_75t_R place4570 (.A(_15191_),
    .Y(net4570));
 BUFx3_ASAP7_75t_R place4571 (.A(_14648_),
    .Y(net4571));
 BUFx3_ASAP7_75t_R place4572 (.A(_14319_),
    .Y(net4572));
 BUFx6f_ASAP7_75t_R place4573 (.A(_13772_),
    .Y(net4573));
 BUFx6f_ASAP7_75t_R place4574 (.A(_13659_),
    .Y(net4574));
 BUFx3_ASAP7_75t_R place4575 (.A(_13659_),
    .Y(net4575));
 BUFx3_ASAP7_75t_R place4576 (.A(_13147_),
    .Y(net4576));
 BUFx6f_ASAP7_75t_R place4577 (.A(_13100_),
    .Y(net4577));
 BUFx3_ASAP7_75t_R place4578 (.A(_13032_),
    .Y(net4578));
 BUFx3_ASAP7_75t_R place4579 (.A(_13030_),
    .Y(net4579));
 BUFx6f_ASAP7_75t_R place4580 (.A(_13030_),
    .Y(net4580));
 BUFx3_ASAP7_75t_R place4581 (.A(_12925_),
    .Y(net4581));
 BUFx3_ASAP7_75t_R place4582 (.A(_12925_),
    .Y(net4582));
 BUFx3_ASAP7_75t_R place4583 (.A(_12377_),
    .Y(net4583));
 BUFx3_ASAP7_75t_R place4584 (.A(_12350_),
    .Y(net4584));
 BUFx3_ASAP7_75t_R place4585 (.A(_12229_),
    .Y(net4585));
 BUFx6f_ASAP7_75t_R place4586 (.A(_12226_),
    .Y(net4586));
 BUFx3_ASAP7_75t_R place4587 (.A(_12226_),
    .Y(net4587));
 BUFx3_ASAP7_75t_R place4588 (.A(_11697_),
    .Y(net4588));
 BUFx3_ASAP7_75t_R place4589 (.A(_11644_),
    .Y(net4589));
 BUFx3_ASAP7_75t_R place4590 (.A(net4591),
    .Y(net4590));
 BUFx3_ASAP7_75t_R place4591 (.A(_11596_),
    .Y(net4591));
 BUFx3_ASAP7_75t_R place4592 (.A(_10954_),
    .Y(net4592));
 BUFx3_ASAP7_75t_R place4593 (.A(_10920_),
    .Y(net4593));
 BUFx3_ASAP7_75t_R place4594 (.A(_10904_),
    .Y(net4594));
 BUFx6f_ASAP7_75t_R place4595 (.A(_10904_),
    .Y(net4595));
 BUFx3_ASAP7_75t_R place4596 (.A(_09329_),
    .Y(net4596));
 BUFx3_ASAP7_75t_R place4597 (.A(_09168_),
    .Y(net4597));
 BUFx6f_ASAP7_75t_R place4598 (.A(_09168_),
    .Y(net4598));
 BUFx3_ASAP7_75t_R place4599 (.A(_09078_),
    .Y(net4599));
 BUFx3_ASAP7_75t_R place4600 (.A(_09078_),
    .Y(net4600));
 BUFx3_ASAP7_75t_R place4601 (.A(_08297_),
    .Y(net4601));
 BUFx3_ASAP7_75t_R place4602 (.A(_08114_),
    .Y(net4602));
 BUFx3_ASAP7_75t_R place4603 (.A(_08114_),
    .Y(net4603));
 BUFx3_ASAP7_75t_R place4604 (.A(_07300_),
    .Y(net4604));
 BUFx3_ASAP7_75t_R place4605 (.A(_07214_),
    .Y(net4605));
 BUFx3_ASAP7_75t_R place4606 (.A(_07205_),
    .Y(net4606));
 BUFx3_ASAP7_75t_R place4607 (.A(_07041_),
    .Y(net4607));
 BUFx3_ASAP7_75t_R place4608 (.A(_06803_),
    .Y(net4608));
 BUFx3_ASAP7_75t_R place4609 (.A(_06702_),
    .Y(net4609));
 BUFx3_ASAP7_75t_R place4610 (.A(_06666_),
    .Y(net4610));
 BUFx3_ASAP7_75t_R place4611 (.A(_06648_),
    .Y(net4611));
 BUFx3_ASAP7_75t_R place4612 (.A(_06645_),
    .Y(net4612));
 BUFx6f_ASAP7_75t_R place4613 (.A(_06614_),
    .Y(net4613));
 BUFx3_ASAP7_75t_R place4614 (.A(_06606_),
    .Y(net4614));
 BUFx3_ASAP7_75t_R place4615 (.A(_06606_),
    .Y(net4615));
 BUFx3_ASAP7_75t_R place4616 (.A(_06598_),
    .Y(net4616));
 BUFx3_ASAP7_75t_R place4617 (.A(_06584_),
    .Y(net4617));
 BUFx3_ASAP7_75t_R place4618 (.A(_06202_),
    .Y(net4618));
 BUFx3_ASAP7_75t_R place4619 (.A(_05429_),
    .Y(net4619));
 BUFx3_ASAP7_75t_R place4620 (.A(_05429_),
    .Y(net4620));
 BUFx3_ASAP7_75t_R place4621 (.A(_05419_),
    .Y(net4621));
 BUFx6f_ASAP7_75t_R place4622 (.A(_05419_),
    .Y(net4622));
 BUFx3_ASAP7_75t_R place4623 (.A(_05380_),
    .Y(net4623));
 BUFx3_ASAP7_75t_R place4624 (.A(_05336_),
    .Y(net4624));
 BUFx3_ASAP7_75t_R place4625 (.A(_05324_),
    .Y(net4625));
 BUFx3_ASAP7_75t_R place4626 (.A(_05320_),
    .Y(net4626));
 BUFx6f_ASAP7_75t_R place4627 (.A(_05320_),
    .Y(net4627));
 BUFx6f_ASAP7_75t_R place4628 (.A(_05319_),
    .Y(net4628));
 BUFx3_ASAP7_75t_R place4629 (.A(_05287_),
    .Y(net4629));
 BUFx3_ASAP7_75t_R place4630 (.A(_05222_),
    .Y(net4630));
 BUFx3_ASAP7_75t_R place4631 (.A(_04912_),
    .Y(net4631));
 BUFx3_ASAP7_75t_R place4632 (.A(_04772_),
    .Y(net4632));
 BUFx3_ASAP7_75t_R place4633 (.A(_04734_),
    .Y(net4633));
 BUFx3_ASAP7_75t_R place4634 (.A(_04684_),
    .Y(net4634));
 BUFx3_ASAP7_75t_R place4635 (.A(_04641_),
    .Y(net4635));
 BUFx6f_ASAP7_75t_R place4636 (.A(_04590_),
    .Y(net4636));
 BUFx3_ASAP7_75t_R place4637 (.A(_04590_),
    .Y(net4637));
 BUFx3_ASAP7_75t_R place4638 (.A(_04585_),
    .Y(net4638));
 BUFx3_ASAP7_75t_R place4639 (.A(_04566_),
    .Y(net4639));
 BUFx3_ASAP7_75t_R place4640 (.A(_04566_),
    .Y(net4640));
 BUFx3_ASAP7_75t_R place4641 (.A(_04555_),
    .Y(net4641));
 BUFx6f_ASAP7_75t_R place4642 (.A(_03906_),
    .Y(net4642));
 BUFx6f_ASAP7_75t_R place4643 (.A(_03888_),
    .Y(net4643));
 BUFx3_ASAP7_75t_R place4644 (.A(_03888_),
    .Y(net4644));
 BUFx3_ASAP7_75t_R place4645 (.A(_03885_),
    .Y(net4645));
 BUFx3_ASAP7_75t_R place4646 (.A(_03852_),
    .Y(net4646));
 BUFx3_ASAP7_75t_R place4647 (.A(_03803_),
    .Y(net4647));
 BUFx6f_ASAP7_75t_R place4648 (.A(_03795_),
    .Y(net4648));
 BUFx3_ASAP7_75t_R place4649 (.A(_03740_),
    .Y(net4649));
 BUFx3_ASAP7_75t_R place4650 (.A(_03375_),
    .Y(net4650));
 BUFx3_ASAP7_75t_R place4651 (.A(_03254_),
    .Y(net4651));
 BUFx3_ASAP7_75t_R place4652 (.A(_03225_),
    .Y(net4652));
 BUFx3_ASAP7_75t_R place4653 (.A(_03179_),
    .Y(net4653));
 BUFx3_ASAP7_75t_R place4654 (.A(_03160_),
    .Y(net4654));
 BUFx3_ASAP7_75t_R place4655 (.A(_03138_),
    .Y(net4655));
 BUFx3_ASAP7_75t_R place4656 (.A(_03113_),
    .Y(net4656));
 BUFx3_ASAP7_75t_R place4657 (.A(_03113_),
    .Y(net4657));
 BUFx3_ASAP7_75t_R place4658 (.A(_02909_),
    .Y(net4658));
 BUFx3_ASAP7_75t_R place4659 (.A(_02783_),
    .Y(net4659));
 BUFx3_ASAP7_75t_R place4660 (.A(_02651_),
    .Y(net4660));
 BUFx3_ASAP7_75t_R place4661 (.A(_02502_),
    .Y(net4661));
 BUFx3_ASAP7_75t_R place4662 (.A(_02495_),
    .Y(net4662));
 BUFx3_ASAP7_75t_R place4663 (.A(_02495_),
    .Y(net4663));
 BUFx3_ASAP7_75t_R place4664 (.A(_02488_),
    .Y(net4664));
 BUFx3_ASAP7_75t_R place4665 (.A(_02446_),
    .Y(net4665));
 BUFx3_ASAP7_75t_R place4666 (.A(_02395_),
    .Y(net4666));
 BUFx3_ASAP7_75t_R place4667 (.A(_02177_),
    .Y(net4667));
 BUFx6f_ASAP7_75t_R place4668 (.A(_01946_),
    .Y(net4668));
 BUFx3_ASAP7_75t_R place4669 (.A(_01716_),
    .Y(net4669));
 BUFx3_ASAP7_75t_R place4670 (.A(_01707_),
    .Y(net4670));
 BUFx3_ASAP7_75t_R place4671 (.A(_15381_),
    .Y(net4671));
 BUFx3_ASAP7_75t_R place4672 (.A(_15291_),
    .Y(net4672));
 BUFx3_ASAP7_75t_R place4673 (.A(_15142_),
    .Y(net4673));
 BUFx3_ASAP7_75t_R place4674 (.A(_15094_),
    .Y(net4674));
 BUFx3_ASAP7_75t_R place4675 (.A(_15071_),
    .Y(net4675));
 BUFx3_ASAP7_75t_R place4676 (.A(_15069_),
    .Y(net4676));
 BUFx3_ASAP7_75t_R place4677 (.A(_15005_),
    .Y(net4677));
 BUFx3_ASAP7_75t_R place4678 (.A(_14521_),
    .Y(net4678));
 BUFx3_ASAP7_75t_R place4679 (.A(_14454_),
    .Y(net4679));
 BUFx3_ASAP7_75t_R place4680 (.A(_13904_),
    .Y(net4680));
 BUFx3_ASAP7_75t_R place4681 (.A(_13791_),
    .Y(net4681));
 BUFx3_ASAP7_75t_R place4682 (.A(_13754_),
    .Y(net4682));
 BUFx3_ASAP7_75t_R place4683 (.A(_13616_),
    .Y(net4683));
 BUFx3_ASAP7_75t_R place4684 (.A(net4685),
    .Y(net4684));
 BUFx6f_ASAP7_75t_R place4685 (.A(_13616_),
    .Y(net4685));
 BUFx3_ASAP7_75t_R place4686 (.A(_13614_),
    .Y(net4686));
 BUFx3_ASAP7_75t_R place4687 (.A(_13379_),
    .Y(net4687));
 BUFx3_ASAP7_75t_R place4688 (.A(_13212_),
    .Y(net4688));
 BUFx6f_ASAP7_75t_R place4689 (.A(_13172_),
    .Y(net4689));
 BUFx3_ASAP7_75t_R place4690 (.A(_13110_),
    .Y(net4690));
 BUFx3_ASAP7_75t_R place4691 (.A(_12993_),
    .Y(net4691));
 BUFx3_ASAP7_75t_R place4692 (.A(_12988_),
    .Y(net4692));
 BUFx3_ASAP7_75t_R place4693 (.A(_12953_),
    .Y(net4693));
 BUFx3_ASAP7_75t_R place4694 (.A(_12575_),
    .Y(net4694));
 BUFx3_ASAP7_75t_R place4695 (.A(_12529_),
    .Y(net4695));
 BUFx3_ASAP7_75t_R place4696 (.A(_12361_),
    .Y(net4696));
 BUFx3_ASAP7_75t_R place4697 (.A(_12305_),
    .Y(net4697));
 BUFx3_ASAP7_75t_R place4698 (.A(_12287_),
    .Y(net4698));
 BUFx3_ASAP7_75t_R place4699 (.A(_12207_),
    .Y(net4699));
 BUFx3_ASAP7_75t_R place4700 (.A(_12205_),
    .Y(net4700));
 BUFx3_ASAP7_75t_R place4701 (.A(_11841_),
    .Y(net4701));
 BUFx3_ASAP7_75t_R place4702 (.A(_11696_),
    .Y(net4702));
 BUFx3_ASAP7_75t_R place4703 (.A(_11589_),
    .Y(net4703));
 BUFx3_ASAP7_75t_R place4704 (.A(_11138_),
    .Y(net4704));
 BUFx3_ASAP7_75t_R place4705 (.A(_11117_),
    .Y(net4705));
 BUFx3_ASAP7_75t_R place4706 (.A(_11009_),
    .Y(net4706));
 BUFx3_ASAP7_75t_R place4707 (.A(_11003_),
    .Y(net4707));
 BUFx3_ASAP7_75t_R place4708 (.A(_10900_),
    .Y(net4708));
 BUFx3_ASAP7_75t_R place4709 (.A(_10793_),
    .Y(net4709));
 BUFx3_ASAP7_75t_R place4710 (.A(_10375_),
    .Y(net4710));
 BUFx3_ASAP7_75t_R place4711 (.A(_09375_),
    .Y(net4711));
 BUFx3_ASAP7_75t_R place4712 (.A(_09336_),
    .Y(net4712));
 BUFx6f_ASAP7_75t_R place4713 (.A(_09252_),
    .Y(net4713));
 BUFx6f_ASAP7_75t_R place4714 (.A(_09090_),
    .Y(net4714));
 BUFx3_ASAP7_75t_R place4715 (.A(_08255_),
    .Y(net4715));
 BUFx3_ASAP7_75t_R place4716 (.A(_08255_),
    .Y(net4716));
 BUFx3_ASAP7_75t_R place4717 (.A(_08249_),
    .Y(net4717));
 BUFx3_ASAP7_75t_R place4718 (.A(_08218_),
    .Y(net4718));
 BUFx3_ASAP7_75t_R place4719 (.A(_08107_),
    .Y(net4719));
 BUFx3_ASAP7_75t_R place4720 (.A(_01366_),
    .Y(net4720));
 BUFx3_ASAP7_75t_R place4721 (.A(_01324_),
    .Y(net4721));
 BUFx3_ASAP7_75t_R place4722 (.A(net4723),
    .Y(net4722));
 BUFx3_ASAP7_75t_R place4723 (.A(_01232_),
    .Y(net4723));
 BUFx6f_ASAP7_75t_R place4724 (.A(_07566_),
    .Y(net4724));
 BUFx3_ASAP7_75t_R place4725 (.A(_07267_),
    .Y(net4725));
 BUFx6f_ASAP7_75t_R place4726 (.A(_07253_),
    .Y(net4726));
 BUFx6f_ASAP7_75t_R place4727 (.A(_07212_),
    .Y(net4727));
 BUFx3_ASAP7_75t_R place4728 (.A(_05882_),
    .Y(net4728));
 BUFx3_ASAP7_75t_R place4729 (.A(_05810_),
    .Y(net4729));
 BUFx3_ASAP7_75t_R place4730 (.A(_04460_),
    .Y(net4730));
 BUFx3_ASAP7_75t_R place4731 (.A(_04460_),
    .Y(net4731));
 BUFx6f_ASAP7_75t_R place4732 (.A(_03894_),
    .Y(net4732));
 BUFx3_ASAP7_75t_R place4733 (.A(_03894_),
    .Y(net4733));
 BUFx3_ASAP7_75t_R place4734 (.A(_03894_),
    .Y(net4734));
 BUFx3_ASAP7_75t_R place4735 (.A(_03853_),
    .Y(net4735));
 BUFx3_ASAP7_75t_R place4736 (.A(_03830_),
    .Y(net4736));
 BUFx3_ASAP7_75t_R place4737 (.A(_03732_),
    .Y(net4737));
 BUFx3_ASAP7_75t_R place4738 (.A(_03142_),
    .Y(net4738));
 BUFx3_ASAP7_75t_R place4739 (.A(_03107_),
    .Y(net4739));
 BUFx6f_ASAP7_75t_R place4740 (.A(_03080_),
    .Y(net4740));
 BUFx3_ASAP7_75t_R place4741 (.A(_01917_),
    .Y(net4741));
 BUFx3_ASAP7_75t_R place4742 (.A(_01828_),
    .Y(net4742));
 BUFx6f_ASAP7_75t_R place4743 (.A(_01794_),
    .Y(net4743));
 BUFx3_ASAP7_75t_R place4744 (.A(_01794_),
    .Y(net4744));
 BUFx3_ASAP7_75t_R place4745 (.A(_01767_),
    .Y(net4745));
 BUFx3_ASAP7_75t_R place4746 (.A(_01745_),
    .Y(net4746));
 BUFx6f_ASAP7_75t_R place4747 (.A(_01722_),
    .Y(net4747));
 BUFx3_ASAP7_75t_R place4748 (.A(_15355_),
    .Y(net4748));
 BUFx3_ASAP7_75t_R place4749 (.A(_15238_),
    .Y(net4749));
 BUFx3_ASAP7_75t_R place4750 (.A(_15185_),
    .Y(net4750));
 BUFx3_ASAP7_75t_R place4751 (.A(_15185_),
    .Y(net4751));
 BUFx3_ASAP7_75t_R place4752 (.A(net4753),
    .Y(net4752));
 BUFx6f_ASAP7_75t_R place4753 (.A(_15035_),
    .Y(net4753));
 BUFx3_ASAP7_75t_R place4754 (.A(net4755),
    .Y(net4754));
 BUFx3_ASAP7_75t_R place4755 (.A(_15035_),
    .Y(net4755));
 BUFx3_ASAP7_75t_R place4756 (.A(_14554_),
    .Y(net4756));
 BUFx3_ASAP7_75t_R place4757 (.A(_14477_),
    .Y(net4757));
 BUFx6f_ASAP7_75t_R place4758 (.A(_14403_),
    .Y(net4758));
 BUFx3_ASAP7_75t_R place4759 (.A(_14318_),
    .Y(net4759));
 BUFx3_ASAP7_75t_R place4760 (.A(_14318_),
    .Y(net4760));
 BUFx3_ASAP7_75t_R place4761 (.A(net4763),
    .Y(net4761));
 BUFx3_ASAP7_75t_R place4762 (.A(net4763),
    .Y(net4762));
 BUFx3_ASAP7_75t_R place4763 (.A(_13619_),
    .Y(net4763));
 BUFx3_ASAP7_75t_R place4764 (.A(_13021_),
    .Y(net4764));
 BUFx3_ASAP7_75t_R place4765 (.A(_12947_),
    .Y(net4765));
 BUFx3_ASAP7_75t_R place4766 (.A(_12924_),
    .Y(net4766));
 BUFx3_ASAP7_75t_R place4767 (.A(_12349_),
    .Y(net4767));
 BUFx3_ASAP7_75t_R place4768 (.A(_12185_),
    .Y(net4768));
 BUFx3_ASAP7_75t_R place4769 (.A(_11920_),
    .Y(net4769));
 BUFx3_ASAP7_75t_R place4770 (.A(_11762_),
    .Y(net4770));
 BUFx3_ASAP7_75t_R place4771 (.A(_11628_),
    .Y(net4771));
 BUFx3_ASAP7_75t_R place4772 (.A(_11619_),
    .Y(net4772));
 BUFx3_ASAP7_75t_R place4773 (.A(net4775),
    .Y(net4773));
 BUFx3_ASAP7_75t_R place4774 (.A(net4775),
    .Y(net4774));
 BUFx6f_ASAP7_75t_R place4775 (.A(_11595_),
    .Y(net4775));
 BUFx3_ASAP7_75t_R place4776 (.A(_11141_),
    .Y(net4776));
 BUFx3_ASAP7_75t_R place4777 (.A(_11038_),
    .Y(net4777));
 BUFx3_ASAP7_75t_R place4778 (.A(_10919_),
    .Y(net4778));
 BUFx3_ASAP7_75t_R place4779 (.A(_10902_),
    .Y(net4779));
 BUFx3_ASAP7_75t_R place4780 (.A(net4781),
    .Y(net4780));
 BUFx3_ASAP7_75t_R place4781 (.A(_10902_),
    .Y(net4781));
 BUFx3_ASAP7_75t_R place4782 (.A(_09891_),
    .Y(net4782));
 BUFx6f_ASAP7_75t_R place4783 (.A(_09828_),
    .Y(net4783));
 BUFx6f_ASAP7_75t_R place4784 (.A(_09605_),
    .Y(net4784));
 BUFx3_ASAP7_75t_R place4785 (.A(_09605_),
    .Y(net4785));
 BUFx3_ASAP7_75t_R place4786 (.A(_09384_),
    .Y(net4786));
 BUFx6f_ASAP7_75t_R place4787 (.A(_09115_),
    .Y(net4787));
 BUFx3_ASAP7_75t_R place4788 (.A(_09077_),
    .Y(net4788));
 BUFx3_ASAP7_75t_R place4789 (.A(_08340_),
    .Y(net4789));
 BUFx3_ASAP7_75t_R place4790 (.A(_08124_),
    .Y(net4790));
 BUFx3_ASAP7_75t_R place4791 (.A(_08124_),
    .Y(net4791));
 BUFx3_ASAP7_75t_R place4792 (.A(_08113_),
    .Y(net4792));
 BUFx3_ASAP7_75t_R place4793 (.A(_01374_),
    .Y(net4793));
 BUFx6f_ASAP7_75t_R place4794 (.A(net4795),
    .Y(net4794));
 BUFx3_ASAP7_75t_R place4795 (.A(_01372_),
    .Y(net4795));
 BUFx3_ASAP7_75t_R place4796 (.A(_01370_),
    .Y(net4796));
 BUFx3_ASAP7_75t_R place4797 (.A(net4798),
    .Y(net4797));
 BUFx3_ASAP7_75t_R place4798 (.A(_01367_),
    .Y(net4798));
 BUFx3_ASAP7_75t_R place4799 (.A(_01332_),
    .Y(net4799));
 BUFx6f_ASAP7_75t_R place4800 (.A(_01330_),
    .Y(net4800));
 BUFx3_ASAP7_75t_R place4801 (.A(_01328_),
    .Y(net4801));
 BUFx3_ASAP7_75t_R place4802 (.A(_01327_),
    .Y(net4802));
 BUFx3_ASAP7_75t_R place4803 (.A(_01325_),
    .Y(net4803));
 BUFx3_ASAP7_75t_R place4804 (.A(net4805),
    .Y(net4804));
 BUFx3_ASAP7_75t_R place4805 (.A(_01236_),
    .Y(net4805));
 BUFx3_ASAP7_75t_R place4806 (.A(_01235_),
    .Y(net4806));
 BUFx3_ASAP7_75t_R place4807 (.A(_01233_),
    .Y(net4807));
 BUFx3_ASAP7_75t_R place4808 (.A(_01233_),
    .Y(net4808));
 BUFx3_ASAP7_75t_R place4809 (.A(_01231_),
    .Y(net4809));
 BUFx3_ASAP7_75t_R place4810 (.A(_07475_),
    .Y(net4810));
 BUFx3_ASAP7_75t_R place4811 (.A(_07458_),
    .Y(net4811));
 BUFx3_ASAP7_75t_R place4812 (.A(_07458_),
    .Y(net4812));
 BUFx3_ASAP7_75t_R place4813 (.A(_07428_),
    .Y(net4813));
 BUFx3_ASAP7_75t_R place4814 (.A(_07409_),
    .Y(net4814));
 BUFx3_ASAP7_75t_R place4815 (.A(_07358_),
    .Y(net4815));
 BUFx3_ASAP7_75t_R place4816 (.A(net4817),
    .Y(net4816));
 BUFx6f_ASAP7_75t_R place4817 (.A(_07331_),
    .Y(net4817));
 BUFx3_ASAP7_75t_R place4818 (.A(_07304_),
    .Y(net4818));
 BUFx3_ASAP7_75t_R place4819 (.A(_07264_),
    .Y(net4819));
 BUFx3_ASAP7_75t_R place4820 (.A(_07261_),
    .Y(net4820));
 BUFx3_ASAP7_75t_R place4821 (.A(_07204_),
    .Y(net4821));
 BUFx6f_ASAP7_75t_R place4822 (.A(_06693_),
    .Y(net4822));
 BUFx3_ASAP7_75t_R place4823 (.A(_06618_),
    .Y(net4823));
 BUFx3_ASAP7_75t_R place4824 (.A(_06587_),
    .Y(net4824));
 BUFx3_ASAP7_75t_R place4825 (.A(_06568_),
    .Y(net4825));
 BUFx6f_ASAP7_75t_R place4826 (.A(_06568_),
    .Y(net4826));
 BUFx3_ASAP7_75t_R place4827 (.A(_06567_),
    .Y(net4827));
 BUFx3_ASAP7_75t_R place4828 (.A(net4829),
    .Y(net4828));
 BUFx3_ASAP7_75t_R place4829 (.A(_06142_),
    .Y(net4829));
 BUFx3_ASAP7_75t_R place4830 (.A(_06142_),
    .Y(net4830));
 BUFx3_ASAP7_75t_R place4831 (.A(_06103_),
    .Y(net4831));
 BUFx6f_ASAP7_75t_R place4832 (.A(_05991_),
    .Y(net4832));
 BUFx6f_ASAP7_75t_R place4833 (.A(_05984_),
    .Y(net4833));
 BUFx3_ASAP7_75t_R place4834 (.A(_05938_),
    .Y(net4834));
 BUFx3_ASAP7_75t_R place4835 (.A(_05928_),
    .Y(net4835));
 BUFx3_ASAP7_75t_R place4836 (.A(_05928_),
    .Y(net4836));
 BUFx6f_ASAP7_75t_R place4837 (.A(_05928_),
    .Y(net4837));
 BUFx3_ASAP7_75t_R place4838 (.A(_05911_),
    .Y(net4838));
 BUFx3_ASAP7_75t_R place4839 (.A(_05893_),
    .Y(net4839));
 BUFx3_ASAP7_75t_R place4840 (.A(_05403_),
    .Y(net4840));
 BUFx6f_ASAP7_75t_R place4841 (.A(net4842),
    .Y(net4841));
 BUFx3_ASAP7_75t_R place4842 (.A(_05379_),
    .Y(net4842));
 BUFx3_ASAP7_75t_R place4843 (.A(_05379_),
    .Y(net4843));
 BUFx3_ASAP7_75t_R place4844 (.A(_05363_),
    .Y(net4844));
 BUFx3_ASAP7_75t_R place4845 (.A(_05225_),
    .Y(net4845));
 BUFx3_ASAP7_75t_R place4846 (.A(_05225_),
    .Y(net4846));
 BUFx3_ASAP7_75t_R place4847 (.A(_05206_),
    .Y(net4847));
 BUFx3_ASAP7_75t_R place4848 (.A(_05203_),
    .Y(net4848));
 BUFx3_ASAP7_75t_R place4849 (.A(_04669_),
    .Y(net4849));
 BUFx3_ASAP7_75t_R place4850 (.A(_04640_),
    .Y(net4850));
 BUFx3_ASAP7_75t_R place4851 (.A(net4852),
    .Y(net4851));
 BUFx3_ASAP7_75t_R place4852 (.A(_04627_),
    .Y(net4852));
 BUFx6f_ASAP7_75t_R place4853 (.A(_04610_),
    .Y(net4853));
 BUFx3_ASAP7_75t_R place4854 (.A(_04610_),
    .Y(net4854));
 BUFx3_ASAP7_75t_R place4855 (.A(_04606_),
    .Y(net4855));
 BUFx6f_ASAP7_75t_R place4856 (.A(_04584_),
    .Y(net4856));
 BUFx3_ASAP7_75t_R place4857 (.A(_04565_),
    .Y(net4857));
 BUFx6f_ASAP7_75t_R place4858 (.A(_04556_),
    .Y(net4858));
 BUFx3_ASAP7_75t_R place4859 (.A(_04552_),
    .Y(net4859));
 BUFx3_ASAP7_75t_R place4860 (.A(_04546_),
    .Y(net4860));
 BUFx3_ASAP7_75t_R place4861 (.A(_04542_),
    .Y(net4861));
 BUFx6f_ASAP7_75t_R place4862 (.A(_04483_),
    .Y(net4862));
 BUFx3_ASAP7_75t_R place4863 (.A(_04483_),
    .Y(net4863));
 BUFx3_ASAP7_75t_R place4864 (.A(_04481_),
    .Y(net4864));
 BUFx3_ASAP7_75t_R place4865 (.A(_03877_),
    .Y(net4865));
 BUFx3_ASAP7_75t_R place4866 (.A(_03840_),
    .Y(net4866));
 BUFx3_ASAP7_75t_R place4867 (.A(_03838_),
    .Y(net4867));
 BUFx3_ASAP7_75t_R place4868 (.A(_03802_),
    .Y(net4868));
 BUFx3_ASAP7_75t_R place4869 (.A(_03793_),
    .Y(net4869));
 BUFx3_ASAP7_75t_R place4870 (.A(_03793_),
    .Y(net4870));
 BUFx3_ASAP7_75t_R place4871 (.A(_03759_),
    .Y(net4871));
 BUFx3_ASAP7_75t_R place4872 (.A(_03739_),
    .Y(net4872));
 BUFx3_ASAP7_75t_R place4873 (.A(_03459_),
    .Y(net4873));
 BUFx3_ASAP7_75t_R place4874 (.A(_03358_),
    .Y(net4874));
 BUFx3_ASAP7_75t_R place4875 (.A(_03178_),
    .Y(net4875));
 BUFx3_ASAP7_75t_R place4876 (.A(_03154_),
    .Y(net4876));
 BUFx3_ASAP7_75t_R place4877 (.A(_03137_),
    .Y(net4877));
 BUFx3_ASAP7_75t_R place4878 (.A(_03112_),
    .Y(net4878));
 BUFx3_ASAP7_75t_R place4879 (.A(_02600_),
    .Y(net4879));
 BUFx6f_ASAP7_75t_R place4880 (.A(_02536_),
    .Y(net4880));
 BUFx6f_ASAP7_75t_R place4881 (.A(_02471_),
    .Y(net4881));
 BUFx3_ASAP7_75t_R place4882 (.A(_02453_),
    .Y(net4882));
 BUFx3_ASAP7_75t_R place4883 (.A(_02453_),
    .Y(net4883));
 BUFx3_ASAP7_75t_R place4884 (.A(_02445_),
    .Y(net4884));
 BUFx3_ASAP7_75t_R place4885 (.A(_02430_),
    .Y(net4885));
 BUFx3_ASAP7_75t_R place4886 (.A(_02122_),
    .Y(net4886));
 BUFx3_ASAP7_75t_R place4887 (.A(_01956_),
    .Y(net4887));
 BUFx3_ASAP7_75t_R place4888 (.A(_01945_),
    .Y(net4888));
 BUFx3_ASAP7_75t_R place4889 (.A(_01925_),
    .Y(net4889));
 BUFx6f_ASAP7_75t_R place4890 (.A(_01824_),
    .Y(net4890));
 BUFx3_ASAP7_75t_R place4891 (.A(net4892),
    .Y(net4891));
 BUFx3_ASAP7_75t_R place4892 (.A(_01764_),
    .Y(net4892));
 BUFx3_ASAP7_75t_R place4893 (.A(_01764_),
    .Y(net4893));
 BUFx3_ASAP7_75t_R place4894 (.A(_01715_),
    .Y(net4894));
 BUFx3_ASAP7_75t_R place4895 (.A(_01706_),
    .Y(net4895));
 BUFx3_ASAP7_75t_R place4896 (.A(_01688_),
    .Y(net4896));
 BUFx3_ASAP7_75t_R place4897 (.A(_01679_),
    .Y(net4897));
 BUFx3_ASAP7_75t_R place4898 (.A(_15307_),
    .Y(net4898));
 BUFx3_ASAP7_75t_R place4899 (.A(_15197_),
    .Y(net4899));
 BUFx6f_ASAP7_75t_R place4900 (.A(_15174_),
    .Y(net4900));
 BUFx3_ASAP7_75t_R place4901 (.A(_15164_),
    .Y(net4901));
 BUFx3_ASAP7_75t_R place4902 (.A(_15093_),
    .Y(net4902));
 BUFx3_ASAP7_75t_R place4903 (.A(_15068_),
    .Y(net4903));
 BUFx3_ASAP7_75t_R place4904 (.A(_14993_),
    .Y(net4904));
 BUFx3_ASAP7_75t_R place4905 (.A(_14589_),
    .Y(net4905));
 BUFx3_ASAP7_75t_R place4906 (.A(_14528_),
    .Y(net4906));
 BUFx3_ASAP7_75t_R place4907 (.A(_14501_),
    .Y(net4907));
 BUFx3_ASAP7_75t_R place4908 (.A(_14453_),
    .Y(net4908));
 BUFx3_ASAP7_75t_R place4909 (.A(_14441_),
    .Y(net4909));
 BUFx3_ASAP7_75t_R place4910 (.A(_14405_),
    .Y(net4910));
 BUFx3_ASAP7_75t_R place4911 (.A(_14401_),
    .Y(net4911));
 BUFx3_ASAP7_75t_R place4912 (.A(_14399_),
    .Y(net4912));
 BUFx3_ASAP7_75t_R place4913 (.A(_14386_),
    .Y(net4913));
 BUFx3_ASAP7_75t_R place4914 (.A(_14347_),
    .Y(net4914));
 BUFx3_ASAP7_75t_R place4915 (.A(_14113_),
    .Y(net4915));
 BUFx3_ASAP7_75t_R place4916 (.A(_13983_),
    .Y(net4916));
 BUFx3_ASAP7_75t_R place4917 (.A(_13908_),
    .Y(net4917));
 BUFx3_ASAP7_75t_R place4918 (.A(_13908_),
    .Y(net4918));
 BUFx3_ASAP7_75t_R place4919 (.A(_13822_),
    .Y(net4919));
 BUFx3_ASAP7_75t_R place4920 (.A(_13735_),
    .Y(net4920));
 BUFx3_ASAP7_75t_R place4921 (.A(_13701_),
    .Y(net4921));
 BUFx3_ASAP7_75t_R place4922 (.A(_13682_),
    .Y(net4922));
 BUFx3_ASAP7_75t_R place4923 (.A(net4924),
    .Y(net4923));
 BUFx6f_ASAP7_75t_R place4924 (.A(_13682_),
    .Y(net4924));
 BUFx3_ASAP7_75t_R place4925 (.A(_13648_),
    .Y(net4925));
 BUFx3_ASAP7_75t_R place4926 (.A(_13641_),
    .Y(net4926));
 BUFx3_ASAP7_75t_R place4927 (.A(_13615_),
    .Y(net4927));
 BUFx3_ASAP7_75t_R place4928 (.A(_13598_),
    .Y(net4928));
 BUFx6f_ASAP7_75t_R place4929 (.A(_13366_),
    .Y(net4929));
 BUFx3_ASAP7_75t_R place4930 (.A(_13079_),
    .Y(net4930));
 BUFx3_ASAP7_75t_R place4931 (.A(_13055_),
    .Y(net4931));
 BUFx3_ASAP7_75t_R place4932 (.A(_12980_),
    .Y(net4932));
 BUFx3_ASAP7_75t_R place4933 (.A(_12973_),
    .Y(net4933));
 BUFx3_ASAP7_75t_R place4934 (.A(_12951_),
    .Y(net4934));
 BUFx6f_ASAP7_75t_R place4935 (.A(_12951_),
    .Y(net4935));
 BUFx3_ASAP7_75t_R place4936 (.A(_12939_),
    .Y(net4936));
 BUFx3_ASAP7_75t_R place4937 (.A(_12878_),
    .Y(net4937));
 BUFx3_ASAP7_75t_R place4938 (.A(_12470_),
    .Y(net4938));
 BUFx3_ASAP7_75t_R place4939 (.A(_12444_),
    .Y(net4939));
 BUFx6f_ASAP7_75t_R place4940 (.A(_12365_),
    .Y(net4940));
 BUFx3_ASAP7_75t_R place4941 (.A(_12359_),
    .Y(net4941));
 BUFx3_ASAP7_75t_R place4942 (.A(_12335_),
    .Y(net4942));
 BUFx3_ASAP7_75t_R place4943 (.A(_12330_),
    .Y(net4943));
 BUFx3_ASAP7_75t_R place4944 (.A(_12304_),
    .Y(net4944));
 BUFx3_ASAP7_75t_R place4945 (.A(_12294_),
    .Y(net4945));
 BUFx3_ASAP7_75t_R place4946 (.A(_12286_),
    .Y(net4946));
 BUFx3_ASAP7_75t_R place4947 (.A(_12264_),
    .Y(net4947));
 BUFx3_ASAP7_75t_R place4948 (.A(_11675_),
    .Y(net4948));
 BUFx3_ASAP7_75t_R place4949 (.A(_11654_),
    .Y(net4949));
 BUFx3_ASAP7_75t_R place4950 (.A(_11603_),
    .Y(net4950));
 BUFx3_ASAP7_75t_R place4951 (.A(_11588_),
    .Y(net4951));
 BUFx3_ASAP7_75t_R place4952 (.A(_11541_),
    .Y(net4952));
 BUFx3_ASAP7_75t_R place4953 (.A(_11497_),
    .Y(net4953));
 BUFx3_ASAP7_75t_R place4954 (.A(_11160_),
    .Y(net4954));
 BUFx3_ASAP7_75t_R place4955 (.A(_11046_),
    .Y(net4955));
 BUFx3_ASAP7_75t_R place4956 (.A(_10986_),
    .Y(net4956));
 BUFx3_ASAP7_75t_R place4957 (.A(_10961_),
    .Y(net4957));
 BUFx3_ASAP7_75t_R place4958 (.A(_10935_),
    .Y(net4958));
 BUFx3_ASAP7_75t_R place4959 (.A(_10897_),
    .Y(net4959));
 BUFx3_ASAP7_75t_R place4960 (.A(_10879_),
    .Y(net4960));
 BUFx3_ASAP7_75t_R place4961 (.A(_10213_),
    .Y(net4961));
 BUFx3_ASAP7_75t_R place4962 (.A(_10158_),
    .Y(net4962));
 BUFx3_ASAP7_75t_R place4963 (.A(_10130_),
    .Y(net4963));
 BUFx3_ASAP7_75t_R place4964 (.A(_10122_),
    .Y(net4964));
 BUFx3_ASAP7_75t_R place4965 (.A(_10119_),
    .Y(net4965));
 BUFx3_ASAP7_75t_R place4966 (.A(_09862_),
    .Y(net4966));
 BUFx3_ASAP7_75t_R place4967 (.A(_09705_),
    .Y(net4967));
 BUFx3_ASAP7_75t_R place4968 (.A(_09686_),
    .Y(net4968));
 BUFx3_ASAP7_75t_R place4969 (.A(_09626_),
    .Y(net4969));
 BUFx3_ASAP7_75t_R place4970 (.A(_09264_),
    .Y(net4970));
 BUFx3_ASAP7_75t_R place4971 (.A(_09251_),
    .Y(net4971));
 BUFx3_ASAP7_75t_R place4972 (.A(_09180_),
    .Y(net4972));
 BUFx3_ASAP7_75t_R place4973 (.A(_09159_),
    .Y(net4973));
 BUFx3_ASAP7_75t_R place4974 (.A(_09135_),
    .Y(net4974));
 BUFx3_ASAP7_75t_R place4975 (.A(_09100_),
    .Y(net4975));
 BUFx3_ASAP7_75t_R place4976 (.A(_09089_),
    .Y(net4976));
 BUFx3_ASAP7_75t_R place4977 (.A(_09065_),
    .Y(net4977));
 BUFx3_ASAP7_75t_R place4978 (.A(_08390_),
    .Y(net4978));
 BUFx3_ASAP7_75t_R place4979 (.A(_08353_),
    .Y(net4979));
 BUFx3_ASAP7_75t_R place4980 (.A(_08289_),
    .Y(net4980));
 BUFx3_ASAP7_75t_R place4981 (.A(_08226_),
    .Y(net4981));
 BUFx6f_ASAP7_75t_R place4982 (.A(_08176_),
    .Y(net4982));
 BUFx3_ASAP7_75t_R place4983 (.A(_08116_),
    .Y(net4983));
 BUFx3_ASAP7_75t_R place4984 (.A(_08105_),
    .Y(net4984));
 BUFx3_ASAP7_75t_R place4985 (.A(_08100_),
    .Y(net4985));
 BUFx3_ASAP7_75t_R place4986 (.A(net4987),
    .Y(net4986));
 BUFx3_ASAP7_75t_R place4987 (.A(_01278_),
    .Y(net4987));
 BUFx3_ASAP7_75t_R place4988 (.A(_01148_),
    .Y(net4988));
 BUFx3_ASAP7_75t_R place4989 (.A(net4990),
    .Y(net4989));
 BUFx3_ASAP7_75t_R place4990 (.A(_01127_),
    .Y(net4990));
 BUFx3_ASAP7_75t_R place4991 (.A(_01106_),
    .Y(net4991));
 BUFx3_ASAP7_75t_R place4992 (.A(_07310_),
    .Y(net4992));
 BUFx3_ASAP7_75t_R place4993 (.A(_05966_),
    .Y(net4993));
 BUFx3_ASAP7_75t_R place4994 (.A(_05895_),
    .Y(net4994));
 BUFx3_ASAP7_75t_R place4995 (.A(_05809_),
    .Y(net4995));
 BUFx3_ASAP7_75t_R place4996 (.A(_01766_),
    .Y(net4996));
 BUFx6f_ASAP7_75t_R place4997 (.A(_01766_),
    .Y(net4997));
 BUFx3_ASAP7_75t_R place4998 (.A(_01766_),
    .Y(net4998));
 BUFx3_ASAP7_75t_R place4999 (.A(_01744_),
    .Y(net4999));
 BUFx3_ASAP7_75t_R place5000 (.A(_01744_),
    .Y(net5000));
 BUFx6f_ASAP7_75t_R place5001 (.A(net5002),
    .Y(net5001));
 BUFx6f_ASAP7_75t_R place5002 (.A(_15231_),
    .Y(net5002));
 BUFx3_ASAP7_75t_R place5003 (.A(_15099_),
    .Y(net5003));
 BUFx3_ASAP7_75t_R place5004 (.A(_15034_),
    .Y(net5004));
 BUFx3_ASAP7_75t_R place5005 (.A(_14476_),
    .Y(net5005));
 BUFx6f_ASAP7_75t_R place5006 (.A(_14474_),
    .Y(net5006));
 BUFx3_ASAP7_75t_R place5007 (.A(_14474_),
    .Y(net5007));
 BUFx3_ASAP7_75t_R place5008 (.A(_14449_),
    .Y(net5008));
 BUFx3_ASAP7_75t_R place5009 (.A(_11617_),
    .Y(net5009));
 BUFx3_ASAP7_75t_R place5010 (.A(net5011),
    .Y(net5010));
 BUFx6f_ASAP7_75t_R place5011 (.A(_11557_),
    .Y(net5011));
 BUFx3_ASAP7_75t_R place5012 (.A(_10912_),
    .Y(net5012));
 BUFx3_ASAP7_75t_R place5013 (.A(_10912_),
    .Y(net5013));
 BUFx3_ASAP7_75t_R place5014 (.A(net5015),
    .Y(net5014));
 BUFx3_ASAP7_75t_R place5015 (.A(_10901_),
    .Y(net5015));
 BUFx6f_ASAP7_75t_R place5016 (.A(_10849_),
    .Y(net5016));
 BUFx3_ASAP7_75t_R place5017 (.A(_10226_),
    .Y(net5017));
 BUFx3_ASAP7_75t_R place5018 (.A(_10209_),
    .Y(net5018));
 BUFx3_ASAP7_75t_R place5019 (.A(_10209_),
    .Y(net5019));
 BUFx3_ASAP7_75t_R place5020 (.A(_09692_),
    .Y(net5020));
 BUFx6f_ASAP7_75t_R place5021 (.A(_09680_),
    .Y(net5021));
 BUFx3_ASAP7_75t_R place5022 (.A(net5023),
    .Y(net5022));
 BUFx3_ASAP7_75t_R place5023 (.A(_09604_),
    .Y(net5023));
 BUFx3_ASAP7_75t_R place5024 (.A(_09127_),
    .Y(net5024));
 BUFx6f_ASAP7_75t_R place5025 (.A(_09127_),
    .Y(net5025));
 BUFx3_ASAP7_75t_R place5026 (.A(_09127_),
    .Y(net5026));
 BUFx3_ASAP7_75t_R place5027 (.A(_09035_),
    .Y(net5027));
 BUFx3_ASAP7_75t_R place5028 (.A(_08266_),
    .Y(net5028));
 BUFx3_ASAP7_75t_R place5029 (.A(_08112_),
    .Y(net5029));
 BUFx3_ASAP7_75t_R place5030 (.A(_01391_),
    .Y(net5030));
 BUFx3_ASAP7_75t_R place5031 (.A(_01391_),
    .Y(net5031));
 BUFx3_ASAP7_75t_R place5032 (.A(_01310_),
    .Y(net5032));
 BUFx3_ASAP7_75t_R place5033 (.A(_01309_),
    .Y(net5033));
 BUFx3_ASAP7_75t_R place5034 (.A(_01308_),
    .Y(net5034));
 BUFx3_ASAP7_75t_R place5035 (.A(net5036),
    .Y(net5035));
 BUFx3_ASAP7_75t_R place5036 (.A(_01307_),
    .Y(net5036));
 BUFx3_ASAP7_75t_R place5037 (.A(_01305_),
    .Y(net5037));
 BUFx3_ASAP7_75t_R place5038 (.A(_01304_),
    .Y(net5038));
 BUFx3_ASAP7_75t_R place5039 (.A(_01302_),
    .Y(net5039));
 BUFx3_ASAP7_75t_R place5040 (.A(net5041),
    .Y(net5040));
 BUFx3_ASAP7_75t_R place5041 (.A(_01287_),
    .Y(net5041));
 BUFx3_ASAP7_75t_R place5042 (.A(_01286_),
    .Y(net5042));
 BUFx3_ASAP7_75t_R place5043 (.A(_01285_),
    .Y(net5043));
 BUFx3_ASAP7_75t_R place5044 (.A(net5045),
    .Y(net5044));
 BUFx3_ASAP7_75t_R place5045 (.A(_01285_),
    .Y(net5045));
 BUFx3_ASAP7_75t_R place5046 (.A(_01284_),
    .Y(net5046));
 BUFx3_ASAP7_75t_R place5047 (.A(_01282_),
    .Y(net5047));
 BUFx3_ASAP7_75t_R place5048 (.A(_01281_),
    .Y(net5048));
 BUFx3_ASAP7_75t_R place5049 (.A(_01264_),
    .Y(net5049));
 BUFx3_ASAP7_75t_R place5050 (.A(_01263_),
    .Y(net5050));
 BUFx3_ASAP7_75t_R place5051 (.A(_01262_),
    .Y(net5051));
 BUFx3_ASAP7_75t_R place5052 (.A(_01262_),
    .Y(net5052));
 BUFx3_ASAP7_75t_R place5053 (.A(_01261_),
    .Y(net5053));
 BUFx3_ASAP7_75t_R place5054 (.A(_01259_),
    .Y(net5054));
 BUFx3_ASAP7_75t_R place5055 (.A(_01258_),
    .Y(net5055));
 BUFx3_ASAP7_75t_R place5056 (.A(_01256_),
    .Y(net5056));
 BUFx3_ASAP7_75t_R place5057 (.A(_01254_),
    .Y(net5057));
 BUFx3_ASAP7_75t_R place5058 (.A(_01241_),
    .Y(net5058));
 BUFx3_ASAP7_75t_R place5059 (.A(_01240_),
    .Y(net5059));
 BUFx3_ASAP7_75t_R place5060 (.A(_01239_),
    .Y(net5060));
 BUFx3_ASAP7_75t_R place5061 (.A(_01198_),
    .Y(net5061));
 BUFx3_ASAP7_75t_R place5062 (.A(_01196_),
    .Y(net5062));
 BUFx3_ASAP7_75t_R place5063 (.A(_01195_),
    .Y(net5063));
 BUFx3_ASAP7_75t_R place5064 (.A(_01151_),
    .Y(net5064));
 BUFx3_ASAP7_75t_R place5065 (.A(_01149_),
    .Y(net5065));
 BUFx3_ASAP7_75t_R place5066 (.A(net5067),
    .Y(net5066));
 BUFx3_ASAP7_75t_R place5067 (.A(_01133_),
    .Y(net5067));
 BUFx3_ASAP7_75t_R place5068 (.A(_01132_),
    .Y(net5068));
 BUFx3_ASAP7_75t_R place5069 (.A(_01128_),
    .Y(net5069));
 BUFx3_ASAP7_75t_R place5070 (.A(_01112_),
    .Y(net5070));
 BUFx3_ASAP7_75t_R place5071 (.A(_01107_),
    .Y(net5071));
 BUFx3_ASAP7_75t_R place5072 (.A(_01105_),
    .Y(net5072));
 BUFx3_ASAP7_75t_R place5073 (.A(_07474_),
    .Y(net5073));
 BUFx3_ASAP7_75t_R place5074 (.A(_07322_),
    .Y(net5074));
 BUFx3_ASAP7_75t_R place5075 (.A(_07230_),
    .Y(net5075));
 BUFx3_ASAP7_75t_R place5076 (.A(_07227_),
    .Y(net5076));
 BUFx3_ASAP7_75t_R place5077 (.A(_07174_),
    .Y(net5077));
 BUFx3_ASAP7_75t_R place5078 (.A(_07170_),
    .Y(net5078));
 BUFx3_ASAP7_75t_R place5079 (.A(net5081),
    .Y(net5079));
 BUFx3_ASAP7_75t_R place5080 (.A(net5081),
    .Y(net5080));
 BUFx3_ASAP7_75t_R place5081 (.A(_06492_),
    .Y(net5081));
 BUFx3_ASAP7_75t_R place5082 (.A(_06472_),
    .Y(net5082));
 BUFx3_ASAP7_75t_R place5083 (.A(_06472_),
    .Y(net5083));
 BUFx3_ASAP7_75t_R place5084 (.A(_06229_),
    .Y(net5084));
 BUFx3_ASAP7_75t_R place5085 (.A(_06141_),
    .Y(net5085));
 BUFx3_ASAP7_75t_R place5086 (.A(_06071_),
    .Y(net5086));
 BUFx3_ASAP7_75t_R place5087 (.A(_06009_),
    .Y(net5087));
 BUFx3_ASAP7_75t_R place5088 (.A(net5089),
    .Y(net5088));
 BUFx6f_ASAP7_75t_R place5089 (.A(_06009_),
    .Y(net5089));
 BUFx3_ASAP7_75t_R place5090 (.A(_06002_),
    .Y(net5090));
 BUFx3_ASAP7_75t_R place5091 (.A(_05960_),
    .Y(net5091));
 BUFx3_ASAP7_75t_R place5092 (.A(_05927_),
    .Y(net5092));
 BUFx3_ASAP7_75t_R place5093 (.A(_05826_),
    .Y(net5093));
 BUFx6f_ASAP7_75t_R place5094 (.A(_05344_),
    .Y(net5094));
 BUFx3_ASAP7_75t_R place5095 (.A(net5096),
    .Y(net5095));
 BUFx3_ASAP7_75t_R place5096 (.A(_05123_),
    .Y(net5096));
 BUFx3_ASAP7_75t_R place5097 (.A(net5098),
    .Y(net5097));
 BUFx3_ASAP7_75t_R place5098 (.A(_05103_),
    .Y(net5098));
 BUFx3_ASAP7_75t_R place5099 (.A(_05103_),
    .Y(net5099));
 BUFx3_ASAP7_75t_R place5100 (.A(net5101),
    .Y(net5100));
 BUFx3_ASAP7_75t_R place5101 (.A(_04434_),
    .Y(net5101));
 BUFx6f_ASAP7_75t_R place5102 (.A(_04434_),
    .Y(net5102));
 BUFx6f_ASAP7_75t_R place5103 (.A(_04428_),
    .Y(net5103));
 BUFx3_ASAP7_75t_R place5104 (.A(_04428_),
    .Y(net5104));
 BUFx3_ASAP7_75t_R place5105 (.A(_03980_),
    .Y(net5105));
 BUFx3_ASAP7_75t_R place5106 (.A(_03980_),
    .Y(net5106));
 BUFx3_ASAP7_75t_R place5107 (.A(_03805_),
    .Y(net5107));
 BUFx3_ASAP7_75t_R place5108 (.A(_03800_),
    .Y(net5108));
 BUFx3_ASAP7_75t_R place5109 (.A(_03743_),
    .Y(net5109));
 BUFx3_ASAP7_75t_R place5110 (.A(_03036_),
    .Y(net5110));
 BUFx3_ASAP7_75t_R place5111 (.A(_03036_),
    .Y(net5111));
 BUFx3_ASAP7_75t_R place5112 (.A(_02429_),
    .Y(net5112));
 BUFx3_ASAP7_75t_R place5113 (.A(net5114),
    .Y(net5113));
 BUFx3_ASAP7_75t_R place5114 (.A(_02387_),
    .Y(net5114));
 BUFx3_ASAP7_75t_R place5115 (.A(_02191_),
    .Y(net5115));
 BUFx3_ASAP7_75t_R place5116 (.A(_01924_),
    .Y(net5116));
 BUFx6f_ASAP7_75t_R place5117 (.A(_01918_),
    .Y(net5117));
 BUFx3_ASAP7_75t_R place5118 (.A(_01918_),
    .Y(net5118));
 BUFx3_ASAP7_75t_R place5119 (.A(_01896_),
    .Y(net5119));
 BUFx3_ASAP7_75t_R place5120 (.A(_01869_),
    .Y(net5120));
 BUFx3_ASAP7_75t_R place5121 (.A(_01853_),
    .Y(net5121));
 BUFx3_ASAP7_75t_R place5122 (.A(_01841_),
    .Y(net5122));
 BUFx3_ASAP7_75t_R place5123 (.A(_01834_),
    .Y(net5123));
 BUFx6f_ASAP7_75t_R place5124 (.A(_01759_),
    .Y(net5124));
 BUFx3_ASAP7_75t_R place5125 (.A(_01756_),
    .Y(net5125));
 BUFx3_ASAP7_75t_R place5126 (.A(_01747_),
    .Y(net5126));
 BUFx3_ASAP7_75t_R place5127 (.A(_01708_),
    .Y(net5127));
 BUFx3_ASAP7_75t_R place5128 (.A(_01705_),
    .Y(net5128));
 BUFx3_ASAP7_75t_R place5129 (.A(net5130),
    .Y(net5129));
 BUFx3_ASAP7_75t_R place5130 (.A(_01687_),
    .Y(net5130));
 BUFx3_ASAP7_75t_R place5131 (.A(_01678_),
    .Y(net5131));
 BUFx6f_ASAP7_75t_R place5132 (.A(_01671_),
    .Y(net5132));
 BUFx3_ASAP7_75t_R place5133 (.A(_15306_),
    .Y(net5133));
 BUFx6f_ASAP7_75t_R place5134 (.A(_15255_),
    .Y(net5134));
 BUFx3_ASAP7_75t_R place5135 (.A(_15214_),
    .Y(net5135));
 BUFx3_ASAP7_75t_R place5136 (.A(_15210_),
    .Y(net5136));
 BUFx6f_ASAP7_75t_R place5137 (.A(_15205_),
    .Y(net5137));
 BUFx3_ASAP7_75t_R place5138 (.A(_15190_),
    .Y(net5138));
 BUFx3_ASAP7_75t_R place5139 (.A(_15190_),
    .Y(net5139));
 BUFx6f_ASAP7_75t_R place5140 (.A(_15187_),
    .Y(net5140));
 BUFx3_ASAP7_75t_R place5141 (.A(_15187_),
    .Y(net5141));
 BUFx3_ASAP7_75t_R place5142 (.A(_15173_),
    .Y(net5142));
 BUFx6f_ASAP7_75t_R place5143 (.A(_15162_),
    .Y(net5143));
 BUFx3_ASAP7_75t_R place5144 (.A(_15121_),
    .Y(net5144));
 BUFx6f_ASAP7_75t_R place5145 (.A(_15121_),
    .Y(net5145));
 BUFx3_ASAP7_75t_R place5146 (.A(_15061_),
    .Y(net5146));
 BUFx3_ASAP7_75t_R place5147 (.A(_15061_),
    .Y(net5147));
 BUFx3_ASAP7_75t_R place5148 (.A(_15037_),
    .Y(net5148));
 BUFx3_ASAP7_75t_R place5149 (.A(net5151),
    .Y(net5149));
 BUFx3_ASAP7_75t_R place5150 (.A(net5151),
    .Y(net5150));
 BUFx6f_ASAP7_75t_R place5151 (.A(_15037_),
    .Y(net5151));
 BUFx3_ASAP7_75t_R place5152 (.A(net5154),
    .Y(net5152));
 BUFx3_ASAP7_75t_R place5153 (.A(net5154),
    .Y(net5153));
 BUFx6f_ASAP7_75t_R place5154 (.A(_15037_),
    .Y(net5154));
 BUFx3_ASAP7_75t_R place5155 (.A(_15037_),
    .Y(net5155));
 BUFx3_ASAP7_75t_R place5156 (.A(_14992_),
    .Y(net5156));
 BUFx3_ASAP7_75t_R place5157 (.A(net5158),
    .Y(net5157));
 BUFx6f_ASAP7_75t_R place5158 (.A(_14975_),
    .Y(net5158));
 BUFx3_ASAP7_75t_R place5159 (.A(_14774_),
    .Y(net5159));
 BUFx3_ASAP7_75t_R place5160 (.A(_14632_),
    .Y(net5160));
 BUFx3_ASAP7_75t_R place5161 (.A(_14580_),
    .Y(net5161));
 BUFx3_ASAP7_75t_R place5162 (.A(_14440_),
    .Y(net5162));
 BUFx3_ASAP7_75t_R place5163 (.A(net5164),
    .Y(net5163));
 BUFx3_ASAP7_75t_R place5164 (.A(_14404_),
    .Y(net5164));
 BUFx3_ASAP7_75t_R place5165 (.A(_14385_),
    .Y(net5165));
 BUFx3_ASAP7_75t_R place5166 (.A(_14380_),
    .Y(net5166));
 BUFx3_ASAP7_75t_R place5167 (.A(_14311_),
    .Y(net5167));
 BUFx3_ASAP7_75t_R place5168 (.A(_14270_),
    .Y(net5168));
 BUFx3_ASAP7_75t_R place5169 (.A(_13907_),
    .Y(net5169));
 BUFx3_ASAP7_75t_R place5170 (.A(_13906_),
    .Y(net5170));
 BUFx3_ASAP7_75t_R place5171 (.A(_13876_),
    .Y(net5171));
 BUFx3_ASAP7_75t_R place5172 (.A(net5173),
    .Y(net5172));
 BUFx3_ASAP7_75t_R place5173 (.A(_13842_),
    .Y(net5173));
 BUFx3_ASAP7_75t_R place5174 (.A(_13805_),
    .Y(net5174));
 BUFx3_ASAP7_75t_R place5175 (.A(_13792_),
    .Y(net5175));
 BUFx3_ASAP7_75t_R place5176 (.A(_13768_),
    .Y(net5176));
 BUFx6f_ASAP7_75t_R place5177 (.A(_13764_),
    .Y(net5177));
 BUFx3_ASAP7_75t_R place5178 (.A(_13731_),
    .Y(net5178));
 BUFx6f_ASAP7_75t_R place5179 (.A(_13712_),
    .Y(net5179));
 BUFx3_ASAP7_75t_R place5180 (.A(_13692_),
    .Y(net5180));
 BUFx3_ASAP7_75t_R place5181 (.A(_13686_),
    .Y(net5181));
 BUFx3_ASAP7_75t_R place5182 (.A(_13635_),
    .Y(net5182));
 BUFx6f_ASAP7_75t_R place5183 (.A(net5184),
    .Y(net5183));
 BUFx3_ASAP7_75t_R place5184 (.A(_13597_),
    .Y(net5184));
 BUFx6f_ASAP7_75t_R place5185 (.A(_13053_),
    .Y(net5185));
 BUFx3_ASAP7_75t_R place5186 (.A(_13045_),
    .Y(net5186));
 BUFx3_ASAP7_75t_R place5187 (.A(_13015_),
    .Y(net5187));
 BUFx3_ASAP7_75t_R place5188 (.A(_12970_),
    .Y(net5188));
 BUFx3_ASAP7_75t_R place5189 (.A(_12945_),
    .Y(net5189));
 BUFx3_ASAP7_75t_R place5190 (.A(net5191),
    .Y(net5190));
 BUFx3_ASAP7_75t_R place5191 (.A(_12938_),
    .Y(net5191));
 BUFx3_ASAP7_75t_R place5192 (.A(_12475_),
    .Y(net5192));
 BUFx3_ASAP7_75t_R place5193 (.A(_12469_),
    .Y(net5193));
 BUFx3_ASAP7_75t_R place5194 (.A(_12428_),
    .Y(net5194));
 BUFx3_ASAP7_75t_R place5195 (.A(_12329_),
    .Y(net5195));
 BUFx3_ASAP7_75t_R place5196 (.A(_12313_),
    .Y(net5196));
 BUFx3_ASAP7_75t_R place5197 (.A(_12285_),
    .Y(net5197));
 BUFx3_ASAP7_75t_R place5198 (.A(_12262_),
    .Y(net5198));
 BUFx3_ASAP7_75t_R place5199 (.A(_11795_),
    .Y(net5199));
 BUFx3_ASAP7_75t_R place5200 (.A(_11792_),
    .Y(net5200));
 BUFx3_ASAP7_75t_R place5201 (.A(_11755_),
    .Y(net5201));
 BUFx3_ASAP7_75t_R place5202 (.A(_11678_),
    .Y(net5202));
 BUFx3_ASAP7_75t_R place5203 (.A(_11664_),
    .Y(net5203));
 BUFx3_ASAP7_75t_R place5204 (.A(_11606_),
    .Y(net5204));
 BUFx3_ASAP7_75t_R place5205 (.A(_11554_),
    .Y(net5205));
 BUFx6f_ASAP7_75t_R place5206 (.A(_11554_),
    .Y(net5206));
 BUFx3_ASAP7_75t_R place5207 (.A(_11549_),
    .Y(net5207));
 BUFx3_ASAP7_75t_R place5208 (.A(_11543_),
    .Y(net5208));
 BUFx3_ASAP7_75t_R place5209 (.A(_11101_),
    .Y(net5209));
 BUFx3_ASAP7_75t_R place5210 (.A(_11060_),
    .Y(net5210));
 BUFx3_ASAP7_75t_R place5211 (.A(_11045_),
    .Y(net5211));
 BUFx3_ASAP7_75t_R place5212 (.A(_10898_),
    .Y(net5212));
 BUFx3_ASAP7_75t_R place5213 (.A(_10882_),
    .Y(net5213));
 BUFx3_ASAP7_75t_R place5214 (.A(_10874_),
    .Y(net5214));
 BUFx3_ASAP7_75t_R place5215 (.A(_10871_),
    .Y(net5215));
 BUFx3_ASAP7_75t_R place5216 (.A(_10831_),
    .Y(net5216));
 BUFx3_ASAP7_75t_R place5217 (.A(_10831_),
    .Y(net5217));
 BUFx3_ASAP7_75t_R place5218 (.A(_10821_),
    .Y(net5218));
 BUFx3_ASAP7_75t_R place5219 (.A(_10814_),
    .Y(net5219));
 BUFx3_ASAP7_75t_R place5220 (.A(_10814_),
    .Y(net5220));
 BUFx3_ASAP7_75t_R place5221 (.A(_10814_),
    .Y(net5221));
 BUFx3_ASAP7_75t_R place5222 (.A(_10790_),
    .Y(net5222));
 BUFx3_ASAP7_75t_R place5223 (.A(_10239_),
    .Y(net5223));
 BUFx3_ASAP7_75t_R place5224 (.A(_10180_),
    .Y(net5224));
 BUFx3_ASAP7_75t_R place5225 (.A(_10143_),
    .Y(net5225));
 BUFx3_ASAP7_75t_R place5226 (.A(_10143_),
    .Y(net5226));
 BUFx3_ASAP7_75t_R place5227 (.A(net5228),
    .Y(net5227));
 BUFx3_ASAP7_75t_R place5228 (.A(_10118_),
    .Y(net5228));
 BUFx3_ASAP7_75t_R place5229 (.A(_09723_),
    .Y(net5229));
 BUFx3_ASAP7_75t_R place5230 (.A(_09703_),
    .Y(net5230));
 BUFx3_ASAP7_75t_R place5231 (.A(_09643_),
    .Y(net5231));
 BUFx3_ASAP7_75t_R place5232 (.A(_09635_),
    .Y(net5232));
 BUFx6f_ASAP7_75t_R place5233 (.A(_09609_),
    .Y(net5233));
 BUFx3_ASAP7_75t_R place5234 (.A(_09602_),
    .Y(net5234));
 BUFx3_ASAP7_75t_R place5235 (.A(_09256_),
    .Y(net5235));
 BUFx6f_ASAP7_75t_R place5236 (.A(_09156_),
    .Y(net5236));
 BUFx3_ASAP7_75t_R place5237 (.A(_09145_),
    .Y(net5237));
 BUFx6f_ASAP7_75t_R place5238 (.A(_09105_),
    .Y(net5238));
 BUFx3_ASAP7_75t_R place5239 (.A(_09094_),
    .Y(net5239));
 BUFx3_ASAP7_75t_R place5240 (.A(_09092_),
    .Y(net5240));
 BUFx3_ASAP7_75t_R place5241 (.A(_09039_),
    .Y(net5241));
 BUFx3_ASAP7_75t_R place5242 (.A(_08397_),
    .Y(net5242));
 BUFx3_ASAP7_75t_R place5243 (.A(_08302_),
    .Y(net5243));
 BUFx3_ASAP7_75t_R place5244 (.A(net5245),
    .Y(net5244));
 BUFx6f_ASAP7_75t_R place5245 (.A(_08225_),
    .Y(net5245));
 BUFx3_ASAP7_75t_R place5246 (.A(_08185_),
    .Y(net5246));
 BUFx3_ASAP7_75t_R place5247 (.A(_08157_),
    .Y(net5247));
 BUFx3_ASAP7_75t_R place5248 (.A(_08151_),
    .Y(net5248));
 BUFx3_ASAP7_75t_R place5249 (.A(_08143_),
    .Y(net5249));
 BUFx6f_ASAP7_75t_R place5250 (.A(_08132_),
    .Y(net5250));
 BUFx3_ASAP7_75t_R place5251 (.A(_08115_),
    .Y(net5251));
 BUFx3_ASAP7_75t_R place5252 (.A(_08099_),
    .Y(net5252));
 BUFx3_ASAP7_75t_R place5253 (.A(_01345_),
    .Y(net5253));
 BUFx3_ASAP7_75t_R place5254 (.A(_01211_),
    .Y(net5254));
 BUFx3_ASAP7_75t_R place5255 (.A(_01190_),
    .Y(net5255));
 BUFx3_ASAP7_75t_R place5256 (.A(net5257),
    .Y(net5256));
 BUFx3_ASAP7_75t_R place5257 (.A(_01169_),
    .Y(net5257));
 BUFx3_ASAP7_75t_R place5258 (.A(_01085_),
    .Y(net5258));
 BUFx3_ASAP7_75t_R place5259 (.A(_01064_),
    .Y(net5259));
 BUFx3_ASAP7_75t_R place5260 (.A(_00998_),
    .Y(net5260));
 BUFx3_ASAP7_75t_R place5261 (.A(_00975_),
    .Y(net5261));
 BUFx6f_ASAP7_75t_R place5262 (.A(net5263),
    .Y(net5262));
 BUFx6f_ASAP7_75t_R place5263 (.A(_10173_),
    .Y(net5263));
 BUFx3_ASAP7_75t_R place5264 (.A(_10155_),
    .Y(net5264));
 BUFx3_ASAP7_75t_R place5265 (.A(_10147_),
    .Y(net5265));
 BUFx3_ASAP7_75t_R place5266 (.A(_09666_),
    .Y(net5266));
 BUFx3_ASAP7_75t_R place5267 (.A(_09631_),
    .Y(net5267));
 BUFx3_ASAP7_75t_R place5268 (.A(_09631_),
    .Y(net5268));
 BUFx3_ASAP7_75t_R place5269 (.A(_01393_),
    .Y(net5269));
 BUFx3_ASAP7_75t_R place5270 (.A(_01393_),
    .Y(net5270));
 BUFx3_ASAP7_75t_R place5271 (.A(_01388_),
    .Y(net5271));
 BUFx3_ASAP7_75t_R place5272 (.A(_01353_),
    .Y(net5272));
 BUFx3_ASAP7_75t_R place5273 (.A(net5274),
    .Y(net5273));
 BUFx3_ASAP7_75t_R place5274 (.A(_01351_),
    .Y(net5274));
 BUFx3_ASAP7_75t_R place5275 (.A(_01349_),
    .Y(net5275));
 BUFx3_ASAP7_75t_R place5276 (.A(_01344_),
    .Y(net5276));
 BUFx3_ASAP7_75t_R place5277 (.A(_01219_),
    .Y(net5277));
 BUFx3_ASAP7_75t_R place5278 (.A(_01218_),
    .Y(net5278));
 BUFx3_ASAP7_75t_R place5279 (.A(_01217_),
    .Y(net5279));
 BUFx3_ASAP7_75t_R place5280 (.A(_01216_),
    .Y(net5280));
 BUFx3_ASAP7_75t_R place5281 (.A(_01214_),
    .Y(net5281));
 BUFx3_ASAP7_75t_R place5282 (.A(_01212_),
    .Y(net5282));
 BUFx3_ASAP7_75t_R place5283 (.A(_01193_),
    .Y(net5283));
 BUFx3_ASAP7_75t_R place5284 (.A(_01191_),
    .Y(net5284));
 BUFx3_ASAP7_75t_R place5285 (.A(_01191_),
    .Y(net5285));
 BUFx6f_ASAP7_75t_R place5286 (.A(_01177_),
    .Y(net5286));
 BUFx3_ASAP7_75t_R place5287 (.A(_01175_),
    .Y(net5287));
 BUFx3_ASAP7_75t_R place5288 (.A(_01174_),
    .Y(net5288));
 BUFx3_ASAP7_75t_R place5289 (.A(_01172_),
    .Y(net5289));
 BUFx3_ASAP7_75t_R place5290 (.A(_01170_),
    .Y(net5290));
 BUFx3_ASAP7_75t_R place5291 (.A(_01156_),
    .Y(net5291));
 BUFx3_ASAP7_75t_R place5292 (.A(_01154_),
    .Y(net5292));
 BUFx3_ASAP7_75t_R place5293 (.A(_01153_),
    .Y(net5293));
 BUFx3_ASAP7_75t_R place5294 (.A(_01135_),
    .Y(net5294));
 BUFx3_ASAP7_75t_R place5295 (.A(_01130_),
    .Y(net5295));
 BUFx6f_ASAP7_75t_R place5296 (.A(_01114_),
    .Y(net5296));
 BUFx3_ASAP7_75t_R place5297 (.A(net5298),
    .Y(net5297));
 BUFx3_ASAP7_75t_R place5298 (.A(_01109_),
    .Y(net5298));
 BUFx3_ASAP7_75t_R place5299 (.A(_01093_),
    .Y(net5299));
 BUFx3_ASAP7_75t_R place5300 (.A(_01091_),
    .Y(net5300));
 BUFx3_ASAP7_75t_R place5301 (.A(_01090_),
    .Y(net5301));
 BUFx3_ASAP7_75t_R place5302 (.A(_01088_),
    .Y(net5302));
 BUFx3_ASAP7_75t_R place5303 (.A(_01086_),
    .Y(net5303));
 BUFx3_ASAP7_75t_R place5304 (.A(_01072_),
    .Y(net5304));
 BUFx3_ASAP7_75t_R place5305 (.A(_01069_),
    .Y(net5305));
 BUFx3_ASAP7_75t_R place5306 (.A(_01069_),
    .Y(net5306));
 BUFx6f_ASAP7_75t_R place5307 (.A(net5308),
    .Y(net5307));
 BUFx3_ASAP7_75t_R place5308 (.A(_01067_),
    .Y(net5308));
 BUFx6f_ASAP7_75t_R place5309 (.A(_01065_),
    .Y(net5309));
 BUFx3_ASAP7_75t_R place5310 (.A(_01051_),
    .Y(net5310));
 BUFx3_ASAP7_75t_R place5311 (.A(_01049_),
    .Y(net5311));
 BUFx3_ASAP7_75t_R place5312 (.A(_01029_),
    .Y(net5312));
 BUFx3_ASAP7_75t_R place5313 (.A(_01028_),
    .Y(net5313));
 BUFx3_ASAP7_75t_R place5314 (.A(_01027_),
    .Y(net5314));
 BUFx3_ASAP7_75t_R place5315 (.A(_01026_),
    .Y(net5315));
 BUFx3_ASAP7_75t_R place5316 (.A(_01007_),
    .Y(net5316));
 BUFx3_ASAP7_75t_R place5317 (.A(net5318),
    .Y(net5317));
 BUFx3_ASAP7_75t_R place5318 (.A(_01002_),
    .Y(net5318));
 BUFx3_ASAP7_75t_R place5319 (.A(_01001_),
    .Y(net5319));
 BUFx3_ASAP7_75t_R place5320 (.A(_00999_),
    .Y(net5320));
 BUFx3_ASAP7_75t_R place5321 (.A(_00978_),
    .Y(net5321));
 BUFx3_ASAP7_75t_R place5322 (.A(_00976_),
    .Y(net5322));
 BUFx3_ASAP7_75t_R place5323 (.A(_00974_),
    .Y(net5323));
 BUFx3_ASAP7_75t_R place5324 (.A(_07463_),
    .Y(net5324));
 BUFx3_ASAP7_75t_R place5325 (.A(_07345_),
    .Y(net5325));
 BUFx3_ASAP7_75t_R place5326 (.A(_07342_),
    .Y(net5326));
 BUFx3_ASAP7_75t_R place5327 (.A(_07342_),
    .Y(net5327));
 BUFx6f_ASAP7_75t_R place5328 (.A(_07298_),
    .Y(net5328));
 BUFx3_ASAP7_75t_R place5329 (.A(_07289_),
    .Y(net5329));
 BUFx3_ASAP7_75t_R place5330 (.A(_07231_),
    .Y(net5330));
 BUFx3_ASAP7_75t_R place5331 (.A(_07200_),
    .Y(net5331));
 BUFx3_ASAP7_75t_R place5332 (.A(net5333),
    .Y(net5332));
 BUFx3_ASAP7_75t_R place5333 (.A(_07186_),
    .Y(net5333));
 BUFx3_ASAP7_75t_R place5334 (.A(_07183_),
    .Y(net5334));
 BUFx6f_ASAP7_75t_R place5335 (.A(_07169_),
    .Y(net5335));
 BUFx3_ASAP7_75t_R place5336 (.A(_01389_),
    .Y(net5336));
 BUFx3_ASAP7_75t_R place5337 (.A(_01389_),
    .Y(net5337));
 BUFx3_ASAP7_75t_R place5338 (.A(_06866_),
    .Y(net5338));
 BUFx3_ASAP7_75t_R place5339 (.A(_06781_),
    .Y(net5339));
 BUFx3_ASAP7_75t_R place5340 (.A(_06707_),
    .Y(net5340));
 BUFx3_ASAP7_75t_R place5341 (.A(_06707_),
    .Y(net5341));
 BUFx3_ASAP7_75t_R place5342 (.A(_06678_),
    .Y(net5342));
 BUFx3_ASAP7_75t_R place5343 (.A(_06632_),
    .Y(net5343));
 BUFx3_ASAP7_75t_R place5344 (.A(_06632_),
    .Y(net5344));
 BUFx3_ASAP7_75t_R place5345 (.A(_06632_),
    .Y(net5345));
 BUFx6f_ASAP7_75t_R place5346 (.A(_06595_),
    .Y(net5346));
 BUFx3_ASAP7_75t_R place5347 (.A(_06583_),
    .Y(net5347));
 BUFx3_ASAP7_75t_R place5348 (.A(net5350),
    .Y(net5348));
 BUFx3_ASAP7_75t_R place5349 (.A(net5350),
    .Y(net5349));
 BUFx6f_ASAP7_75t_R place5350 (.A(_06551_),
    .Y(net5350));
 BUFx6f_ASAP7_75t_R place5351 (.A(_06534_),
    .Y(net5351));
 BUFx3_ASAP7_75t_R place5352 (.A(_06054_),
    .Y(net5352));
 BUFx3_ASAP7_75t_R place5353 (.A(_06054_),
    .Y(net5353));
 BUFx3_ASAP7_75t_R place5354 (.A(_05977_),
    .Y(net5354));
 BUFx6f_ASAP7_75t_R place5355 (.A(_05969_),
    .Y(net5355));
 BUFx3_ASAP7_75t_R place5356 (.A(_05944_),
    .Y(net5356));
 BUFx6f_ASAP7_75t_R place5357 (.A(_05933_),
    .Y(net5357));
 BUFx3_ASAP7_75t_R place5358 (.A(_05932_),
    .Y(net5358));
 BUFx3_ASAP7_75t_R place5359 (.A(net5360),
    .Y(net5359));
 BUFx6f_ASAP7_75t_R place5360 (.A(_05918_),
    .Y(net5360));
 BUFx3_ASAP7_75t_R place5361 (.A(_05885_),
    .Y(net5361));
 BUFx3_ASAP7_75t_R place5362 (.A(_05851_),
    .Y(net5362));
 BUFx3_ASAP7_75t_R place5363 (.A(_05846_),
    .Y(net5363));
 BUFx6f_ASAP7_75t_R place5364 (.A(_05806_),
    .Y(net5364));
 BUFx3_ASAP7_75t_R place5365 (.A(_05305_),
    .Y(net5365));
 BUFx3_ASAP7_75t_R place5366 (.A(_05266_),
    .Y(net5366));
 BUFx6f_ASAP7_75t_R place5367 (.A(_05266_),
    .Y(net5367));
 BUFx3_ASAP7_75t_R place5368 (.A(_05262_),
    .Y(net5368));
 BUFx3_ASAP7_75t_R place5369 (.A(net5371),
    .Y(net5369));
 BUFx6f_ASAP7_75t_R place5370 (.A(net5371),
    .Y(net5370));
 BUFx3_ASAP7_75t_R place5371 (.A(_05248_),
    .Y(net5371));
 BUFx3_ASAP7_75t_R place5372 (.A(_05242_),
    .Y(net5372));
 BUFx3_ASAP7_75t_R place5373 (.A(net5374),
    .Y(net5373));
 BUFx3_ASAP7_75t_R place5374 (.A(_01321_),
    .Y(net5374));
 BUFx3_ASAP7_75t_R place5375 (.A(_05161_),
    .Y(net5375));
 BUFx3_ASAP7_75t_R place5376 (.A(_05161_),
    .Y(net5376));
 BUFx3_ASAP7_75t_R place5377 (.A(_05161_),
    .Y(net5377));
 BUFx3_ASAP7_75t_R place5378 (.A(net5379),
    .Y(net5378));
 BUFx3_ASAP7_75t_R place5379 (.A(_04500_),
    .Y(net5379));
 BUFx3_ASAP7_75t_R place5380 (.A(_04472_),
    .Y(net5380));
 BUFx3_ASAP7_75t_R place5381 (.A(_04432_),
    .Y(net5381));
 BUFx3_ASAP7_75t_R place5382 (.A(_04421_),
    .Y(net5382));
 BUFx3_ASAP7_75t_R place5383 (.A(_01303_),
    .Y(net5383));
 BUFx6f_ASAP7_75t_R place5384 (.A(net5385),
    .Y(net5384));
 BUFx3_ASAP7_75t_R place5385 (.A(_03796_),
    .Y(net5385));
 BUFx3_ASAP7_75t_R place5386 (.A(_03720_),
    .Y(net5386));
 BUFx6f_ASAP7_75t_R place5387 (.A(_03720_),
    .Y(net5387));
 BUFx6f_ASAP7_75t_R place5388 (.A(_03713_),
    .Y(net5388));
 BUFx3_ASAP7_75t_R place5389 (.A(_01280_),
    .Y(net5389));
 BUFx3_ASAP7_75t_R place5390 (.A(_01280_),
    .Y(net5390));
 BUFx3_ASAP7_75t_R place5391 (.A(_03163_),
    .Y(net5391));
 BUFx3_ASAP7_75t_R place5392 (.A(_03163_),
    .Y(net5392));
 BUFx3_ASAP7_75t_R place5393 (.A(_03163_),
    .Y(net5393));
 BUFx3_ASAP7_75t_R place5394 (.A(_03163_),
    .Y(net5394));
 BUFx3_ASAP7_75t_R place5395 (.A(_01253_),
    .Y(net5395));
 BUFx6f_ASAP7_75t_R place5396 (.A(_03035_),
    .Y(net5396));
 BUFx3_ASAP7_75t_R place5397 (.A(net5398),
    .Y(net5397));
 BUFx6f_ASAP7_75t_R place5398 (.A(_03035_),
    .Y(net5398));
 BUFx3_ASAP7_75t_R place5399 (.A(_03031_),
    .Y(net5399));
 BUFx3_ASAP7_75t_R place5400 (.A(_03031_),
    .Y(net5400));
 BUFx3_ASAP7_75t_R place5401 (.A(_03011_),
    .Y(net5401));
 BUFx3_ASAP7_75t_R place5402 (.A(net5403),
    .Y(net5402));
 BUFx6f_ASAP7_75t_R place5403 (.A(_03011_),
    .Y(net5403));
 BUFx6f_ASAP7_75t_R place5404 (.A(_02413_),
    .Y(net5404));
 BUFx3_ASAP7_75t_R place5405 (.A(_02413_),
    .Y(net5405));
 BUFx6f_ASAP7_75t_R place5406 (.A(_02376_),
    .Y(net5406));
 BUFx3_ASAP7_75t_R place5407 (.A(_02376_),
    .Y(net5407));
 BUFx6f_ASAP7_75t_R place5408 (.A(net5409),
    .Y(net5408));
 BUFx6f_ASAP7_75t_R place5409 (.A(_02376_),
    .Y(net5409));
 BUFx3_ASAP7_75t_R place5410 (.A(_02376_),
    .Y(net5410));
 BUFx3_ASAP7_75t_R place5411 (.A(_02376_),
    .Y(net5411));
 BUFx6f_ASAP7_75t_R place5412 (.A(_02342_),
    .Y(net5412));
 BUFx6f_ASAP7_75t_R place5413 (.A(_02336_),
    .Y(net5413));
 BUFx3_ASAP7_75t_R place5414 (.A(_02336_),
    .Y(net5414));
 BUFx3_ASAP7_75t_R place5415 (.A(_01237_),
    .Y(net5415));
 BUFx3_ASAP7_75t_R place5416 (.A(_01237_),
    .Y(net5416));
 BUFx3_ASAP7_75t_R place5417 (.A(_02219_),
    .Y(net5417));
 BUFx3_ASAP7_75t_R place5418 (.A(_01785_),
    .Y(net5418));
 BUFx3_ASAP7_75t_R place5419 (.A(_01785_),
    .Y(net5419));
 BUFx3_ASAP7_75t_R place5420 (.A(_01758_),
    .Y(net5420));
 BUFx3_ASAP7_75t_R place5421 (.A(_01753_),
    .Y(net5421));
 BUFx6f_ASAP7_75t_R place5422 (.A(_01753_),
    .Y(net5422));
 BUFx3_ASAP7_75t_R place5423 (.A(_01702_),
    .Y(net5423));
 BUFx6f_ASAP7_75t_R place5424 (.A(_01702_),
    .Y(net5424));
 BUFx3_ASAP7_75t_R place5425 (.A(_01675_),
    .Y(net5425));
 BUFx6f_ASAP7_75t_R place5426 (.A(_01675_),
    .Y(net5426));
 BUFx3_ASAP7_75t_R place5427 (.A(_01654_),
    .Y(net5427));
 BUFx6f_ASAP7_75t_R place5428 (.A(_01654_),
    .Y(net5428));
 BUFx6f_ASAP7_75t_R place5429 (.A(_01654_),
    .Y(net5429));
 BUFx3_ASAP7_75t_R place5430 (.A(net5433),
    .Y(net5430));
 BUFx6f_ASAP7_75t_R place5431 (.A(net5433),
    .Y(net5431));
 BUFx3_ASAP7_75t_R place5432 (.A(net5433),
    .Y(net5432));
 BUFx6f_ASAP7_75t_R place5433 (.A(_01639_),
    .Y(net5433));
 BUFx3_ASAP7_75t_R place5434 (.A(_01634_),
    .Y(net5434));
 BUFx6f_ASAP7_75t_R place5435 (.A(_01634_),
    .Y(net5435));
 BUFx3_ASAP7_75t_R place5436 (.A(net5437),
    .Y(net5436));
 BUFx6f_ASAP7_75t_R place5437 (.A(_01634_),
    .Y(net5437));
 BUFx3_ASAP7_75t_R place5438 (.A(_15213_),
    .Y(net5438));
 BUFx3_ASAP7_75t_R place5439 (.A(_15171_),
    .Y(net5439));
 BUFx6f_ASAP7_75t_R place5440 (.A(_15060_),
    .Y(net5440));
 BUFx3_ASAP7_75t_R place5441 (.A(_15060_),
    .Y(net5441));
 BUFx3_ASAP7_75t_R place5442 (.A(net5443),
    .Y(net5442));
 BUFx6f_ASAP7_75t_R place5443 (.A(_15030_),
    .Y(net5443));
 BUFx6f_ASAP7_75t_R place5444 (.A(_14974_),
    .Y(net5444));
 BUFx6f_ASAP7_75t_R place5445 (.A(_14974_),
    .Y(net5445));
 BUFx3_ASAP7_75t_R place5446 (.A(_14974_),
    .Y(net5446));
 BUFx6f_ASAP7_75t_R place5447 (.A(_14974_),
    .Y(net5447));
 BUFx6f_ASAP7_75t_R place5448 (.A(_14967_),
    .Y(net5448));
 BUFx6f_ASAP7_75t_R place5449 (.A(_14967_),
    .Y(net5449));
 BUFx6f_ASAP7_75t_R place5450 (.A(net5451),
    .Y(net5450));
 BUFx6f_ASAP7_75t_R place5451 (.A(_14967_),
    .Y(net5451));
 BUFx3_ASAP7_75t_R place5452 (.A(_01194_),
    .Y(net5452));
 BUFx3_ASAP7_75t_R place5453 (.A(_14541_),
    .Y(net5453));
 BUFx3_ASAP7_75t_R place5454 (.A(_14541_),
    .Y(net5454));
 BUFx3_ASAP7_75t_R place5455 (.A(_14517_),
    .Y(net5455));
 BUFx3_ASAP7_75t_R place5456 (.A(_14515_),
    .Y(net5456));
 BUFx3_ASAP7_75t_R place5457 (.A(_14388_),
    .Y(net5457));
 BUFx3_ASAP7_75t_R place5458 (.A(_14388_),
    .Y(net5458));
 BUFx3_ASAP7_75t_R place5459 (.A(_14348_),
    .Y(net5459));
 BUFx3_ASAP7_75t_R place5460 (.A(_14339_),
    .Y(net5460));
 BUFx6f_ASAP7_75t_R place5461 (.A(_14339_),
    .Y(net5461));
 BUFx3_ASAP7_75t_R place5462 (.A(_14310_),
    .Y(net5462));
 BUFx3_ASAP7_75t_R place5463 (.A(net5465),
    .Y(net5463));
 BUFx6f_ASAP7_75t_R place5464 (.A(net5465),
    .Y(net5464));
 BUFx6f_ASAP7_75t_R place5465 (.A(_13678_),
    .Y(net5465));
 BUFx6f_ASAP7_75t_R place5466 (.A(net5475),
    .Y(net5466));
 BUFx3_ASAP7_75t_R place5467 (.A(net5475),
    .Y(net5467));
 BUFx6f_ASAP7_75t_R place5468 (.A(net5475),
    .Y(net5468));
 BUFx3_ASAP7_75t_R place5469 (.A(net5475),
    .Y(net5469));
 BUFx3_ASAP7_75t_R place5470 (.A(net5475),
    .Y(net5470));
 BUFx3_ASAP7_75t_R place5471 (.A(net5475),
    .Y(net5471));
 BUFx3_ASAP7_75t_R place5472 (.A(net5475),
    .Y(net5472));
 BUFx3_ASAP7_75t_R place5473 (.A(net5474),
    .Y(net5473));
 BUFx6f_ASAP7_75t_R place5474 (.A(net5475),
    .Y(net5474));
 BUFx6f_ASAP7_75t_R place5475 (.A(_13639_),
    .Y(net5475));
 BUFx6f_ASAP7_75t_R place5476 (.A(_13613_),
    .Y(net5476));
 BUFx3_ASAP7_75t_R place5477 (.A(_13613_),
    .Y(net5477));
 BUFx3_ASAP7_75t_R place5478 (.A(_13613_),
    .Y(net5478));
 BUFx6f_ASAP7_75t_R place5479 (.A(_13613_),
    .Y(net5479));
 BUFx6f_ASAP7_75t_R place5480 (.A(net5482),
    .Y(net5480));
 BUFx3_ASAP7_75t_R place5481 (.A(net5482),
    .Y(net5481));
 BUFx6f_ASAP7_75t_R place5482 (.A(_13580_),
    .Y(net5482));
 BUFx3_ASAP7_75t_R place5483 (.A(net5484),
    .Y(net5483));
 BUFx3_ASAP7_75t_R place5484 (.A(_13576_),
    .Y(net5484));
 BUFx3_ASAP7_75t_R place5485 (.A(net5486),
    .Y(net5485));
 BUFx6f_ASAP7_75t_R place5486 (.A(_13571_),
    .Y(net5486));
 BUFx3_ASAP7_75t_R place5487 (.A(_13571_),
    .Y(net5487));
 BUFx3_ASAP7_75t_R place5488 (.A(_13160_),
    .Y(net5488));
 BUFx3_ASAP7_75t_R place5489 (.A(_13132_),
    .Y(net5489));
 BUFx3_ASAP7_75t_R place5490 (.A(_13099_),
    .Y(net5490));
 BUFx3_ASAP7_75t_R place5491 (.A(_13099_),
    .Y(net5491));
 BUFx3_ASAP7_75t_R place5492 (.A(_13099_),
    .Y(net5492));
 BUFx3_ASAP7_75t_R place5493 (.A(_13073_),
    .Y(net5493));
 BUFx3_ASAP7_75t_R place5494 (.A(_13073_),
    .Y(net5494));
 BUFx3_ASAP7_75t_R place5495 (.A(_13073_),
    .Y(net5495));
 BUFx3_ASAP7_75t_R place5496 (.A(_01125_),
    .Y(net5496));
 BUFx3_ASAP7_75t_R place5497 (.A(_13062_),
    .Y(net5497));
 BUFx3_ASAP7_75t_R place5498 (.A(_13062_),
    .Y(net5498));
 BUFx3_ASAP7_75t_R place5499 (.A(_13062_),
    .Y(net5499));
 BUFx3_ASAP7_75t_R place5500 (.A(_13062_),
    .Y(net5500));
 BUFx3_ASAP7_75t_R place5501 (.A(_13052_),
    .Y(net5501));
 BUFx3_ASAP7_75t_R place5502 (.A(_13043_),
    .Y(net5502));
 BUFx6f_ASAP7_75t_R place5503 (.A(_12990_),
    .Y(net5503));
 BUFx3_ASAP7_75t_R place5504 (.A(_12944_),
    .Y(net5504));
 BUFx3_ASAP7_75t_R place5505 (.A(_12943_),
    .Y(net5505));
 BUFx3_ASAP7_75t_R place5506 (.A(_12507_),
    .Y(net5506));
 BUFx3_ASAP7_75t_R place5507 (.A(net5508),
    .Y(net5507));
 BUFx3_ASAP7_75t_R place5508 (.A(_01104_),
    .Y(net5508));
 BUFx3_ASAP7_75t_R place5509 (.A(_12353_),
    .Y(net5509));
 BUFx3_ASAP7_75t_R place5510 (.A(_12336_),
    .Y(net5510));
 BUFx3_ASAP7_75t_R place5511 (.A(_12311_),
    .Y(net5511));
 BUFx6f_ASAP7_75t_R place5512 (.A(_12263_),
    .Y(net5512));
 BUFx3_ASAP7_75t_R place5513 (.A(net5514),
    .Y(net5513));
 BUFx3_ASAP7_75t_R place5514 (.A(_12263_),
    .Y(net5514));
 BUFx3_ASAP7_75t_R place5515 (.A(_12250_),
    .Y(net5515));
 BUFx3_ASAP7_75t_R place5516 (.A(_12250_),
    .Y(net5516));
 BUFx6f_ASAP7_75t_R place5517 (.A(_12224_),
    .Y(net5517));
 BUFx6f_ASAP7_75t_R place5518 (.A(_12174_),
    .Y(net5518));
 BUFx3_ASAP7_75t_R place5519 (.A(_11700_),
    .Y(net5519));
 BUFx3_ASAP7_75t_R place5520 (.A(_11642_),
    .Y(net5520));
 BUFx3_ASAP7_75t_R place5521 (.A(_11636_),
    .Y(net5521));
 BUFx6f_ASAP7_75t_R place5522 (.A(_11586_),
    .Y(net5522));
 BUFx3_ASAP7_75t_R place5523 (.A(_11452_),
    .Y(net5523));
 BUFx6f_ASAP7_75t_R place5524 (.A(_11452_),
    .Y(net5524));
 BUFx6f_ASAP7_75t_R place5525 (.A(_10999_),
    .Y(net5525));
 BUFx3_ASAP7_75t_R place5526 (.A(_10952_),
    .Y(net5526));
 BUFx3_ASAP7_75t_R place5527 (.A(_10944_),
    .Y(net5527));
 BUFx3_ASAP7_75t_R place5528 (.A(_10891_),
    .Y(net5528));
 BUFx3_ASAP7_75t_R place5529 (.A(_10885_),
    .Y(net5529));
 BUFx6f_ASAP7_75t_R place5530 (.A(_10870_),
    .Y(net5530));
 BUFx3_ASAP7_75t_R place5531 (.A(_10836_),
    .Y(net5531));
 BUFx3_ASAP7_75t_R place5532 (.A(_10836_),
    .Y(net5532));
 BUFx3_ASAP7_75t_R place5533 (.A(_10813_),
    .Y(net5533));
 BUFx3_ASAP7_75t_R place5534 (.A(_10236_),
    .Y(net5534));
 BUFx3_ASAP7_75t_R place5535 (.A(_10197_),
    .Y(net5535));
 BUFx3_ASAP7_75t_R place5536 (.A(_10187_),
    .Y(net5536));
 BUFx3_ASAP7_75t_R place5537 (.A(_10165_),
    .Y(net5537));
 BUFx3_ASAP7_75t_R place5538 (.A(_10138_),
    .Y(net5538));
 BUFx3_ASAP7_75t_R place5539 (.A(_10126_),
    .Y(net5539));
 BUFx6f_ASAP7_75t_R place5540 (.A(_10126_),
    .Y(net5540));
 BUFx6f_ASAP7_75t_R place5541 (.A(_10126_),
    .Y(net5541));
 BUFx3_ASAP7_75t_R place5542 (.A(_09653_),
    .Y(net5542));
 BUFx3_ASAP7_75t_R place5543 (.A(_09653_),
    .Y(net5543));
 BUFx3_ASAP7_75t_R place5544 (.A(_09621_),
    .Y(net5544));
 BUFx3_ASAP7_75t_R place5545 (.A(_09621_),
    .Y(net5545));
 BUFx3_ASAP7_75t_R place5546 (.A(_09608_),
    .Y(net5546));
 BUFx6f_ASAP7_75t_R place5547 (.A(_09607_),
    .Y(net5547));
 BUFx3_ASAP7_75t_R place5548 (.A(_09577_),
    .Y(net5548));
 BUFx3_ASAP7_75t_R place5549 (.A(_09143_),
    .Y(net5549));
 BUFx6f_ASAP7_75t_R place5550 (.A(_09121_),
    .Y(net5550));
 BUFx3_ASAP7_75t_R place5551 (.A(_09114_),
    .Y(net5551));
 BUFx3_ASAP7_75t_R place5552 (.A(net5553),
    .Y(net5552));
 BUFx6f_ASAP7_75t_R place5553 (.A(_09114_),
    .Y(net5553));
 BUFx6f_ASAP7_75t_R place5554 (.A(_09073_),
    .Y(net5554));
 BUFx3_ASAP7_75t_R place5555 (.A(_09060_),
    .Y(net5555));
 BUFx3_ASAP7_75t_R place5556 (.A(_09054_),
    .Y(net5556));
 BUFx3_ASAP7_75t_R place5557 (.A(_09034_),
    .Y(net5557));
 BUFx6f_ASAP7_75t_R place5558 (.A(_09027_),
    .Y(net5558));
 BUFx3_ASAP7_75t_R place5559 (.A(_08414_),
    .Y(net5559));
 BUFx3_ASAP7_75t_R place5560 (.A(_08320_),
    .Y(net5560));
 BUFx3_ASAP7_75t_R place5561 (.A(_08137_),
    .Y(net5561));
 BUFx3_ASAP7_75t_R place5562 (.A(_01042_),
    .Y(net5562));
 BUFx3_ASAP7_75t_R place5563 (.A(_01020_),
    .Y(net5563));
 BUFx3_ASAP7_75t_R place5564 (.A(_01046_),
    .Y(net5564));
 BUFx3_ASAP7_75t_R place5565 (.A(_01045_),
    .Y(net5565));
 BUFx3_ASAP7_75t_R place5566 (.A(_01043_),
    .Y(net5566));
 BUFx3_ASAP7_75t_R place5567 (.A(_01041_),
    .Y(net5567));
 BUFx3_ASAP7_75t_R place5568 (.A(_01024_),
    .Y(net5568));
 BUFx3_ASAP7_75t_R place5569 (.A(_01023_),
    .Y(net5569));
 BUFx3_ASAP7_75t_R place5570 (.A(_01005_),
    .Y(net5570));
 BUFx3_ASAP7_75t_R place5571 (.A(_01004_),
    .Y(net5571));
 BUFx3_ASAP7_75t_R place5572 (.A(_00984_),
    .Y(net5572));
 BUFx3_ASAP7_75t_R place5573 (.A(_07352_),
    .Y(net5573));
 BUFx6f_ASAP7_75t_R place5574 (.A(_07243_),
    .Y(net5574));
 BUFx3_ASAP7_75t_R place5575 (.A(_01384_),
    .Y(net5575));
 BUFx6f_ASAP7_75t_R place5576 (.A(_07158_),
    .Y(net5576));
 BUFx3_ASAP7_75t_R place5577 (.A(net5580),
    .Y(net5577));
 BUFx3_ASAP7_75t_R place5578 (.A(net5580),
    .Y(net5578));
 BUFx3_ASAP7_75t_R place5579 (.A(net5580),
    .Y(net5579));
 BUFx6f_ASAP7_75t_R place5580 (.A(_07158_),
    .Y(net5580));
 BUFx6f_ASAP7_75t_R place5581 (.A(_07153_),
    .Y(net5581));
 BUFx6f_ASAP7_75t_R place5582 (.A(_07153_),
    .Y(net5582));
 BUFx3_ASAP7_75t_R place5583 (.A(net5585),
    .Y(net5583));
 BUFx3_ASAP7_75t_R place5584 (.A(net5585),
    .Y(net5584));
 BUFx3_ASAP7_75t_R place5585 (.A(_07136_),
    .Y(net5585));
 BUFx3_ASAP7_75t_R place5586 (.A(_07123_),
    .Y(net5586));
 BUFx3_ASAP7_75t_R place5587 (.A(_07123_),
    .Y(net5587));
 BUFx3_ASAP7_75t_R place5588 (.A(_06622_),
    .Y(net5588));
 BUFx3_ASAP7_75t_R place5589 (.A(_06622_),
    .Y(net5589));
 BUFx3_ASAP7_75t_R place5590 (.A(_06582_),
    .Y(net5590));
 BUFx6f_ASAP7_75t_R place5591 (.A(_06550_),
    .Y(net5591));
 BUFx3_ASAP7_75t_R place5592 (.A(_06538_),
    .Y(net5592));
 BUFx3_ASAP7_75t_R place5593 (.A(_06538_),
    .Y(net5593));
 BUFx6f_ASAP7_75t_R place5594 (.A(_06538_),
    .Y(net5594));
 BUFx6f_ASAP7_75t_R place5595 (.A(net5597),
    .Y(net5595));
 BUFx3_ASAP7_75t_R place5596 (.A(net5597),
    .Y(net5596));
 BUFx6f_ASAP7_75t_R place5597 (.A(_06496_),
    .Y(net5597));
 BUFx3_ASAP7_75t_R place5598 (.A(net5599),
    .Y(net5598));
 BUFx6f_ASAP7_75t_R place5599 (.A(_06496_),
    .Y(net5599));
 BUFx6f_ASAP7_75t_R place5600 (.A(_06489_),
    .Y(net5600));
 BUFx3_ASAP7_75t_R place5601 (.A(_06464_),
    .Y(net5601));
 BUFx3_ASAP7_75t_R place5602 (.A(_06457_),
    .Y(net5602));
 BUFx3_ASAP7_75t_R place5603 (.A(_06457_),
    .Y(net5603));
 BUFx6f_ASAP7_75t_R place5604 (.A(_05880_),
    .Y(net5604));
 BUFx3_ASAP7_75t_R place5605 (.A(net5606),
    .Y(net5605));
 BUFx6f_ASAP7_75t_R place5606 (.A(_05870_),
    .Y(net5606));
 BUFx3_ASAP7_75t_R place5607 (.A(net5608),
    .Y(net5607));
 BUFx3_ASAP7_75t_R place5608 (.A(_05845_),
    .Y(net5608));
 BUFx3_ASAP7_75t_R place5609 (.A(_05839_),
    .Y(net5609));
 BUFx6f_ASAP7_75t_R place5610 (.A(_05839_),
    .Y(net5610));
 BUFx6f_ASAP7_75t_R place5611 (.A(_05839_),
    .Y(net5611));
 BUFx3_ASAP7_75t_R place5612 (.A(net5614),
    .Y(net5612));
 BUFx3_ASAP7_75t_R place5613 (.A(net5614),
    .Y(net5613));
 BUFx6f_ASAP7_75t_R place5614 (.A(_05839_),
    .Y(net5614));
 BUFx3_ASAP7_75t_R place5615 (.A(net5616),
    .Y(net5615));
 BUFx6f_ASAP7_75t_R place5616 (.A(_05805_),
    .Y(net5616));
 BUFx3_ASAP7_75t_R place5617 (.A(net5619),
    .Y(net5617));
 BUFx3_ASAP7_75t_R place5618 (.A(net5619),
    .Y(net5618));
 BUFx3_ASAP7_75t_R place5619 (.A(_05800_),
    .Y(net5619));
 BUFx6f_ASAP7_75t_R place5620 (.A(net5623),
    .Y(net5620));
 BUFx3_ASAP7_75t_R place5621 (.A(net5623),
    .Y(net5621));
 BUFx3_ASAP7_75t_R place5622 (.A(net5623),
    .Y(net5622));
 BUFx6f_ASAP7_75t_R place5623 (.A(_05793_),
    .Y(net5623));
 BUFx3_ASAP7_75t_R place5624 (.A(_05777_),
    .Y(net5624));
 BUFx3_ASAP7_75t_R place5625 (.A(_05777_),
    .Y(net5625));
 BUFx3_ASAP7_75t_R place5626 (.A(_05777_),
    .Y(net5626));
 BUFx3_ASAP7_75t_R place5627 (.A(net5628),
    .Y(net5627));
 BUFx3_ASAP7_75t_R place5628 (.A(net5629),
    .Y(net5628));
 BUFx3_ASAP7_75t_R place5629 (.A(_05766_),
    .Y(net5629));
 BUFx3_ASAP7_75t_R place5630 (.A(_05766_),
    .Y(net5630));
 BUFx3_ASAP7_75t_R place5631 (.A(_05237_),
    .Y(net5631));
 BUFx3_ASAP7_75t_R place5632 (.A(net5635),
    .Y(net5632));
 BUFx3_ASAP7_75t_R place5633 (.A(net5635),
    .Y(net5633));
 BUFx3_ASAP7_75t_R place5634 (.A(net5635),
    .Y(net5634));
 BUFx6f_ASAP7_75t_R place5635 (.A(_05186_),
    .Y(net5635));
 BUFx6f_ASAP7_75t_R place5636 (.A(_05127_),
    .Y(net5636));
 BUFx6f_ASAP7_75t_R place5637 (.A(_05127_),
    .Y(net5637));
 BUFx6f_ASAP7_75t_R place5638 (.A(_05119_),
    .Y(net5638));
 BUFx3_ASAP7_75t_R place5639 (.A(_05119_),
    .Y(net5639));
 BUFx3_ASAP7_75t_R place5640 (.A(net5642),
    .Y(net5640));
 BUFx3_ASAP7_75t_R place5641 (.A(net5642),
    .Y(net5641));
 BUFx3_ASAP7_75t_R place5642 (.A(_05087_),
    .Y(net5642));
 BUFx3_ASAP7_75t_R place5643 (.A(_04849_),
    .Y(net5643));
 BUFx6f_ASAP7_75t_R place5644 (.A(_04536_),
    .Y(net5644));
 BUFx3_ASAP7_75t_R place5645 (.A(_04498_),
    .Y(net5645));
 BUFx3_ASAP7_75t_R place5646 (.A(_04492_),
    .Y(net5646));
 BUFx3_ASAP7_75t_R place5647 (.A(net5649),
    .Y(net5647));
 BUFx3_ASAP7_75t_R place5648 (.A(net5649),
    .Y(net5648));
 BUFx6f_ASAP7_75t_R place5649 (.A(_04492_),
    .Y(net5649));
 BUFx6f_ASAP7_75t_R place5650 (.A(net5655),
    .Y(net5650));
 BUFx3_ASAP7_75t_R place5651 (.A(net5655),
    .Y(net5651));
 BUFx3_ASAP7_75t_R place5652 (.A(net5655),
    .Y(net5652));
 BUFx3_ASAP7_75t_R place5653 (.A(net5655),
    .Y(net5653));
 BUFx6f_ASAP7_75t_R place5654 (.A(net5655),
    .Y(net5654));
 BUFx6f_ASAP7_75t_R place5655 (.A(_04492_),
    .Y(net5655));
 BUFx3_ASAP7_75t_R place5656 (.A(_04475_),
    .Y(net5656));
 BUFx3_ASAP7_75t_R place5657 (.A(_04469_),
    .Y(net5657));
 BUFx6f_ASAP7_75t_R place5658 (.A(_04469_),
    .Y(net5658));
 BUFx6f_ASAP7_75t_R place5659 (.A(_04456_),
    .Y(net5659));
 BUFx3_ASAP7_75t_R place5660 (.A(_04456_),
    .Y(net5660));
 BUFx6f_ASAP7_75t_R place5661 (.A(_04456_),
    .Y(net5661));
 BUFx3_ASAP7_75t_R place5662 (.A(_04433_),
    .Y(net5662));
 BUFx3_ASAP7_75t_R place5663 (.A(_04431_),
    .Y(net5663));
 BUFx3_ASAP7_75t_R place5664 (.A(_04427_),
    .Y(net5664));
 BUFx3_ASAP7_75t_R place5665 (.A(_01306_),
    .Y(net5665));
 BUFx3_ASAP7_75t_R place5666 (.A(_01306_),
    .Y(net5666));
 BUFx6f_ASAP7_75t_R place5667 (.A(_03880_),
    .Y(net5667));
 BUFx3_ASAP7_75t_R place5668 (.A(_03880_),
    .Y(net5668));
 BUFx3_ASAP7_75t_R place5669 (.A(_03789_),
    .Y(net5669));
 BUFx6f_ASAP7_75t_R place5670 (.A(net5672),
    .Y(net5670));
 BUFx3_ASAP7_75t_R place5671 (.A(net5672),
    .Y(net5671));
 BUFx6f_ASAP7_75t_R place5672 (.A(_03779_),
    .Y(net5672));
 BUFx3_ASAP7_75t_R place5673 (.A(_03765_),
    .Y(net5673));
 BUFx3_ASAP7_75t_R place5674 (.A(_03735_),
    .Y(net5674));
 BUFx3_ASAP7_75t_R place5675 (.A(_01275_),
    .Y(net5675));
 BUFx3_ASAP7_75t_R place5676 (.A(_03706_),
    .Y(net5676));
 BUFx3_ASAP7_75t_R place5677 (.A(net5678),
    .Y(net5677));
 BUFx3_ASAP7_75t_R place5678 (.A(_01283_),
    .Y(net5678));
 BUFx6f_ASAP7_75t_R place5679 (.A(_03208_),
    .Y(net5679));
 BUFx3_ASAP7_75t_R place5680 (.A(_03166_),
    .Y(net5680));
 BUFx6f_ASAP7_75t_R place5681 (.A(_03095_),
    .Y(net5681));
 BUFx3_ASAP7_75t_R place5682 (.A(_03073_),
    .Y(net5682));
 BUFx3_ASAP7_75t_R place5683 (.A(_03066_),
    .Y(net5683));
 BUFx3_ASAP7_75t_R place5684 (.A(_03066_),
    .Y(net5684));
 BUFx6f_ASAP7_75t_R place5685 (.A(_03066_),
    .Y(net5685));
 BUFx6f_ASAP7_75t_R place5686 (.A(_03066_),
    .Y(net5686));
 BUFx6f_ASAP7_75t_R place5687 (.A(_03066_),
    .Y(net5687));
 BUFx3_ASAP7_75t_R place5688 (.A(_03038_),
    .Y(net5688));
 BUFx3_ASAP7_75t_R place5689 (.A(_03033_),
    .Y(net5689));
 BUFx3_ASAP7_75t_R place5690 (.A(net5691),
    .Y(net5690));
 BUFx3_ASAP7_75t_R place5691 (.A(_03032_),
    .Y(net5691));
 BUFx3_ASAP7_75t_R place5692 (.A(_03024_),
    .Y(net5692));
 BUFx3_ASAP7_75t_R place5693 (.A(_01260_),
    .Y(net5693));
 BUFx3_ASAP7_75t_R place5694 (.A(net5695),
    .Y(net5694));
 BUFx6f_ASAP7_75t_R place5695 (.A(_01260_),
    .Y(net5695));
 BUFx3_ASAP7_75t_R place5696 (.A(_02463_),
    .Y(net5696));
 BUFx6f_ASAP7_75t_R place5697 (.A(_02463_),
    .Y(net5697));
 BUFx3_ASAP7_75t_R place5698 (.A(_02463_),
    .Y(net5698));
 BUFx3_ASAP7_75t_R place5699 (.A(_02463_),
    .Y(net5699));
 BUFx6f_ASAP7_75t_R place5700 (.A(_02412_),
    .Y(net5700));
 BUFx3_ASAP7_75t_R place5701 (.A(_02412_),
    .Y(net5701));
 BUFx6f_ASAP7_75t_R place5702 (.A(net5706),
    .Y(net5702));
 BUFx6f_ASAP7_75t_R place5703 (.A(net5706),
    .Y(net5703));
 BUFx3_ASAP7_75t_R place5704 (.A(net5706),
    .Y(net5704));
 BUFx3_ASAP7_75t_R place5705 (.A(net5706),
    .Y(net5705));
 BUFx6f_ASAP7_75t_R place5706 (.A(_02370_),
    .Y(net5706));
 BUFx3_ASAP7_75t_R place5707 (.A(net5708),
    .Y(net5707));
 BUFx6f_ASAP7_75t_R place5708 (.A(_02357_),
    .Y(net5708));
 BUFx6f_ASAP7_75t_R place5709 (.A(_02357_),
    .Y(net5709));
 BUFx3_ASAP7_75t_R place5710 (.A(_02339_),
    .Y(net5710));
 BUFx3_ASAP7_75t_R place5711 (.A(_01230_),
    .Y(net5711));
 BUFx3_ASAP7_75t_R place5712 (.A(_02329_),
    .Y(net5712));
 BUFx3_ASAP7_75t_R place5713 (.A(_02297_),
    .Y(net5713));
 BUFx3_ASAP7_75t_R place5714 (.A(_02297_),
    .Y(net5714));
 BUFx6f_ASAP7_75t_R place5715 (.A(_01733_),
    .Y(net5715));
 BUFx3_ASAP7_75t_R place5716 (.A(net5717),
    .Y(net5716));
 BUFx3_ASAP7_75t_R place5717 (.A(net5718),
    .Y(net5717));
 BUFx6f_ASAP7_75t_R place5718 (.A(_01684_),
    .Y(net5718));
 BUFx6f_ASAP7_75t_R place5719 (.A(_01684_),
    .Y(net5719));
 BUFx3_ASAP7_75t_R place5720 (.A(net5721),
    .Y(net5720));
 BUFx3_ASAP7_75t_R place5721 (.A(_01684_),
    .Y(net5721));
 BUFx3_ASAP7_75t_R place5722 (.A(net5723),
    .Y(net5722));
 BUFx6f_ASAP7_75t_R place5723 (.A(_01684_),
    .Y(net5723));
 BUFx3_ASAP7_75t_R place5724 (.A(_01674_),
    .Y(net5724));
 BUFx6f_ASAP7_75t_R place5725 (.A(net5727),
    .Y(net5725));
 BUFx6f_ASAP7_75t_R place5726 (.A(net5727),
    .Y(net5726));
 BUFx6f_ASAP7_75t_R place5727 (.A(_01670_),
    .Y(net5727));
 BUFx6f_ASAP7_75t_R place5728 (.A(_01670_),
    .Y(net5728));
 BUFx3_ASAP7_75t_R place5729 (.A(_01670_),
    .Y(net5729));
 BUFx3_ASAP7_75t_R place5730 (.A(net5733),
    .Y(net5730));
 BUFx3_ASAP7_75t_R place5731 (.A(net5733),
    .Y(net5731));
 BUFx6f_ASAP7_75t_R place5732 (.A(net5733),
    .Y(net5732));
 BUFx6f_ASAP7_75t_R place5733 (.A(_01670_),
    .Y(net5733));
 BUFx6f_ASAP7_75t_R place5734 (.A(_01670_),
    .Y(net5734));
 BUFx3_ASAP7_75t_R place5735 (.A(net5736),
    .Y(net5735));
 BUFx6f_ASAP7_75t_R place5736 (.A(net5740),
    .Y(net5736));
 BUFx6f_ASAP7_75t_R place5737 (.A(net5740),
    .Y(net5737));
 BUFx3_ASAP7_75t_R place5738 (.A(net5740),
    .Y(net5738));
 BUFx6f_ASAP7_75t_R place5739 (.A(net5740),
    .Y(net5739));
 BUFx6f_ASAP7_75t_R place5740 (.A(_01653_),
    .Y(net5740));
 BUFx3_ASAP7_75t_R place5741 (.A(_01637_),
    .Y(net5741));
 BUFx3_ASAP7_75t_R place5742 (.A(_01636_),
    .Y(net5742));
 BUFx3_ASAP7_75t_R place5743 (.A(_01624_),
    .Y(net5743));
 BUFx6f_ASAP7_75t_R place5744 (.A(_01215_),
    .Y(net5744));
 BUFx3_ASAP7_75t_R place5745 (.A(_01599_),
    .Y(net5745));
 BUFx3_ASAP7_75t_R place5746 (.A(net5747),
    .Y(net5746));
 BUFx3_ASAP7_75t_R place5747 (.A(_01599_),
    .Y(net5747));
 BUFx3_ASAP7_75t_R place5748 (.A(_15102_),
    .Y(net5748));
 BUFx6f_ASAP7_75t_R place5749 (.A(_15102_),
    .Y(net5749));
 BUFx3_ASAP7_75t_R place5750 (.A(_15080_),
    .Y(net5750));
 BUFx6f_ASAP7_75t_R place5751 (.A(_15051_),
    .Y(net5751));
 BUFx3_ASAP7_75t_R place5752 (.A(_15051_),
    .Y(net5752));
 BUFx6f_ASAP7_75t_R place5753 (.A(net5763),
    .Y(net5753));
 BUFx6f_ASAP7_75t_R place5754 (.A(net5763),
    .Y(net5754));
 BUFx6f_ASAP7_75t_R place5755 (.A(net5763),
    .Y(net5755));
 BUFx3_ASAP7_75t_R place5756 (.A(net5763),
    .Y(net5756));
 BUFx3_ASAP7_75t_R place5757 (.A(net5763),
    .Y(net5757));
 BUFx3_ASAP7_75t_R place5758 (.A(net5763),
    .Y(net5758));
 BUFx6f_ASAP7_75t_R place5759 (.A(net5760),
    .Y(net5759));
 BUFx6f_ASAP7_75t_R place5760 (.A(net5763),
    .Y(net5760));
 BUFx3_ASAP7_75t_R place5761 (.A(net5763),
    .Y(net5761));
 BUFx3_ASAP7_75t_R place5762 (.A(net5763),
    .Y(net5762));
 BUFx6f_ASAP7_75t_R place5763 (.A(_14999_),
    .Y(net5763));
 BUFx6f_ASAP7_75t_R place5764 (.A(_14989_),
    .Y(net5764));
 BUFx3_ASAP7_75t_R place5765 (.A(net5767),
    .Y(net5765));
 BUFx3_ASAP7_75t_R place5766 (.A(net5767),
    .Y(net5766));
 BUFx3_ASAP7_75t_R place5767 (.A(_14989_),
    .Y(net5767));
 BUFx3_ASAP7_75t_R place5768 (.A(net5776),
    .Y(net5768));
 BUFx3_ASAP7_75t_R place5769 (.A(net5776),
    .Y(net5769));
 BUFx3_ASAP7_75t_R place5770 (.A(net5776),
    .Y(net5770));
 BUFx3_ASAP7_75t_R place5771 (.A(net5776),
    .Y(net5771));
 BUFx3_ASAP7_75t_R place5772 (.A(net5776),
    .Y(net5772));
 BUFx6f_ASAP7_75t_R place5773 (.A(net5776),
    .Y(net5773));
 BUFx3_ASAP7_75t_R place5774 (.A(net5776),
    .Y(net5774));
 BUFx3_ASAP7_75t_R place5775 (.A(net5776),
    .Y(net5775));
 BUFx6f_ASAP7_75t_R place5776 (.A(_14989_),
    .Y(net5776));
 BUFx3_ASAP7_75t_R place5777 (.A(_14972_),
    .Y(net5777));
 BUFx3_ASAP7_75t_R place5778 (.A(_14971_),
    .Y(net5778));
 BUFx3_ASAP7_75t_R place5779 (.A(_14956_),
    .Y(net5779));
 BUFx3_ASAP7_75t_R place5780 (.A(_14393_),
    .Y(net5780));
 BUFx3_ASAP7_75t_R place5781 (.A(_14393_),
    .Y(net5781));
 BUFx6f_ASAP7_75t_R place5782 (.A(_14393_),
    .Y(net5782));
 BUFx6f_ASAP7_75t_R place5783 (.A(net5784),
    .Y(net5783));
 BUFx6f_ASAP7_75t_R place5784 (.A(net5791),
    .Y(net5784));
 BUFx6f_ASAP7_75t_R place5785 (.A(net5791),
    .Y(net5785));
 BUFx3_ASAP7_75t_R place5786 (.A(net5791),
    .Y(net5786));
 BUFx3_ASAP7_75t_R place5787 (.A(net5791),
    .Y(net5787));
 BUFx3_ASAP7_75t_R place5788 (.A(net5791),
    .Y(net5788));
 BUFx3_ASAP7_75t_R place5789 (.A(net5791),
    .Y(net5789));
 BUFx6f_ASAP7_75t_R place5790 (.A(net5791),
    .Y(net5790));
 BUFx6f_ASAP7_75t_R place5791 (.A(_14346_),
    .Y(net5791));
 BUFx6f_ASAP7_75t_R place5792 (.A(_14338_),
    .Y(net5792));
 BUFx6f_ASAP7_75t_R place5793 (.A(_14323_),
    .Y(net5793));
 BUFx3_ASAP7_75t_R place5794 (.A(net5797),
    .Y(net5794));
 BUFx3_ASAP7_75t_R place5795 (.A(net5797),
    .Y(net5795));
 BUFx3_ASAP7_75t_R place5796 (.A(net5797),
    .Y(net5796));
 BUFx6f_ASAP7_75t_R place5797 (.A(_14323_),
    .Y(net5797));
 BUFx3_ASAP7_75t_R place5798 (.A(_14307_),
    .Y(net5798));
 BUFx6f_ASAP7_75t_R place5799 (.A(_14307_),
    .Y(net5799));
 BUFx6f_ASAP7_75t_R place5800 (.A(_14307_),
    .Y(net5800));
 BUFx3_ASAP7_75t_R place5801 (.A(net5810),
    .Y(net5801));
 BUFx3_ASAP7_75t_R place5802 (.A(net5810),
    .Y(net5802));
 BUFx3_ASAP7_75t_R place5803 (.A(net5810),
    .Y(net5803));
 BUFx6f_ASAP7_75t_R place5804 (.A(net5810),
    .Y(net5804));
 BUFx3_ASAP7_75t_R place5805 (.A(net5810),
    .Y(net5805));
 BUFx6f_ASAP7_75t_R place5806 (.A(net5810),
    .Y(net5806));
 BUFx3_ASAP7_75t_R place5807 (.A(net5810),
    .Y(net5807));
 BUFx3_ASAP7_75t_R place5808 (.A(net5810),
    .Y(net5808));
 BUFx6f_ASAP7_75t_R place5809 (.A(net5810),
    .Y(net5809));
 BUFx6f_ASAP7_75t_R place5810 (.A(_14287_),
    .Y(net5810));
 BUFx3_ASAP7_75t_R place5811 (.A(_14266_),
    .Y(net5811));
 BUFx3_ASAP7_75t_R place5812 (.A(net5813),
    .Y(net5812));
 BUFx6f_ASAP7_75t_R place5813 (.A(_14266_),
    .Y(net5813));
 BUFx3_ASAP7_75t_R place5814 (.A(_14266_),
    .Y(net5814));
 BUFx3_ASAP7_75t_R place5815 (.A(_14266_),
    .Y(net5815));
 BUFx3_ASAP7_75t_R place5816 (.A(_14266_),
    .Y(net5816));
 BUFx3_ASAP7_75t_R place5817 (.A(_14263_),
    .Y(net5817));
 BUFx6f_ASAP7_75t_R place5818 (.A(_14260_),
    .Y(net5818));
 BUFx3_ASAP7_75t_R place5819 (.A(_14260_),
    .Y(net5819));
 BUFx3_ASAP7_75t_R place5820 (.A(_14260_),
    .Y(net5820));
 BUFx6f_ASAP7_75t_R place5821 (.A(_14260_),
    .Y(net5821));
 BUFx3_ASAP7_75t_R place5822 (.A(_14242_),
    .Y(net5822));
 BUFx3_ASAP7_75t_R place5823 (.A(_14242_),
    .Y(net5823));
 BUFx3_ASAP7_75t_R place5824 (.A(_13759_),
    .Y(net5824));
 BUFx3_ASAP7_75t_R place5825 (.A(_13759_),
    .Y(net5825));
 BUFx3_ASAP7_75t_R place5826 (.A(_13759_),
    .Y(net5826));
 BUFx3_ASAP7_75t_R place5827 (.A(_13759_),
    .Y(net5827));
 BUFx6f_ASAP7_75t_R place5828 (.A(_13677_),
    .Y(net5828));
 BUFx3_ASAP7_75t_R place5829 (.A(net5834),
    .Y(net5829));
 BUFx6f_ASAP7_75t_R place5830 (.A(net5834),
    .Y(net5830));
 BUFx3_ASAP7_75t_R place5831 (.A(net5834),
    .Y(net5831));
 BUFx3_ASAP7_75t_R place5832 (.A(net5834),
    .Y(net5832));
 BUFx3_ASAP7_75t_R place5833 (.A(net5834),
    .Y(net5833));
 BUFx6f_ASAP7_75t_R place5834 (.A(_13612_),
    .Y(net5834));
 BUFx6f_ASAP7_75t_R place5835 (.A(net5840),
    .Y(net5835));
 BUFx6f_ASAP7_75t_R place5836 (.A(net5840),
    .Y(net5836));
 BUFx3_ASAP7_75t_R place5837 (.A(net5840),
    .Y(net5837));
 BUFx3_ASAP7_75t_R place5838 (.A(net5840),
    .Y(net5838));
 BUFx3_ASAP7_75t_R place5839 (.A(net5840),
    .Y(net5839));
 BUFx6f_ASAP7_75t_R place5840 (.A(_13595_),
    .Y(net5840));
 BUFx3_ASAP7_75t_R place5841 (.A(net5843),
    .Y(net5841));
 BUFx3_ASAP7_75t_R place5842 (.A(net5843),
    .Y(net5842));
 BUFx6f_ASAP7_75t_R place5843 (.A(_13595_),
    .Y(net5843));
 BUFx3_ASAP7_75t_R place5844 (.A(_13578_),
    .Y(net5844));
 BUFx3_ASAP7_75t_R place5845 (.A(_13567_),
    .Y(net5845));
 BUFx3_ASAP7_75t_R place5846 (.A(_01152_),
    .Y(net5846));
 BUFx3_ASAP7_75t_R place5847 (.A(_01152_),
    .Y(net5847));
 BUFx6f_ASAP7_75t_R place5848 (.A(_12966_),
    .Y(net5848));
 BUFx3_ASAP7_75t_R place5849 (.A(_12935_),
    .Y(net5849));
 BUFx3_ASAP7_75t_R place5850 (.A(_12935_),
    .Y(net5850));
 BUFx3_ASAP7_75t_R place5851 (.A(_12916_),
    .Y(net5851));
 BUFx3_ASAP7_75t_R place5852 (.A(_12916_),
    .Y(net5852));
 BUFx6f_ASAP7_75t_R place5853 (.A(_12916_),
    .Y(net5853));
 BUFx3_ASAP7_75t_R place5854 (.A(net5856),
    .Y(net5854));
 BUFx6f_ASAP7_75t_R place5855 (.A(net5856),
    .Y(net5855));
 BUFx6f_ASAP7_75t_R place5856 (.A(_12916_),
    .Y(net5856));
 BUFx6f_ASAP7_75t_R place5857 (.A(_12874_),
    .Y(net5857));
 BUFx6f_ASAP7_75t_R place5858 (.A(_12874_),
    .Y(net5858));
 BUFx3_ASAP7_75t_R place5859 (.A(_12870_),
    .Y(net5859));
 BUFx6f_ASAP7_75t_R place5860 (.A(_12866_),
    .Y(net5860));
 BUFx3_ASAP7_75t_R place5861 (.A(net5862),
    .Y(net5861));
 BUFx6f_ASAP7_75t_R place5862 (.A(_12866_),
    .Y(net5862));
 BUFx3_ASAP7_75t_R place5863 (.A(_12849_),
    .Y(net5863));
 BUFx3_ASAP7_75t_R place5864 (.A(_12832_),
    .Y(net5864));
 BUFx3_ASAP7_75t_R place5865 (.A(_12277_),
    .Y(net5865));
 BUFx3_ASAP7_75t_R place5866 (.A(_12245_),
    .Y(net5866));
 BUFx3_ASAP7_75t_R place5867 (.A(_12245_),
    .Y(net5867));
 BUFx6f_ASAP7_75t_R place5868 (.A(_12182_),
    .Y(net5868));
 BUFx3_ASAP7_75t_R place5869 (.A(_12182_),
    .Y(net5869));
 BUFx3_ASAP7_75t_R place5870 (.A(_12178_),
    .Y(net5870));
 BUFx3_ASAP7_75t_R place5871 (.A(_12172_),
    .Y(net5871));
 BUFx3_ASAP7_75t_R place5872 (.A(_01110_),
    .Y(net5872));
 BUFx3_ASAP7_75t_R place5873 (.A(_01110_),
    .Y(net5873));
 BUFx3_ASAP7_75t_R place5874 (.A(_12139_),
    .Y(net5874));
 BUFx3_ASAP7_75t_R place5875 (.A(_11576_),
    .Y(net5875));
 BUFx3_ASAP7_75t_R place5876 (.A(_11576_),
    .Y(net5876));
 BUFx3_ASAP7_75t_R place5877 (.A(net5878),
    .Y(net5877));
 BUFx3_ASAP7_75t_R place5878 (.A(_11553_),
    .Y(net5878));
 BUFx6f_ASAP7_75t_R place5879 (.A(_11519_),
    .Y(net5879));
 BUFx3_ASAP7_75t_R place5880 (.A(_11465_),
    .Y(net5880));
 BUFx3_ASAP7_75t_R place5881 (.A(_11448_),
    .Y(net5881));
 BUFx6f_ASAP7_75t_R place5882 (.A(_11446_),
    .Y(net5882));
 BUFx3_ASAP7_75t_R place5883 (.A(_11443_),
    .Y(net5883));
 BUFx3_ASAP7_75t_R place5884 (.A(_11443_),
    .Y(net5884));
 BUFx3_ASAP7_75t_R place5885 (.A(_11443_),
    .Y(net5885));
 BUFx3_ASAP7_75t_R place5886 (.A(_11443_),
    .Y(net5886));
 BUFx3_ASAP7_75t_R place5887 (.A(_11426_),
    .Y(net5887));
 BUFx3_ASAP7_75t_R place5888 (.A(_11426_),
    .Y(net5888));
 BUFx3_ASAP7_75t_R place5889 (.A(net5890),
    .Y(net5889));
 BUFx3_ASAP7_75t_R place5890 (.A(_11409_),
    .Y(net5890));
 BUFx3_ASAP7_75t_R place5891 (.A(_11409_),
    .Y(net5891));
 BUFx3_ASAP7_75t_R place5892 (.A(net5894),
    .Y(net5892));
 BUFx3_ASAP7_75t_R place5893 (.A(net5894),
    .Y(net5893));
 BUFx6f_ASAP7_75t_R place5894 (.A(_10835_),
    .Y(net5894));
 BUFx6f_ASAP7_75t_R place5895 (.A(_10753_),
    .Y(net5895));
 BUFx3_ASAP7_75t_R place5896 (.A(net5898),
    .Y(net5896));
 BUFx3_ASAP7_75t_R place5897 (.A(net5898),
    .Y(net5897));
 BUFx6f_ASAP7_75t_R place5898 (.A(_10741_),
    .Y(net5898));
 BUFx3_ASAP7_75t_R place5899 (.A(_10741_),
    .Y(net5899));
 BUFx3_ASAP7_75t_R place5900 (.A(net5901),
    .Y(net5900));
 BUFx3_ASAP7_75t_R place5901 (.A(_10736_),
    .Y(net5901));
 BUFx6f_ASAP7_75t_R place5902 (.A(net5905),
    .Y(net5902));
 BUFx6f_ASAP7_75t_R place5903 (.A(net5905),
    .Y(net5903));
 BUFx3_ASAP7_75t_R place5904 (.A(net5905),
    .Y(net5904));
 BUFx6f_ASAP7_75t_R place5905 (.A(_10732_),
    .Y(net5905));
 BUFx3_ASAP7_75t_R place5906 (.A(_10715_),
    .Y(net5906));
 BUFx3_ASAP7_75t_R place5907 (.A(_10715_),
    .Y(net5907));
 BUFx3_ASAP7_75t_R place5908 (.A(_10695_),
    .Y(net5908));
 BUFx3_ASAP7_75t_R place5909 (.A(_10695_),
    .Y(net5909));
 BUFx3_ASAP7_75t_R place5910 (.A(_10695_),
    .Y(net5910));
 BUFx3_ASAP7_75t_R place5911 (.A(_10140_),
    .Y(net5911));
 BUFx3_ASAP7_75t_R place5912 (.A(net5916),
    .Y(net5912));
 BUFx3_ASAP7_75t_R place5913 (.A(net5916),
    .Y(net5913));
 BUFx3_ASAP7_75t_R place5914 (.A(net5916),
    .Y(net5914));
 BUFx3_ASAP7_75t_R place5915 (.A(net5916),
    .Y(net5915));
 BUFx6f_ASAP7_75t_R place5916 (.A(_10140_),
    .Y(net5916));
 BUFx3_ASAP7_75t_R place5917 (.A(_10140_),
    .Y(net5917));
 BUFx3_ASAP7_75t_R place5918 (.A(_09688_),
    .Y(net5918));
 BUFx3_ASAP7_75t_R place5919 (.A(net5920),
    .Y(net5919));
 BUFx6f_ASAP7_75t_R place5920 (.A(_09594_),
    .Y(net5920));
 BUFx3_ASAP7_75t_R place5921 (.A(_09580_),
    .Y(net5921));
 BUFx3_ASAP7_75t_R place5922 (.A(_09187_),
    .Y(net5922));
 BUFx3_ASAP7_75t_R place5923 (.A(_09151_),
    .Y(net5923));
 BUFx3_ASAP7_75t_R place5924 (.A(_09124_),
    .Y(net5924));
 BUFx3_ASAP7_75t_R place5925 (.A(_09043_),
    .Y(net5925));
 BUFx6f_ASAP7_75t_R place5926 (.A(_09043_),
    .Y(net5926));
 BUFx3_ASAP7_75t_R place5927 (.A(_09043_),
    .Y(net5927));
 BUFx3_ASAP7_75t_R place5928 (.A(_09043_),
    .Y(net5928));
 BUFx3_ASAP7_75t_R place5929 (.A(_09043_),
    .Y(net5929));
 BUFx3_ASAP7_75t_R place5930 (.A(_09043_),
    .Y(net5930));
 BUFx3_ASAP7_75t_R place5931 (.A(_00995_),
    .Y(net5931));
 BUFx3_ASAP7_75t_R place5932 (.A(_09030_),
    .Y(net5932));
 BUFx6f_ASAP7_75t_R place5933 (.A(_09026_),
    .Y(net5933));
 BUFx3_ASAP7_75t_R place5934 (.A(_09016_),
    .Y(net5934));
 BUFx6f_ASAP7_75t_R place5935 (.A(net5937),
    .Y(net5935));
 BUFx6f_ASAP7_75t_R place5936 (.A(net5937),
    .Y(net5936));
 BUFx6f_ASAP7_75t_R place5937 (.A(_09016_),
    .Y(net5937));
 BUFx3_ASAP7_75t_R place5938 (.A(_09007_),
    .Y(net5938));
 BUFx3_ASAP7_75t_R place5939 (.A(_09007_),
    .Y(net5939));
 BUFx3_ASAP7_75t_R place5940 (.A(_01047_),
    .Y(net5940));
 BUFx3_ASAP7_75t_R place5941 (.A(_01047_),
    .Y(net5941));
 BUFx3_ASAP7_75t_R place5942 (.A(_08984_),
    .Y(net5942));
 BUFx6f_ASAP7_75t_R place5943 (.A(_08980_),
    .Y(net5943));
 BUFx6f_ASAP7_75t_R place5944 (.A(net5945),
    .Y(net5944));
 BUFx6f_ASAP7_75t_R place5945 (.A(_08968_),
    .Y(net5945));
 BUFx3_ASAP7_75t_R place5946 (.A(_08968_),
    .Y(net5946));
 BUFx3_ASAP7_75t_R place5947 (.A(net5948),
    .Y(net5947));
 BUFx6f_ASAP7_75t_R place5948 (.A(_08968_),
    .Y(net5948));
 BUFx3_ASAP7_75t_R place5949 (.A(_08962_),
    .Y(net5949));
 BUFx3_ASAP7_75t_R place5950 (.A(_08962_),
    .Y(net5950));
 BUFx3_ASAP7_75t_R place5951 (.A(_08962_),
    .Y(net5951));
 BUFx3_ASAP7_75t_R place5952 (.A(_01000_),
    .Y(net5952));
 BUFx3_ASAP7_75t_R place5953 (.A(_08944_),
    .Y(net5953));
 BUFx3_ASAP7_75t_R place5954 (.A(_08940_),
    .Y(net5954));
 BUFx6f_ASAP7_75t_R place5955 (.A(net5957),
    .Y(net5955));
 BUFx3_ASAP7_75t_R place5956 (.A(net5957),
    .Y(net5956));
 BUFx6f_ASAP7_75t_R place5957 (.A(_08929_),
    .Y(net5957));
 BUFx3_ASAP7_75t_R place5958 (.A(_08929_),
    .Y(net5958));
 BUFx6f_ASAP7_75t_R place5959 (.A(net5960),
    .Y(net5959));
 BUFx6f_ASAP7_75t_R place5960 (.A(_08929_),
    .Y(net5960));
 BUFx3_ASAP7_75t_R place5961 (.A(net5962),
    .Y(net5961));
 BUFx6f_ASAP7_75t_R place5962 (.A(_08929_),
    .Y(net5962));
 BUFx3_ASAP7_75t_R place5963 (.A(_08923_),
    .Y(net5963));
 BUFx3_ASAP7_75t_R place5964 (.A(_08923_),
    .Y(net5964));
 BUFx3_ASAP7_75t_R place5965 (.A(net5966),
    .Y(net5965));
 BUFx3_ASAP7_75t_R place5966 (.A(_01025_),
    .Y(net5966));
 BUFx3_ASAP7_75t_R place5967 (.A(_08233_),
    .Y(net5967));
 BUFx6f_ASAP7_75t_R place5968 (.A(_08215_),
    .Y(net5968));
 BUFx3_ASAP7_75t_R place5969 (.A(net5970),
    .Y(net5969));
 BUFx6f_ASAP7_75t_R place5970 (.A(_08193_),
    .Y(net5970));
 BUFx3_ASAP7_75t_R place5971 (.A(_08172_),
    .Y(net5971));
 BUFx6f_ASAP7_75t_R place5972 (.A(_08169_),
    .Y(net5972));
 BUFx3_ASAP7_75t_R place5973 (.A(_08130_),
    .Y(net5973));
 BUFx3_ASAP7_75t_R place5974 (.A(_08127_),
    .Y(net5974));
 BUFx3_ASAP7_75t_R place5975 (.A(_08121_),
    .Y(net5975));
 BUFx3_ASAP7_75t_R place5976 (.A(_08117_),
    .Y(net5976));
 BUFx3_ASAP7_75t_R place5977 (.A(_08117_),
    .Y(net5977));
 BUFx6f_ASAP7_75t_R place5978 (.A(net5980),
    .Y(net5978));
 BUFx6f_ASAP7_75t_R place5979 (.A(net5980),
    .Y(net5979));
 BUFx6f_ASAP7_75t_R place5980 (.A(_08117_),
    .Y(net5980));
 BUFx3_ASAP7_75t_R place5981 (.A(_00973_),
    .Y(net5981));
 BUFx3_ASAP7_75t_R place5982 (.A(_00972_),
    .Y(net5982));
 BUFx3_ASAP7_75t_R place5983 (.A(_00972_),
    .Y(net5983));
 BUFx3_ASAP7_75t_R place5984 (.A(_07251_),
    .Y(net5984));
 BUFx6f_ASAP7_75t_R place5985 (.A(_07242_),
    .Y(net5985));
 BUFx3_ASAP7_75t_R place5986 (.A(_07234_),
    .Y(net5986));
 BUFx6f_ASAP7_75t_R place5987 (.A(_07234_),
    .Y(net5987));
 BUFx6f_ASAP7_75t_R place5988 (.A(_07224_),
    .Y(net5988));
 BUFx6f_ASAP7_75t_R place5989 (.A(_07224_),
    .Y(net5989));
 BUFx3_ASAP7_75t_R place5990 (.A(_07224_),
    .Y(net5990));
 BUFx3_ASAP7_75t_R place5991 (.A(_07224_),
    .Y(net5991));
 BUFx3_ASAP7_75t_R place5992 (.A(_07194_),
    .Y(net5992));
 BUFx3_ASAP7_75t_R place5993 (.A(_07194_),
    .Y(net5993));
 BUFx6f_ASAP7_75t_R place5994 (.A(_07179_),
    .Y(net5994));
 BUFx3_ASAP7_75t_R place5995 (.A(net5996),
    .Y(net5995));
 BUFx6f_ASAP7_75t_R place5996 (.A(_07179_),
    .Y(net5996));
 BUFx6f_ASAP7_75t_R place5997 (.A(_07179_),
    .Y(net5997));
 BUFx6f_ASAP7_75t_R place5998 (.A(_07171_),
    .Y(net5998));
 BUFx3_ASAP7_75t_R place5999 (.A(_07171_),
    .Y(net5999));
 BUFx3_ASAP7_75t_R place6000 (.A(_07171_),
    .Y(net6000));
 BUFx3_ASAP7_75t_R place6001 (.A(_07171_),
    .Y(net6001));
 BUFx6f_ASAP7_75t_R place6002 (.A(_07171_),
    .Y(net6002));
 BUFx6f_ASAP7_75t_R place6003 (.A(_07171_),
    .Y(net6003));
 BUFx6f_ASAP7_75t_R place6004 (.A(net6007),
    .Y(net6004));
 BUFx3_ASAP7_75t_R place6005 (.A(net6007),
    .Y(net6005));
 BUFx3_ASAP7_75t_R place6006 (.A(net6007),
    .Y(net6006));
 BUFx6f_ASAP7_75t_R place6007 (.A(_07166_),
    .Y(net6007));
 BUFx3_ASAP7_75t_R place6008 (.A(net6009),
    .Y(net6008));
 BUFx6f_ASAP7_75t_R place6009 (.A(_07166_),
    .Y(net6009));
 BUFx3_ASAP7_75t_R place6010 (.A(_07156_),
    .Y(net6010));
 BUFx3_ASAP7_75t_R place6011 (.A(_07155_),
    .Y(net6011));
 BUFx3_ASAP7_75t_R place6012 (.A(_07151_),
    .Y(net6012));
 BUFx3_ASAP7_75t_R place6013 (.A(_07150_),
    .Y(net6013));
 BUFx3_ASAP7_75t_R place6014 (.A(_06630_),
    .Y(net6014));
 BUFx3_ASAP7_75t_R place6015 (.A(_06529_),
    .Y(net6015));
 BUFx6f_ASAP7_75t_R place6016 (.A(_06529_),
    .Y(net6016));
 BUFx3_ASAP7_75t_R place6017 (.A(_06529_),
    .Y(net6017));
 BUFx3_ASAP7_75t_R place6018 (.A(_06522_),
    .Y(net6018));
 BUFx3_ASAP7_75t_R place6019 (.A(net6021),
    .Y(net6019));
 BUFx3_ASAP7_75t_R place6020 (.A(net6021),
    .Y(net6020));
 BUFx6f_ASAP7_75t_R place6021 (.A(_06522_),
    .Y(net6021));
 BUFx6f_ASAP7_75t_R place6022 (.A(net6023),
    .Y(net6022));
 BUFx6f_ASAP7_75t_R place6023 (.A(_06522_),
    .Y(net6023));
 BUFx3_ASAP7_75t_R place6024 (.A(_06522_),
    .Y(net6024));
 BUFx3_ASAP7_75t_R place6025 (.A(_06514_),
    .Y(net6025));
 BUFx6f_ASAP7_75t_R place6026 (.A(net6031),
    .Y(net6026));
 BUFx3_ASAP7_75t_R place6027 (.A(net6031),
    .Y(net6027));
 BUFx3_ASAP7_75t_R place6028 (.A(net6031),
    .Y(net6028));
 BUFx6f_ASAP7_75t_R place6029 (.A(net6031),
    .Y(net6029));
 BUFx6f_ASAP7_75t_R place6030 (.A(net6031),
    .Y(net6030));
 BUFx6f_ASAP7_75t_R place6031 (.A(_06514_),
    .Y(net6031));
 BUFx3_ASAP7_75t_R place6032 (.A(_06502_),
    .Y(net6032));
 BUFx3_ASAP7_75t_R place6033 (.A(_06494_),
    .Y(net6033));
 BUFx3_ASAP7_75t_R place6034 (.A(_06493_),
    .Y(net6034));
 BUFx3_ASAP7_75t_R place6035 (.A(_06487_),
    .Y(net6035));
 BUFx3_ASAP7_75t_R place6036 (.A(_06486_),
    .Y(net6036));
 BUFx3_ASAP7_75t_R place6037 (.A(_06469_),
    .Y(net6037));
 BUFx3_ASAP7_75t_R place6038 (.A(_05955_),
    .Y(net6038));
 BUFx3_ASAP7_75t_R place6039 (.A(_05879_),
    .Y(net6039));
 BUFx3_ASAP7_75t_R place6040 (.A(net6041),
    .Y(net6040));
 BUFx6f_ASAP7_75t_R place6041 (.A(_05853_),
    .Y(net6041));
 BUFx6f_ASAP7_75t_R place6042 (.A(_05853_),
    .Y(net6042));
 BUFx6f_ASAP7_75t_R place6043 (.A(net6044),
    .Y(net6043));
 BUFx3_ASAP7_75t_R place6044 (.A(_05853_),
    .Y(net6044));
 BUFx6f_ASAP7_75t_R place6045 (.A(_05838_),
    .Y(net6045));
 BUFx3_ASAP7_75t_R place6046 (.A(net6049),
    .Y(net6046));
 BUFx3_ASAP7_75t_R place6047 (.A(net6049),
    .Y(net6047));
 BUFx3_ASAP7_75t_R place6048 (.A(net6049),
    .Y(net6048));
 BUFx6f_ASAP7_75t_R place6049 (.A(_05817_),
    .Y(net6049));
 BUFx3_ASAP7_75t_R place6050 (.A(net6052),
    .Y(net6050));
 BUFx3_ASAP7_75t_R place6051 (.A(net6052),
    .Y(net6051));
 BUFx6f_ASAP7_75t_R place6052 (.A(_05817_),
    .Y(net6052));
 BUFx3_ASAP7_75t_R place6053 (.A(_05804_),
    .Y(net6053));
 BUFx3_ASAP7_75t_R place6054 (.A(_05803_),
    .Y(net6054));
 BUFx3_ASAP7_75t_R place6055 (.A(_05799_),
    .Y(net6055));
 BUFx3_ASAP7_75t_R place6056 (.A(_05794_),
    .Y(net6056));
 BUFx3_ASAP7_75t_R place6057 (.A(_05792_),
    .Y(net6057));
 BUFx3_ASAP7_75t_R place6058 (.A(_05791_),
    .Y(net6058));
 BUFx3_ASAP7_75t_R place6059 (.A(_05276_),
    .Y(net6059));
 BUFx3_ASAP7_75t_R place6060 (.A(_05218_),
    .Y(net6060));
 BUFx6f_ASAP7_75t_R place6061 (.A(net6065),
    .Y(net6061));
 BUFx6f_ASAP7_75t_R place6062 (.A(net6065),
    .Y(net6062));
 BUFx3_ASAP7_75t_R place6063 (.A(net6065),
    .Y(net6063));
 BUFx3_ASAP7_75t_R place6064 (.A(net6065),
    .Y(net6064));
 BUFx6f_ASAP7_75t_R place6065 (.A(_05170_),
    .Y(net6065));
 BUFx3_ASAP7_75t_R place6066 (.A(_05170_),
    .Y(net6066));
 BUFx3_ASAP7_75t_R place6067 (.A(_05170_),
    .Y(net6067));
 BUFx6f_ASAP7_75t_R place6068 (.A(_05157_),
    .Y(net6068));
 BUFx3_ASAP7_75t_R place6069 (.A(_05157_),
    .Y(net6069));
 BUFx3_ASAP7_75t_R place6070 (.A(_05157_),
    .Y(net6070));
 BUFx6f_ASAP7_75t_R place6071 (.A(_05157_),
    .Y(net6071));
 BUFx3_ASAP7_75t_R place6072 (.A(_05147_),
    .Y(net6072));
 BUFx6f_ASAP7_75t_R place6073 (.A(_05147_),
    .Y(net6073));
 BUFx6f_ASAP7_75t_R place6074 (.A(_05147_),
    .Y(net6074));
 BUFx6f_ASAP7_75t_R place6075 (.A(_05147_),
    .Y(net6075));
 BUFx3_ASAP7_75t_R place6076 (.A(net6077),
    .Y(net6076));
 BUFx6f_ASAP7_75t_R place6077 (.A(_05140_),
    .Y(net6077));
 BUFx3_ASAP7_75t_R place6078 (.A(net6082),
    .Y(net6078));
 BUFx6f_ASAP7_75t_R place6079 (.A(net6082),
    .Y(net6079));
 BUFx3_ASAP7_75t_R place6080 (.A(net6082),
    .Y(net6080));
 BUFx6f_ASAP7_75t_R place6081 (.A(net6082),
    .Y(net6081));
 BUFx6f_ASAP7_75t_R place6082 (.A(_05140_),
    .Y(net6082));
 BUFx3_ASAP7_75t_R place6083 (.A(_05126_),
    .Y(net6083));
 BUFx3_ASAP7_75t_R place6084 (.A(_05125_),
    .Y(net6084));
 BUFx3_ASAP7_75t_R place6085 (.A(_05118_),
    .Y(net6085));
 BUFx3_ASAP7_75t_R place6086 (.A(_05117_),
    .Y(net6086));
 BUFx3_ASAP7_75t_R place6087 (.A(_05100_),
    .Y(net6087));
 BUFx3_ASAP7_75t_R place6088 (.A(_04578_),
    .Y(net6088));
 BUFx3_ASAP7_75t_R place6089 (.A(_04535_),
    .Y(net6089));
 BUFx3_ASAP7_75t_R place6090 (.A(_04499_),
    .Y(net6090));
 BUFx6f_ASAP7_75t_R place6091 (.A(net6094),
    .Y(net6091));
 BUFx3_ASAP7_75t_R place6092 (.A(net6094),
    .Y(net6092));
 BUFx3_ASAP7_75t_R place6093 (.A(net6094),
    .Y(net6093));
 BUFx6f_ASAP7_75t_R place6094 (.A(_04485_),
    .Y(net6094));
 BUFx3_ASAP7_75t_R place6095 (.A(net6099),
    .Y(net6095));
 BUFx3_ASAP7_75t_R place6096 (.A(net6099),
    .Y(net6096));
 BUFx3_ASAP7_75t_R place6097 (.A(net6099),
    .Y(net6097));
 BUFx3_ASAP7_75t_R place6098 (.A(net6099),
    .Y(net6098));
 BUFx6f_ASAP7_75t_R place6099 (.A(_04485_),
    .Y(net6099));
 BUFx3_ASAP7_75t_R place6100 (.A(net6101),
    .Y(net6100));
 BUFx6f_ASAP7_75t_R place6101 (.A(_04468_),
    .Y(net6101));
 BUFx3_ASAP7_75t_R place6102 (.A(_04444_),
    .Y(net6102));
 BUFx3_ASAP7_75t_R place6103 (.A(net6105),
    .Y(net6103));
 BUFx3_ASAP7_75t_R place6104 (.A(net6105),
    .Y(net6104));
 BUFx6f_ASAP7_75t_R place6105 (.A(_04444_),
    .Y(net6105));
 BUFx3_ASAP7_75t_R place6106 (.A(net6107),
    .Y(net6106));
 BUFx6f_ASAP7_75t_R place6107 (.A(_04444_),
    .Y(net6107));
 BUFx3_ASAP7_75t_R place6108 (.A(_03823_),
    .Y(net6108));
 BUFx6f_ASAP7_75t_R place6109 (.A(_03798_),
    .Y(net6109));
 BUFx3_ASAP7_75t_R place6110 (.A(_03798_),
    .Y(net6110));
 BUFx6f_ASAP7_75t_R place6111 (.A(net6115),
    .Y(net6111));
 BUFx3_ASAP7_75t_R place6112 (.A(net6115),
    .Y(net6112));
 BUFx6f_ASAP7_75t_R place6113 (.A(net6114),
    .Y(net6113));
 BUFx6f_ASAP7_75t_R place6114 (.A(net6115),
    .Y(net6114));
 BUFx6f_ASAP7_75t_R place6115 (.A(_03798_),
    .Y(net6115));
 BUFx3_ASAP7_75t_R place6116 (.A(_03788_),
    .Y(net6116));
 BUFx3_ASAP7_75t_R place6117 (.A(_03764_),
    .Y(net6117));
 BUFx6f_ASAP7_75t_R place6118 (.A(_03756_),
    .Y(net6118));
 BUFx3_ASAP7_75t_R place6119 (.A(_03756_),
    .Y(net6119));
 BUFx3_ASAP7_75t_R place6120 (.A(_03756_),
    .Y(net6120));
 BUFx3_ASAP7_75t_R place6121 (.A(net6122),
    .Y(net6121));
 BUFx6f_ASAP7_75t_R place6122 (.A(_03756_),
    .Y(net6122));
 BUFx6f_ASAP7_75t_R place6123 (.A(_03752_),
    .Y(net6123));
 BUFx6f_ASAP7_75t_R place6124 (.A(_03752_),
    .Y(net6124));
 BUFx3_ASAP7_75t_R place6125 (.A(_03752_),
    .Y(net6125));
 BUFx6f_ASAP7_75t_R place6126 (.A(_03752_),
    .Y(net6126));
 BUFx3_ASAP7_75t_R place6127 (.A(_03752_),
    .Y(net6127));
 BUFx6f_ASAP7_75t_R place6128 (.A(net6132),
    .Y(net6128));
 BUFx3_ASAP7_75t_R place6129 (.A(net6132),
    .Y(net6129));
 BUFx3_ASAP7_75t_R place6130 (.A(net6132),
    .Y(net6130));
 BUFx3_ASAP7_75t_R place6131 (.A(net6132),
    .Y(net6131));
 BUFx6f_ASAP7_75t_R place6132 (.A(_03731_),
    .Y(net6132));
 BUFx6f_ASAP7_75t_R place6133 (.A(net6136),
    .Y(net6133));
 BUFx3_ASAP7_75t_R place6134 (.A(net6136),
    .Y(net6134));
 BUFx3_ASAP7_75t_R place6135 (.A(net6136),
    .Y(net6135));
 BUFx6f_ASAP7_75t_R place6136 (.A(_03731_),
    .Y(net6136));
 BUFx3_ASAP7_75t_R place6137 (.A(_03719_),
    .Y(net6137));
 BUFx3_ASAP7_75t_R place6138 (.A(_03717_),
    .Y(net6138));
 BUFx3_ASAP7_75t_R place6139 (.A(_03712_),
    .Y(net6139));
 BUFx3_ASAP7_75t_R place6140 (.A(_03694_),
    .Y(net6140));
 BUFx3_ASAP7_75t_R place6141 (.A(_03174_),
    .Y(net6141));
 BUFx3_ASAP7_75t_R place6142 (.A(_03103_),
    .Y(net6142));
 BUFx3_ASAP7_75t_R place6143 (.A(net6144),
    .Y(net6143));
 BUFx6f_ASAP7_75t_R place6144 (.A(_03065_),
    .Y(net6144));
 BUFx3_ASAP7_75t_R place6145 (.A(_03065_),
    .Y(net6145));
 BUFx3_ASAP7_75t_R place6146 (.A(net6150),
    .Y(net6146));
 BUFx6f_ASAP7_75t_R place6147 (.A(net6150),
    .Y(net6147));
 BUFx3_ASAP7_75t_R place6148 (.A(net6150),
    .Y(net6148));
 BUFx3_ASAP7_75t_R place6149 (.A(net6150),
    .Y(net6149));
 BUFx6f_ASAP7_75t_R place6150 (.A(_03055_),
    .Y(net6150));
 BUFx3_ASAP7_75t_R place6151 (.A(net6152),
    .Y(net6151));
 BUFx6f_ASAP7_75t_R place6152 (.A(_03055_),
    .Y(net6152));
 BUFx6f_ASAP7_75t_R place6153 (.A(_03050_),
    .Y(net6153));
 BUFx3_ASAP7_75t_R place6154 (.A(net6155),
    .Y(net6154));
 BUFx6f_ASAP7_75t_R place6155 (.A(_03050_),
    .Y(net6155));
 BUFx3_ASAP7_75t_R place6156 (.A(_03039_),
    .Y(net6156));
 BUFx3_ASAP7_75t_R place6157 (.A(_03034_),
    .Y(net6157));
 BUFx3_ASAP7_75t_R place6158 (.A(_03030_),
    .Y(net6158));
 BUFx3_ASAP7_75t_R place6159 (.A(_03010_),
    .Y(net6159));
 BUFx3_ASAP7_75t_R place6160 (.A(_02995_),
    .Y(net6160));
 BUFx3_ASAP7_75t_R place6161 (.A(_02990_),
    .Y(net6161));
 BUFx24_ASAP7_75t_R place6162 (.A(_02356_),
    .Y(net6162));
 BUFx3_ASAP7_75t_R place6163 (.A(_02348_),
    .Y(net6163));
 BUFx3_ASAP7_75t_R place6164 (.A(_02340_),
    .Y(net6164));
 BUFx3_ASAP7_75t_R place6165 (.A(_02335_),
    .Y(net6165));
 BUFx3_ASAP7_75t_R place6166 (.A(_02311_),
    .Y(net6166));
 BUFx3_ASAP7_75t_R place6167 (.A(_01779_),
    .Y(net6167));
 BUFx3_ASAP7_75t_R place6168 (.A(_01732_),
    .Y(net6168));
 BUFx3_ASAP7_75t_R place6169 (.A(_01638_),
    .Y(net6169));
 BUFx3_ASAP7_75t_R place6170 (.A(_01633_),
    .Y(net6170));
 BUFx3_ASAP7_75t_R place6171 (.A(_01613_),
    .Y(net6171));
 BUFx3_ASAP7_75t_R place6172 (.A(_15161_),
    .Y(net6172));
 BUFx3_ASAP7_75t_R place6173 (.A(_15137_),
    .Y(net6173));
 BUFx3_ASAP7_75t_R place6174 (.A(_15079_),
    .Y(net6174));
 BUFx3_ASAP7_75t_R place6175 (.A(_14997_),
    .Y(net6175));
 BUFx3_ASAP7_75t_R place6176 (.A(_14973_),
    .Y(net6176));
 BUFx3_ASAP7_75t_R place6177 (.A(_14966_),
    .Y(net6177));
 BUFx3_ASAP7_75t_R place6178 (.A(_14927_),
    .Y(net6178));
 BUFx3_ASAP7_75t_R place6179 (.A(_14927_),
    .Y(net6179));
 BUFx3_ASAP7_75t_R place6180 (.A(_14415_),
    .Y(net6180));
 BUFx3_ASAP7_75t_R place6181 (.A(_14368_),
    .Y(net6181));
 BUFx3_ASAP7_75t_R place6182 (.A(_14286_),
    .Y(net6182));
 BUFx3_ASAP7_75t_R place6183 (.A(_14285_),
    .Y(net6183));
 BUFx3_ASAP7_75t_R place6184 (.A(net6185),
    .Y(net6184));
 BUFx3_ASAP7_75t_R place6185 (.A(_14272_),
    .Y(net6185));
 BUFx3_ASAP7_75t_R place6186 (.A(_14265_),
    .Y(net6186));
 BUFx3_ASAP7_75t_R place6187 (.A(_14264_),
    .Y(net6187));
 BUFx3_ASAP7_75t_R place6188 (.A(_14259_),
    .Y(net6188));
 BUFx3_ASAP7_75t_R place6189 (.A(_14252_),
    .Y(net6189));
 BUFx3_ASAP7_75t_R place6190 (.A(_14224_),
    .Y(net6190));
 BUFx3_ASAP7_75t_R place6191 (.A(_14224_),
    .Y(net6191));
 BUFx3_ASAP7_75t_R place6192 (.A(_13724_),
    .Y(net6192));
 BUFx3_ASAP7_75t_R place6193 (.A(_13634_),
    .Y(net6193));
 BUFx3_ASAP7_75t_R place6194 (.A(_13628_),
    .Y(net6194));
 BUFx3_ASAP7_75t_R place6195 (.A(_13579_),
    .Y(net6195));
 BUFx3_ASAP7_75t_R place6196 (.A(_13570_),
    .Y(net6196));
 BUFx6f_ASAP7_75t_R place6197 (.A(net6198),
    .Y(net6197));
 BUFx3_ASAP7_75t_R place6198 (.A(_13533_),
    .Y(net6198));
 BUFx3_ASAP7_75t_R place6199 (.A(_13010_),
    .Y(net6199));
 BUFx3_ASAP7_75t_R place6200 (.A(_12934_),
    .Y(net6200));
 BUFx3_ASAP7_75t_R place6201 (.A(net6202),
    .Y(net6201));
 BUFx6f_ASAP7_75t_R place6202 (.A(_12921_),
    .Y(net6202));
 BUFx3_ASAP7_75t_R place6203 (.A(net6204),
    .Y(net6203));
 BUFx6f_ASAP7_75t_R place6204 (.A(_12921_),
    .Y(net6204));
 BUFx3_ASAP7_75t_R place6205 (.A(net6206),
    .Y(net6205));
 BUFx6f_ASAP7_75t_R place6206 (.A(_12921_),
    .Y(net6206));
 BUFx24_ASAP7_75t_R place6207 (.A(_12915_),
    .Y(net6207));
 BUFx3_ASAP7_75t_R place6208 (.A(net6211),
    .Y(net6208));
 BUFx3_ASAP7_75t_R place6209 (.A(net6211),
    .Y(net6209));
 BUFx3_ASAP7_75t_R place6210 (.A(net6211),
    .Y(net6210));
 BUFx6f_ASAP7_75t_R place6211 (.A(_12894_),
    .Y(net6211));
 BUFx3_ASAP7_75t_R place6212 (.A(_12894_),
    .Y(net6212));
 BUFx6f_ASAP7_75t_R place6213 (.A(_12894_),
    .Y(net6213));
 BUFx3_ASAP7_75t_R place6214 (.A(_12894_),
    .Y(net6214));
 BUFx3_ASAP7_75t_R place6215 (.A(_12873_),
    .Y(net6215));
 BUFx3_ASAP7_75t_R place6216 (.A(_12872_),
    .Y(net6216));
 BUFx3_ASAP7_75t_R place6217 (.A(_12865_),
    .Y(net6217));
 BUFx3_ASAP7_75t_R place6218 (.A(_12864_),
    .Y(net6218));
 BUFx3_ASAP7_75t_R place6219 (.A(_12848_),
    .Y(net6219));
 BUFx3_ASAP7_75t_R place6220 (.A(_12326_),
    .Y(net6220));
 BUFx3_ASAP7_75t_R place6221 (.A(_12276_),
    .Y(net6221));
 BUFx3_ASAP7_75t_R place6222 (.A(_12244_),
    .Y(net6222));
 BUFx3_ASAP7_75t_R place6223 (.A(_12244_),
    .Y(net6223));
 BUFx6f_ASAP7_75t_R place6224 (.A(_12232_),
    .Y(net6224));
 BUFx3_ASAP7_75t_R place6225 (.A(_12232_),
    .Y(net6225));
 BUFx6f_ASAP7_75t_R place6226 (.A(_12232_),
    .Y(net6226));
 BUFx6f_ASAP7_75t_R place6227 (.A(_12220_),
    .Y(net6227));
 BUFx3_ASAP7_75t_R place6228 (.A(_12220_),
    .Y(net6228));
 BUFx6f_ASAP7_75t_R place6229 (.A(_12220_),
    .Y(net6229));
 BUFx6f_ASAP7_75t_R place6230 (.A(net6231),
    .Y(net6230));
 BUFx6f_ASAP7_75t_R place6231 (.A(_12208_),
    .Y(net6231));
 BUFx3_ASAP7_75t_R place6232 (.A(_12208_),
    .Y(net6232));
 BUFx6f_ASAP7_75t_R place6233 (.A(_12208_),
    .Y(net6233));
 BUFx3_ASAP7_75t_R place6234 (.A(_12201_),
    .Y(net6234));
 BUFx3_ASAP7_75t_R place6235 (.A(_12201_),
    .Y(net6235));
 BUFx3_ASAP7_75t_R place6236 (.A(_12201_),
    .Y(net6236));
 BUFx3_ASAP7_75t_R place6237 (.A(net6238),
    .Y(net6237));
 BUFx6f_ASAP7_75t_R place6238 (.A(_12201_),
    .Y(net6238));
 BUFx3_ASAP7_75t_R place6239 (.A(_12181_),
    .Y(net6239));
 BUFx3_ASAP7_75t_R place6240 (.A(_12180_),
    .Y(net6240));
 BUFx3_ASAP7_75t_R place6241 (.A(_12173_),
    .Y(net6241));
 BUFx3_ASAP7_75t_R place6242 (.A(_11552_),
    .Y(net6242));
 BUFx3_ASAP7_75t_R place6243 (.A(_11551_),
    .Y(net6243));
 BUFx6f_ASAP7_75t_R place6244 (.A(_11528_),
    .Y(net6244));
 BUFx6f_ASAP7_75t_R place6245 (.A(_11528_),
    .Y(net6245));
 BUFx3_ASAP7_75t_R place6246 (.A(_11528_),
    .Y(net6246));
 BUFx6f_ASAP7_75t_R place6247 (.A(_11523_),
    .Y(net6247));
 BUFx6f_ASAP7_75t_R place6248 (.A(_11523_),
    .Y(net6248));
 BUFx6f_ASAP7_75t_R place6249 (.A(_11490_),
    .Y(net6249));
 BUFx3_ASAP7_75t_R place6250 (.A(_11490_),
    .Y(net6250));
 BUFx3_ASAP7_75t_R place6251 (.A(net6252),
    .Y(net6251));
 BUFx6f_ASAP7_75t_R place6252 (.A(_11477_),
    .Y(net6252));
 BUFx3_ASAP7_75t_R place6253 (.A(net6256),
    .Y(net6253));
 BUFx6f_ASAP7_75t_R place6254 (.A(net6256),
    .Y(net6254));
 BUFx3_ASAP7_75t_R place6255 (.A(net6256),
    .Y(net6255));
 BUFx6f_ASAP7_75t_R place6256 (.A(_11477_),
    .Y(net6256));
 BUFx3_ASAP7_75t_R place6257 (.A(_11464_),
    .Y(net6257));
 BUFx3_ASAP7_75t_R place6258 (.A(_11450_),
    .Y(net6258));
 BUFx3_ASAP7_75t_R place6259 (.A(_11442_),
    .Y(net6259));
 BUFx3_ASAP7_75t_R place6260 (.A(_11441_),
    .Y(net6260));
 BUFx3_ASAP7_75t_R place6261 (.A(_11408_),
    .Y(net6261));
 BUFx3_ASAP7_75t_R place6262 (.A(_11403_),
    .Y(net6262));
 BUFx3_ASAP7_75t_R place6263 (.A(_10867_),
    .Y(net6263));
 BUFx6f_ASAP7_75t_R place6264 (.A(_10822_),
    .Y(net6264));
 BUFx6f_ASAP7_75t_R place6265 (.A(_10822_),
    .Y(net6265));
 BUFx6f_ASAP7_75t_R place6266 (.A(_10822_),
    .Y(net6266));
 BUFx3_ASAP7_75t_R place6267 (.A(_10818_),
    .Y(net6267));
 BUFx6f_ASAP7_75t_R place6268 (.A(_10818_),
    .Y(net6268));
 BUFx3_ASAP7_75t_R place6269 (.A(net6271),
    .Y(net6269));
 BUFx3_ASAP7_75t_R place6270 (.A(net6271),
    .Y(net6270));
 BUFx6f_ASAP7_75t_R place6271 (.A(_10784_),
    .Y(net6271));
 BUFx6f_ASAP7_75t_R place6272 (.A(_10784_),
    .Y(net6272));
 BUFx3_ASAP7_75t_R place6273 (.A(_10770_),
    .Y(net6273));
 BUFx6f_ASAP7_75t_R place6274 (.A(_10770_),
    .Y(net6274));
 BUFx6f_ASAP7_75t_R place6275 (.A(net6277),
    .Y(net6275));
 BUFx6f_ASAP7_75t_R place6276 (.A(net6277),
    .Y(net6276));
 BUFx6f_ASAP7_75t_R place6277 (.A(_10770_),
    .Y(net6277));
 BUFx6f_ASAP7_75t_R place6278 (.A(_10752_),
    .Y(net6278));
 BUFx3_ASAP7_75t_R place6279 (.A(_10739_),
    .Y(net6279));
 BUFx3_ASAP7_75t_R place6280 (.A(_10738_),
    .Y(net6280));
 BUFx3_ASAP7_75t_R place6281 (.A(_10735_),
    .Y(net6281));
 BUFx3_ASAP7_75t_R place6282 (.A(_10734_),
    .Y(net6282));
 BUFx3_ASAP7_75t_R place6283 (.A(_10731_),
    .Y(net6283));
 BUFx3_ASAP7_75t_R place6284 (.A(_10730_),
    .Y(net6284));
 BUFx3_ASAP7_75t_R place6285 (.A(_10694_),
    .Y(net6285));
 BUFx3_ASAP7_75t_R place6286 (.A(_10686_),
    .Y(net6286));
 BUFx3_ASAP7_75t_R place6287 (.A(_10111_),
    .Y(net6287));
 BUFx3_ASAP7_75t_R place6288 (.A(net6289),
    .Y(net6288));
 BUFx6f_ASAP7_75t_R place6289 (.A(_10106_),
    .Y(net6289));
 BUFx3_ASAP7_75t_R place6290 (.A(_10106_),
    .Y(net6290));
 BUFx3_ASAP7_75t_R place6291 (.A(_10106_),
    .Y(net6291));
 BUFx6f_ASAP7_75t_R place6292 (.A(_10106_),
    .Y(net6292));
 BUFx3_ASAP7_75t_R place6293 (.A(_09591_),
    .Y(net6293));
 BUFx3_ASAP7_75t_R place6294 (.A(net6295),
    .Y(net6294));
 BUFx6f_ASAP7_75t_R place6295 (.A(_09591_),
    .Y(net6295));
 BUFx3_ASAP7_75t_R place6296 (.A(_09567_),
    .Y(net6296));
 BUFx6f_ASAP7_75t_R place6297 (.A(_09021_),
    .Y(net6297));
 BUFx3_ASAP7_75t_R place6298 (.A(_09006_),
    .Y(net6298));
 BUFx3_ASAP7_75t_R place6299 (.A(net6300),
    .Y(net6299));
 BUFx3_ASAP7_75t_R place6300 (.A(_08997_),
    .Y(net6300));
 BUFx3_ASAP7_75t_R place6301 (.A(_08992_),
    .Y(net6301));
 BUFx3_ASAP7_75t_R place6302 (.A(_08992_),
    .Y(net6302));
 BUFx6f_ASAP7_75t_R place6303 (.A(_08976_),
    .Y(net6303));
 BUFx6f_ASAP7_75t_R place6304 (.A(_08972_),
    .Y(net6304));
 BUFx6f_ASAP7_75t_R place6305 (.A(net6307),
    .Y(net6305));
 BUFx6f_ASAP7_75t_R place6306 (.A(net6307),
    .Y(net6306));
 BUFx6f_ASAP7_75t_R place6307 (.A(_08967_),
    .Y(net6307));
 BUFx3_ASAP7_75t_R place6308 (.A(_08961_),
    .Y(net6308));
 BUFx3_ASAP7_75t_R place6309 (.A(_08955_),
    .Y(net6309));
 BUFx3_ASAP7_75t_R place6310 (.A(net6311),
    .Y(net6310));
 BUFx3_ASAP7_75t_R place6311 (.A(_08950_),
    .Y(net6311));
 BUFx3_ASAP7_75t_R place6312 (.A(_08936_),
    .Y(net6312));
 BUFx3_ASAP7_75t_R place6313 (.A(_08936_),
    .Y(net6313));
 BUFx3_ASAP7_75t_R place6314 (.A(net6318),
    .Y(net6314));
 BUFx3_ASAP7_75t_R place6315 (.A(net6318),
    .Y(net6315));
 BUFx3_ASAP7_75t_R place6316 (.A(net6318),
    .Y(net6316));
 BUFx6f_ASAP7_75t_R place6317 (.A(net6318),
    .Y(net6317));
 BUFx6f_ASAP7_75t_R place6318 (.A(_08933_),
    .Y(net6318));
 BUFx3_ASAP7_75t_R place6319 (.A(net6320),
    .Y(net6319));
 BUFx6f_ASAP7_75t_R place6320 (.A(_08928_),
    .Y(net6320));
 BUFx3_ASAP7_75t_R place6321 (.A(_08922_),
    .Y(net6321));
 BUFx3_ASAP7_75t_R place6322 (.A(_08922_),
    .Y(net6322));
 BUFx3_ASAP7_75t_R place6323 (.A(_08916_),
    .Y(net6323));
 BUFx3_ASAP7_75t_R place6324 (.A(_08911_),
    .Y(net6324));
 BUFx3_ASAP7_75t_R place6325 (.A(_08911_),
    .Y(net6325));
 BUFx6f_ASAP7_75t_R place6326 (.A(_08111_),
    .Y(net6326));
 BUFx6f_ASAP7_75t_R place6327 (.A(_08111_),
    .Y(net6327));
 BUFx3_ASAP7_75t_R place6328 (.A(net6330),
    .Y(net6328));
 BUFx3_ASAP7_75t_R place6329 (.A(net6330),
    .Y(net6329));
 BUFx6f_ASAP7_75t_R place6330 (.A(_08111_),
    .Y(net6330));
 BUFx3_ASAP7_75t_R place6331 (.A(_08102_),
    .Y(net6331));
 BUFx3_ASAP7_75t_R place6332 (.A(_08090_),
    .Y(net6332));
 BUFx6f_ASAP7_75t_R place6333 (.A(_08082_),
    .Y(net6333));
 BUFx6f_ASAP7_75t_R place6334 (.A(net6336),
    .Y(net6334));
 BUFx3_ASAP7_75t_R place6335 (.A(net6336),
    .Y(net6335));
 BUFx6f_ASAP7_75t_R place6336 (.A(_08074_),
    .Y(net6336));
 BUFx3_ASAP7_75t_R place6337 (.A(_00980_),
    .Y(net6337));
 BUFx3_ASAP7_75t_R place6338 (.A(_08060_),
    .Y(net6338));
 BUFx3_ASAP7_75t_R place6339 (.A(_08060_),
    .Y(net6339));
 BUFx6f_ASAP7_75t_R place6340 (.A(_08051_),
    .Y(net6340));
 BUFx3_ASAP7_75t_R place6341 (.A(_07121_),
    .Y(net6341));
 BUFx3_ASAP7_75t_R place6342 (.A(_07116_),
    .Y(net6342));
 BUFx3_ASAP7_75t_R place6343 (.A(_06454_),
    .Y(net6343));
 BUFx3_ASAP7_75t_R place6344 (.A(_05763_),
    .Y(net6344));
 BUFx3_ASAP7_75t_R place6345 (.A(_05757_),
    .Y(net6345));
 BUFx3_ASAP7_75t_R place6346 (.A(_04403_),
    .Y(net6346));
 BUFx3_ASAP7_75t_R place6347 (.A(_04392_),
    .Y(net6347));
 BUFx3_ASAP7_75t_R place6348 (.A(_04387_),
    .Y(net6348));
 BUFx3_ASAP7_75t_R place6349 (.A(_03677_),
    .Y(net6349));
 BUFx3_ASAP7_75t_R place6350 (.A(_03672_),
    .Y(net6350));
 BUFx3_ASAP7_75t_R place6351 (.A(_03005_),
    .Y(net6351));
 BUFx3_ASAP7_75t_R place6352 (.A(_02294_),
    .Y(net6352));
 BUFx3_ASAP7_75t_R place6353 (.A(_01597_),
    .Y(net6353));
 BUFx3_ASAP7_75t_R place6354 (.A(_01592_),
    .Y(net6354));
 BUFx3_ASAP7_75t_R place6355 (.A(_14940_),
    .Y(net6355));
 BUFx3_ASAP7_75t_R place6356 (.A(_14926_),
    .Y(net6356));
 BUFx3_ASAP7_75t_R place6357 (.A(_14251_),
    .Y(net6357));
 BUFx3_ASAP7_75t_R place6358 (.A(_14237_),
    .Y(net6358));
 BUFx3_ASAP7_75t_R place6359 (.A(_13532_),
    .Y(net6359));
 BUFx3_ASAP7_75t_R place6360 (.A(_12844_),
    .Y(net6360));
 BUFx3_ASAP7_75t_R place6361 (.A(_12152_),
    .Y(net6361));
 BUFx3_ASAP7_75t_R place6362 (.A(_11406_),
    .Y(net6362));
 BUFx3_ASAP7_75t_R place6363 (.A(_11402_),
    .Y(net6363));
 BUFx3_ASAP7_75t_R place6364 (.A(_10707_),
    .Y(net6364));
 BUFx3_ASAP7_75t_R place6365 (.A(_10692_),
    .Y(net6365));
 BUFx3_ASAP7_75t_R place6366 (.A(_10685_),
    .Y(net6366));
 BUFx3_ASAP7_75t_R place6367 (.A(_08960_),
    .Y(net6367));
 BUFx3_ASAP7_75t_R place6368 (.A(_08921_),
    .Y(net6368));
 BUFx3_ASAP7_75t_R place6369 (.A(_08058_),
    .Y(net6369));
 BUFx3_ASAP7_75t_R place6370 (.A(net6372),
    .Y(net6370));
 BUFx6f_ASAP7_75t_R place6371 (.A(net6372),
    .Y(net6371));
 BUFx6f_ASAP7_75t_R place6372 (.A(_08058_),
    .Y(net6372));
 BUFx6f_ASAP7_75t_R place6373 (.A(_08058_),
    .Y(net6373));
 BUFx3_ASAP7_75t_R place6374 (.A(net6378),
    .Y(net6374));
 BUFx3_ASAP7_75t_R place6375 (.A(net6378),
    .Y(net6375));
 BUFx3_ASAP7_75t_R place6376 (.A(net6378),
    .Y(net6376));
 BUFx3_ASAP7_75t_R place6377 (.A(net6378),
    .Y(net6377));
 BUFx6f_ASAP7_75t_R place6378 (.A(_08043_),
    .Y(net6378));
 BUFx6f_ASAP7_75t_R place6379 (.A(net6380),
    .Y(net6379));
 BUFx3_ASAP7_75t_R place6380 (.A(_08043_),
    .Y(net6380));
 BUFx3_ASAP7_75t_R place6381 (.A(_05762_),
    .Y(net6381));
 BUFx3_ASAP7_75t_R place6382 (.A(_05090_),
    .Y(net6382));
 BUFx3_ASAP7_75t_R place6383 (.A(_08787_),
    .Y(net6383));
 BUFx3_ASAP7_75t_R place6384 (.A(_05772_),
    .Y(net6384));
 BUFx3_ASAP7_75t_R place6385 (.A(_05771_),
    .Y(net6385));
 BUFx3_ASAP7_75t_R place6386 (.A(_03693_),
    .Y(net6386));
 BUFx3_ASAP7_75t_R place6387 (.A(_14239_),
    .Y(net6387));
 BUFx3_ASAP7_75t_R place6388 (.A(_08999_),
    .Y(net6388));
 BUFx3_ASAP7_75t_R place6389 (.A(_08817_),
    .Y(net6389));
 BUFx3_ASAP7_75t_R place6390 (.A(_08793_),
    .Y(net6390));
 BUFx3_ASAP7_75t_R place6391 (.A(_06458_),
    .Y(net6391));
 BUFx3_ASAP7_75t_R place6392 (.A(_06442_),
    .Y(net6392));
 BUFx3_ASAP7_75t_R place6393 (.A(_05752_),
    .Y(net6393));
 BUFx3_ASAP7_75t_R place6394 (.A(_05115_),
    .Y(net6394));
 BUFx3_ASAP7_75t_R place6395 (.A(_04410_),
    .Y(net6395));
 BUFx3_ASAP7_75t_R place6396 (.A(_04396_),
    .Y(net6396));
 BUFx3_ASAP7_75t_R place6397 (.A(_04395_),
    .Y(net6397));
 BUFx3_ASAP7_75t_R place6398 (.A(_03680_),
    .Y(net6398));
 BUFx3_ASAP7_75t_R place6399 (.A(_02996_),
    .Y(net6399));
 BUFx3_ASAP7_75t_R place6400 (.A(_02982_),
    .Y(net6400));
 BUFx3_ASAP7_75t_R place6401 (.A(_02981_),
    .Y(net6401));
 BUFx3_ASAP7_75t_R place6402 (.A(_02282_),
    .Y(net6402));
 BUFx3_ASAP7_75t_R place6403 (.A(_01773_),
    .Y(net6403));
 BUFx3_ASAP7_75t_R place6404 (.A(_01589_),
    .Y(net6404));
 BUFx3_ASAP7_75t_R place6405 (.A(_01585_),
    .Y(net6405));
 BUFx3_ASAP7_75t_R place6406 (.A(_01584_),
    .Y(net6406));
 BUFx3_ASAP7_75t_R place6407 (.A(_01581_),
    .Y(net6407));
 BUFx3_ASAP7_75t_R place6408 (.A(_14936_),
    .Y(net6408));
 BUFx3_ASAP7_75t_R place6409 (.A(_14928_),
    .Y(net6409));
 BUFx3_ASAP7_75t_R place6410 (.A(_14922_),
    .Y(net6410));
 BUFx3_ASAP7_75t_R place6411 (.A(_14918_),
    .Y(net6411));
 BUFx3_ASAP7_75t_R place6412 (.A(_14917_),
    .Y(net6412));
 BUFx3_ASAP7_75t_R place6413 (.A(_14915_),
    .Y(net6413));
 BUFx3_ASAP7_75t_R place6414 (.A(_14218_),
    .Y(net6414));
 BUFx3_ASAP7_75t_R place6415 (.A(_14217_),
    .Y(net6415));
 BUFx3_ASAP7_75t_R place6416 (.A(_13541_),
    .Y(net6416));
 BUFx3_ASAP7_75t_R place6417 (.A(_13528_),
    .Y(net6417));
 BUFx3_ASAP7_75t_R place6418 (.A(_13524_),
    .Y(net6418));
 BUFx3_ASAP7_75t_R place6419 (.A(_13521_),
    .Y(net6419));
 BUFx3_ASAP7_75t_R place6420 (.A(_12853_),
    .Y(net6420));
 BUFx3_ASAP7_75t_R place6421 (.A(_12851_),
    .Y(net6421));
 BUFx3_ASAP7_75t_R place6422 (.A(_12846_),
    .Y(net6422));
 BUFx3_ASAP7_75t_R place6423 (.A(_12838_),
    .Y(net6423));
 BUFx3_ASAP7_75t_R place6424 (.A(_12834_),
    .Y(net6424));
 BUFx3_ASAP7_75t_R place6425 (.A(_12818_),
    .Y(net6425));
 BUFx3_ASAP7_75t_R place6426 (.A(_12815_),
    .Y(net6426));
 BUFx3_ASAP7_75t_R place6427 (.A(_12319_),
    .Y(net6427));
 BUFx3_ASAP7_75t_R place6428 (.A(_12192_),
    .Y(net6428));
 BUFx3_ASAP7_75t_R place6429 (.A(net6430),
    .Y(net6429));
 BUFx3_ASAP7_75t_R place6430 (.A(_12162_),
    .Y(net6430));
 BUFx3_ASAP7_75t_R place6431 (.A(_12160_),
    .Y(net6431));
 BUFx3_ASAP7_75t_R place6432 (.A(_12154_),
    .Y(net6432));
 BUFx3_ASAP7_75t_R place6433 (.A(_12141_),
    .Y(net6433));
 BUFx3_ASAP7_75t_R place6434 (.A(_12140_),
    .Y(net6434));
 BUFx3_ASAP7_75t_R place6435 (.A(_12129_),
    .Y(net6435));
 BUFx6f_ASAP7_75t_R place6436 (.A(_12127_),
    .Y(net6436));
 BUFx3_ASAP7_75t_R place6437 (.A(_12124_),
    .Y(net6437));
 BUFx3_ASAP7_75t_R place6438 (.A(_12123_),
    .Y(net6438));
 BUFx3_ASAP7_75t_R place6439 (.A(_12121_),
    .Y(net6439));
 BUFx3_ASAP7_75t_R place6440 (.A(_11565_),
    .Y(net6440));
 BUFx3_ASAP7_75t_R place6441 (.A(_11428_),
    .Y(net6441));
 BUFx3_ASAP7_75t_R place6442 (.A(_11415_),
    .Y(net6442));
 BUFx3_ASAP7_75t_R place6443 (.A(_11397_),
    .Y(net6443));
 BUFx3_ASAP7_75t_R place6444 (.A(_11396_),
    .Y(net6444));
 BUFx3_ASAP7_75t_R place6445 (.A(_10858_),
    .Y(net6445));
 BUFx3_ASAP7_75t_R place6446 (.A(_10719_),
    .Y(net6446));
 BUFx3_ASAP7_75t_R place6447 (.A(_10717_),
    .Y(net6447));
 BUFx3_ASAP7_75t_R place6448 (.A(_10701_),
    .Y(net6448));
 BUFx3_ASAP7_75t_R place6449 (.A(_10696_),
    .Y(net6449));
 BUFx3_ASAP7_75t_R place6450 (.A(_10682_),
    .Y(net6450));
 BUFx3_ASAP7_75t_R place6451 (.A(_10680_),
    .Y(net6451));
 BUFx3_ASAP7_75t_R place6452 (.A(net6453),
    .Y(net6452));
 BUFx6f_ASAP7_75t_R place6453 (.A(_10679_),
    .Y(net6453));
 BUFx6f_ASAP7_75t_R place6454 (.A(net6455),
    .Y(net6454));
 BUFx3_ASAP7_75t_R place6455 (.A(_10676_),
    .Y(net6455));
 BUFx3_ASAP7_75t_R place6456 (.A(net6460),
    .Y(net6456));
 BUFx3_ASAP7_75t_R place6457 (.A(net6460),
    .Y(net6457));
 BUFx3_ASAP7_75t_R place6458 (.A(net6460),
    .Y(net6458));
 BUFx6f_ASAP7_75t_R place6459 (.A(net6460),
    .Y(net6459));
 BUFx6f_ASAP7_75t_R place6460 (.A(_10676_),
    .Y(net6460));
 BUFx6f_ASAP7_75t_R place6461 (.A(net6464),
    .Y(net6461));
 BUFx6f_ASAP7_75t_R place6462 (.A(net6464),
    .Y(net6462));
 BUFx3_ASAP7_75t_R place6463 (.A(net6464),
    .Y(net6463));
 BUFx3_ASAP7_75t_R place6464 (.A(_10676_),
    .Y(net6464));
 BUFx3_ASAP7_75t_R place6465 (.A(_08956_),
    .Y(net6465));
 BUFx3_ASAP7_75t_R place6466 (.A(_08917_),
    .Y(net6466));
 BUFx3_ASAP7_75t_R place6467 (.A(_08881_),
    .Y(net6467));
 BUFx3_ASAP7_75t_R place6468 (.A(_08841_),
    .Y(net6468));
 BUFx3_ASAP7_75t_R place6469 (.A(_08742_),
    .Y(net6469));
 BUFx3_ASAP7_75t_R place6470 (.A(_08723_),
    .Y(net6470));
 BUFx3_ASAP7_75t_R place6471 (.A(_08720_),
    .Y(net6471));
 BUFx3_ASAP7_75t_R place6472 (.A(_00486_),
    .Y(net6472));
 BUFx3_ASAP7_75t_R place6473 (.A(_00945_),
    .Y(net6473));
 BUFx3_ASAP7_75t_R place6474 (.A(_00942_),
    .Y(net6474));
 BUFx3_ASAP7_75t_R place6475 (.A(_00941_),
    .Y(net6475));
 BUFx3_ASAP7_75t_R place6476 (.A(_00935_),
    .Y(net6476));
 BUFx3_ASAP7_75t_R place6477 (.A(_00934_),
    .Y(net6477));
 BUFx3_ASAP7_75t_R place6478 (.A(_00933_),
    .Y(net6478));
 BUFx3_ASAP7_75t_R place6479 (.A(_00932_),
    .Y(net6479));
 BUFx3_ASAP7_75t_R place6480 (.A(_00924_),
    .Y(net6480));
 BUFx3_ASAP7_75t_R place6481 (.A(_00921_),
    .Y(net6481));
 BUFx3_ASAP7_75t_R place6482 (.A(_00920_),
    .Y(net6482));
 BUFx3_ASAP7_75t_R place6483 (.A(_00919_),
    .Y(net6483));
 BUFx3_ASAP7_75t_R place6484 (.A(_00918_),
    .Y(net6484));
 BUFx3_ASAP7_75t_R place6485 (.A(_00917_),
    .Y(net6485));
 BUFx3_ASAP7_75t_R place6486 (.A(_00914_),
    .Y(net6486));
 BUFx3_ASAP7_75t_R place6487 (.A(_00913_),
    .Y(net6487));
 BUFx3_ASAP7_75t_R place6488 (.A(_00910_),
    .Y(net6488));
 BUFx3_ASAP7_75t_R place6489 (.A(_00909_),
    .Y(net6489));
 BUFx3_ASAP7_75t_R place6490 (.A(_00904_),
    .Y(net6490));
 BUFx3_ASAP7_75t_R place6491 (.A(_00903_),
    .Y(net6491));
 BUFx3_ASAP7_75t_R place6492 (.A(_00902_),
    .Y(net6492));
 BUFx3_ASAP7_75t_R place6493 (.A(_00901_),
    .Y(net6493));
 BUFx3_ASAP7_75t_R place6494 (.A(_00900_),
    .Y(net6494));
 BUFx3_ASAP7_75t_R place6495 (.A(_00898_),
    .Y(net6495));
 BUFx3_ASAP7_75t_R place6496 (.A(_00897_),
    .Y(net6496));
 BUFx3_ASAP7_75t_R place6497 (.A(_00896_),
    .Y(net6497));
 BUFx3_ASAP7_75t_R place6498 (.A(_00895_),
    .Y(net6498));
 BUFx3_ASAP7_75t_R place6499 (.A(_00892_),
    .Y(net6499));
 BUFx3_ASAP7_75t_R place6500 (.A(_00889_),
    .Y(net6500));
 BUFx3_ASAP7_75t_R place6501 (.A(_00888_),
    .Y(net6501));
 BUFx3_ASAP7_75t_R place6502 (.A(_00887_),
    .Y(net6502));
 BUFx3_ASAP7_75t_R place6503 (.A(_00886_),
    .Y(net6503));
 BUFx3_ASAP7_75t_R place6504 (.A(_00885_),
    .Y(net6504));
 BUFx3_ASAP7_75t_R place6505 (.A(_00881_),
    .Y(net6505));
 BUFx3_ASAP7_75t_R place6506 (.A(_00879_),
    .Y(net6506));
 BUFx3_ASAP7_75t_R place6507 (.A(_00878_),
    .Y(net6507));
 BUFx3_ASAP7_75t_R place6508 (.A(_00877_),
    .Y(net6508));
 BUFx3_ASAP7_75t_R place6509 (.A(_00873_),
    .Y(net6509));
 BUFx3_ASAP7_75t_R place6510 (.A(_00872_),
    .Y(net6510));
 BUFx3_ASAP7_75t_R place6511 (.A(_00871_),
    .Y(net6511));
 BUFx3_ASAP7_75t_R place6512 (.A(_00870_),
    .Y(net6512));
 BUFx3_ASAP7_75t_R place6513 (.A(_00869_),
    .Y(net6513));
 BUFx3_ASAP7_75t_R place6514 (.A(_00868_),
    .Y(net6514));
 BUFx3_ASAP7_75t_R place6515 (.A(_00867_),
    .Y(net6515));
 BUFx3_ASAP7_75t_R place6516 (.A(_00866_),
    .Y(net6516));
 BUFx3_ASAP7_75t_R place6517 (.A(_00865_),
    .Y(net6517));
 BUFx3_ASAP7_75t_R place6518 (.A(_00864_),
    .Y(net6518));
 BUFx3_ASAP7_75t_R place6519 (.A(_00863_),
    .Y(net6519));
 BUFx3_ASAP7_75t_R place6520 (.A(_00862_),
    .Y(net6520));
 BUFx3_ASAP7_75t_R place6521 (.A(_00861_),
    .Y(net6521));
 BUFx3_ASAP7_75t_R place6522 (.A(_00860_),
    .Y(net6522));
 BUFx3_ASAP7_75t_R place6523 (.A(_00859_),
    .Y(net6523));
 BUFx3_ASAP7_75t_R place6524 (.A(_00858_),
    .Y(net6524));
 BUFx3_ASAP7_75t_R place6525 (.A(_00857_),
    .Y(net6525));
 BUFx3_ASAP7_75t_R place6526 (.A(_00856_),
    .Y(net6526));
 BUFx3_ASAP7_75t_R place6527 (.A(_00855_),
    .Y(net6527));
 BUFx3_ASAP7_75t_R place6528 (.A(_00854_),
    .Y(net6528));
 BUFx3_ASAP7_75t_R place6529 (.A(_00849_),
    .Y(net6529));
 BUFx3_ASAP7_75t_R place6530 (.A(_00848_),
    .Y(net6530));
 BUFx3_ASAP7_75t_R place6531 (.A(_00847_),
    .Y(net6531));
 BUFx3_ASAP7_75t_R place6532 (.A(_00846_),
    .Y(net6532));
 BUFx3_ASAP7_75t_R place6533 (.A(_00845_),
    .Y(net6533));
 BUFx3_ASAP7_75t_R place6534 (.A(_00843_),
    .Y(net6534));
 BUFx3_ASAP7_75t_R place6535 (.A(_00842_),
    .Y(net6535));
 BUFx3_ASAP7_75t_R place6536 (.A(_00841_),
    .Y(net6536));
 BUFx3_ASAP7_75t_R place6537 (.A(_00840_),
    .Y(net6537));
 BUFx3_ASAP7_75t_R place6538 (.A(_00839_),
    .Y(net6538));
 BUFx3_ASAP7_75t_R place6539 (.A(_00838_),
    .Y(net6539));
 BUFx3_ASAP7_75t_R place6540 (.A(_00421_),
    .Y(net6540));
 BUFx3_ASAP7_75t_R place6541 (.A(_00429_),
    .Y(net6541));
 BUFx3_ASAP7_75t_R place6542 (.A(_00569_),
    .Y(net6542));
 BUFx3_ASAP7_75t_R place6543 (.A(_00699_),
    .Y(net6543));
 BUFx6f_ASAP7_75t_R place6544 (.A(_00697_),
    .Y(net6544));
 BUFx3_ASAP7_75t_R place6545 (.A(net6547),
    .Y(net6545));
 BUFx3_ASAP7_75t_R place6546 (.A(net6547),
    .Y(net6546));
 BUFx6f_ASAP7_75t_R place6547 (.A(_00696_),
    .Y(net6547));
 BUFx3_ASAP7_75t_R place6548 (.A(_00695_),
    .Y(net6548));
 BUFx3_ASAP7_75t_R place6549 (.A(_00694_),
    .Y(net6549));
 BUFx3_ASAP7_75t_R place6550 (.A(_00690_),
    .Y(net6550));
 BUFx3_ASAP7_75t_R place6551 (.A(_00689_),
    .Y(net6551));
 BUFx3_ASAP7_75t_R place6552 (.A(_00688_),
    .Y(net6552));
 BUFx3_ASAP7_75t_R place6553 (.A(_00687_),
    .Y(net6553));
 BUFx3_ASAP7_75t_R place6554 (.A(_00686_),
    .Y(net6554));
 BUFx3_ASAP7_75t_R place6555 (.A(_00684_),
    .Y(net6555));
 BUFx3_ASAP7_75t_R place6556 (.A(_00683_),
    .Y(net6556));
 BUFx3_ASAP7_75t_R place6557 (.A(_00681_),
    .Y(net6557));
 BUFx3_ASAP7_75t_R place6558 (.A(_00680_),
    .Y(net6558));
 BUFx3_ASAP7_75t_R place6559 (.A(_00679_),
    .Y(net6559));
 BUFx3_ASAP7_75t_R place6560 (.A(_00678_),
    .Y(net6560));
 BUFx3_ASAP7_75t_R place6561 (.A(_00676_),
    .Y(net6561));
 BUFx3_ASAP7_75t_R place6562 (.A(_00675_),
    .Y(net6562));
 BUFx3_ASAP7_75t_R place6563 (.A(_00674_),
    .Y(net6563));
 BUFx3_ASAP7_75t_R place6564 (.A(_00673_),
    .Y(net6564));
 BUFx3_ASAP7_75t_R place6565 (.A(_00672_),
    .Y(net6565));
 BUFx3_ASAP7_75t_R place6566 (.A(net6569),
    .Y(net6566));
 BUFx6f_ASAP7_75t_R place6567 (.A(net6569),
    .Y(net6567));
 BUFx3_ASAP7_75t_R place6568 (.A(net6569),
    .Y(net6568));
 BUFx6f_ASAP7_75t_R place6569 (.A(_00671_),
    .Y(net6569));
 BUFx3_ASAP7_75t_R place6570 (.A(net6571),
    .Y(net6570));
 BUFx3_ASAP7_75t_R place6571 (.A(_00670_),
    .Y(net6571));
 BUFx3_ASAP7_75t_R place6572 (.A(_00667_),
    .Y(net6572));
 BUFx3_ASAP7_75t_R place6573 (.A(_00666_),
    .Y(net6573));
 BUFx3_ASAP7_75t_R place6574 (.A(_00665_),
    .Y(net6574));
 BUFx3_ASAP7_75t_R place6575 (.A(_00664_),
    .Y(net6575));
 BUFx3_ASAP7_75t_R place6576 (.A(net6577),
    .Y(net6576));
 BUFx6f_ASAP7_75t_R place6577 (.A(_00663_),
    .Y(net6577));
 BUFx3_ASAP7_75t_R place6578 (.A(_00662_),
    .Y(net6578));
 BUFx3_ASAP7_75t_R place6579 (.A(_00662_),
    .Y(net6579));
 BUFx3_ASAP7_75t_R place6580 (.A(_00662_),
    .Y(net6580));
 BUFx3_ASAP7_75t_R place6581 (.A(_00658_),
    .Y(net6581));
 BUFx3_ASAP7_75t_R place6582 (.A(_00657_),
    .Y(net6582));
 BUFx3_ASAP7_75t_R place6583 (.A(_00657_),
    .Y(net6583));
 BUFx3_ASAP7_75t_R place6584 (.A(_00656_),
    .Y(net6584));
 BUFx3_ASAP7_75t_R place6585 (.A(_00655_),
    .Y(net6585));
 BUFx3_ASAP7_75t_R place6586 (.A(_00655_),
    .Y(net6586));
 BUFx3_ASAP7_75t_R place6587 (.A(_00654_),
    .Y(net6587));
 BUFx3_ASAP7_75t_R place6588 (.A(_00652_),
    .Y(net6588));
 BUFx3_ASAP7_75t_R place6589 (.A(_00649_),
    .Y(net6589));
 BUFx3_ASAP7_75t_R place6590 (.A(net6591),
    .Y(net6590));
 BUFx6f_ASAP7_75t_R place6591 (.A(_00648_),
    .Y(net6591));
 BUFx3_ASAP7_75t_R place6592 (.A(_00646_),
    .Y(net6592));
 BUFx3_ASAP7_75t_R place6593 (.A(_00646_),
    .Y(net6593));
 BUFx3_ASAP7_75t_R place6594 (.A(_00644_),
    .Y(net6594));
 BUFx3_ASAP7_75t_R place6595 (.A(_00642_),
    .Y(net6595));
 BUFx3_ASAP7_75t_R place6596 (.A(_00641_),
    .Y(net6596));
 BUFx3_ASAP7_75t_R place6597 (.A(_00640_),
    .Y(net6597));
 BUFx3_ASAP7_75t_R place6598 (.A(_00639_),
    .Y(net6598));
 BUFx3_ASAP7_75t_R place6599 (.A(_00639_),
    .Y(net6599));
 BUFx3_ASAP7_75t_R place6600 (.A(net6601),
    .Y(net6600));
 BUFx3_ASAP7_75t_R place6601 (.A(_00638_),
    .Y(net6601));
 BUFx3_ASAP7_75t_R place6602 (.A(_00633_),
    .Y(net6602));
 BUFx3_ASAP7_75t_R place6603 (.A(_00631_),
    .Y(net6603));
 BUFx3_ASAP7_75t_R place6604 (.A(net6606),
    .Y(net6604));
 BUFx3_ASAP7_75t_R place6605 (.A(net6606),
    .Y(net6605));
 BUFx3_ASAP7_75t_R place6606 (.A(_00630_),
    .Y(net6606));
 BUFx3_ASAP7_75t_R place6607 (.A(_00629_),
    .Y(net6607));
 BUFx3_ASAP7_75t_R place6608 (.A(_00627_),
    .Y(net6608));
 BUFx3_ASAP7_75t_R place6609 (.A(_00626_),
    .Y(net6609));
 BUFx6f_ASAP7_75t_R place6610 (.A(_00625_),
    .Y(net6610));
 BUFx6f_ASAP7_75t_R place6611 (.A(_00624_),
    .Y(net6611));
 BUFx6f_ASAP7_75t_R place6612 (.A(net6613),
    .Y(net6612));
 BUFx6f_ASAP7_75t_R place6613 (.A(_00623_),
    .Y(net6613));
 BUFx6f_ASAP7_75t_R place6614 (.A(_00622_),
    .Y(net6614));
 BUFx3_ASAP7_75t_R place6615 (.A(_00616_),
    .Y(net6615));
 BUFx3_ASAP7_75t_R place6616 (.A(_00615_),
    .Y(net6616));
 BUFx3_ASAP7_75t_R place6617 (.A(net6618),
    .Y(net6617));
 BUFx6f_ASAP7_75t_R place6618 (.A(_00614_),
    .Y(net6618));
 BUFx3_ASAP7_75t_R place6619 (.A(_00610_),
    .Y(net6619));
 BUFx3_ASAP7_75t_R place6620 (.A(_00609_),
    .Y(net6620));
 BUFx6f_ASAP7_75t_R place6621 (.A(_00608_),
    .Y(net6621));
 BUFx3_ASAP7_75t_R place6622 (.A(net6623),
    .Y(net6622));
 BUFx6f_ASAP7_75t_R place6623 (.A(_00607_),
    .Y(net6623));
 BUFx3_ASAP7_75t_R place6624 (.A(_00606_),
    .Y(net6624));
 BUFx3_ASAP7_75t_R place6625 (.A(_00601_),
    .Y(net6625));
 BUFx3_ASAP7_75t_R place6626 (.A(_00600_),
    .Y(net6626));
 BUFx3_ASAP7_75t_R place6627 (.A(_00600_),
    .Y(net6627));
 BUFx3_ASAP7_75t_R place6628 (.A(_00599_),
    .Y(net6628));
 BUFx3_ASAP7_75t_R place6629 (.A(_00598_),
    .Y(net6629));
 BUFx3_ASAP7_75t_R place6630 (.A(net6631),
    .Y(net6630));
 BUFx6f_ASAP7_75t_R place6631 (.A(_00598_),
    .Y(net6631));
 BUFx3_ASAP7_75t_R place6632 (.A(_00596_),
    .Y(net6632));
 BUFx3_ASAP7_75t_R place6633 (.A(_00594_),
    .Y(net6633));
 BUFx3_ASAP7_75t_R place6634 (.A(_00593_),
    .Y(net6634));
 BUFx3_ASAP7_75t_R place6635 (.A(_00592_),
    .Y(net6635));
 BUFx3_ASAP7_75t_R place6636 (.A(_00592_),
    .Y(net6636));
 BUFx3_ASAP7_75t_R place6637 (.A(_00591_),
    .Y(net6637));
 BUFx3_ASAP7_75t_R place6638 (.A(net6639),
    .Y(net6638));
 BUFx6f_ASAP7_75t_R place6639 (.A(_00591_),
    .Y(net6639));
 BUFx3_ASAP7_75t_R place6640 (.A(_00590_),
    .Y(net6640));
 BUFx3_ASAP7_75t_R place6641 (.A(_00584_),
    .Y(net6641));
 BUFx3_ASAP7_75t_R place6642 (.A(_00583_),
    .Y(net6642));
 BUFx3_ASAP7_75t_R place6643 (.A(_00582_),
    .Y(net6643));
 BUFx6f_ASAP7_75t_R place6644 (.A(_00582_),
    .Y(net6644));
 BUFx3_ASAP7_75t_R place6645 (.A(_00578_),
    .Y(net6645));
 BUFx3_ASAP7_75t_R place6646 (.A(_00577_),
    .Y(net6646));
 BUFx3_ASAP7_75t_R place6647 (.A(net6649),
    .Y(net6647));
 BUFx3_ASAP7_75t_R place6648 (.A(net6649),
    .Y(net6648));
 BUFx6f_ASAP7_75t_R place6649 (.A(_00576_),
    .Y(net6649));
 BUFx3_ASAP7_75t_R place6650 (.A(net6651),
    .Y(net6650));
 BUFx3_ASAP7_75t_R place6651 (.A(_00575_),
    .Y(net6651));
 BUFx3_ASAP7_75t_R place6652 (.A(_00575_),
    .Y(net6652));
 BUFx3_ASAP7_75t_R place6653 (.A(net6664),
    .Y(net6653));
 BUFx3_ASAP7_75t_R place6654 (.A(net6657),
    .Y(net6654));
 BUFx3_ASAP7_75t_R place6655 (.A(net6657),
    .Y(net6655));
 BUFx3_ASAP7_75t_R place6656 (.A(net6657),
    .Y(net6656));
 BUFx6f_ASAP7_75t_R place6657 (.A(net6664),
    .Y(net6657));
 BUFx3_ASAP7_75t_R place6658 (.A(net6660),
    .Y(net6658));
 BUFx3_ASAP7_75t_R place6659 (.A(net6660),
    .Y(net6659));
 BUFx6f_ASAP7_75t_R place6660 (.A(net6664),
    .Y(net6660));
 BUFx3_ASAP7_75t_R place6661 (.A(net6664),
    .Y(net6661));
 BUFx3_ASAP7_75t_R place6662 (.A(net6663),
    .Y(net6662));
 BUFx6f_ASAP7_75t_R place6663 (.A(net6664),
    .Y(net6663));
 BUFx6f_ASAP7_75t_R place6664 (.A(_00574_),
    .Y(net6664));
 BUFx3_ASAP7_75t_R place6665 (.A(net6668),
    .Y(net6665));
 BUFx6f_ASAP7_75t_R place6666 (.A(net6668),
    .Y(net6666));
 BUFx3_ASAP7_75t_R place6667 (.A(net6668),
    .Y(net6667));
 BUFx6f_ASAP7_75t_R place6668 (.A(net6673),
    .Y(net6668));
 BUFx6f_ASAP7_75t_R place6669 (.A(net6673),
    .Y(net6669));
 BUFx3_ASAP7_75t_R place6670 (.A(net6673),
    .Y(net6670));
 BUFx6f_ASAP7_75t_R place6671 (.A(net6673),
    .Y(net6671));
 BUFx3_ASAP7_75t_R place6672 (.A(net6673),
    .Y(net6672));
 BUFx6f_ASAP7_75t_R place6673 (.A(_00574_),
    .Y(net6673));
 BUFx3_ASAP7_75t_R place6674 (.A(_08030_),
    .Y(net6674));
 BUFx3_ASAP7_75t_R place6675 (.A(_08030_),
    .Y(net6675));
 BUFx3_ASAP7_75t_R place6676 (.A(_08030_),
    .Y(net6676));
 BUFx3_ASAP7_75t_R place6677 (.A(_08030_),
    .Y(net6677));
 BUFx3_ASAP7_75t_R place6678 (.A(net6679),
    .Y(net6678));
 BUFx3_ASAP7_75t_R place6679 (.A(_08030_),
    .Y(net6679));
 BUFx6f_ASAP7_75t_R place6680 (.A(net6683),
    .Y(net6680));
 BUFx6f_ASAP7_75t_R place6681 (.A(net6682),
    .Y(net6681));
 BUFx3_ASAP7_75t_R place6682 (.A(net6683),
    .Y(net6682));
 BUFx6f_ASAP7_75t_R place6683 (.A(net129),
    .Y(net6683));
 BUFx3_ASAP7_75t_R place6684 (.A(net129),
    .Y(net6684));
 BUFx3_ASAP7_75t_R place6685 (.A(net129),
    .Y(net6685));
 BUFx3_ASAP7_75t_R place6686 (.A(net6690),
    .Y(net6686));
 BUFx3_ASAP7_75t_R place6687 (.A(net6690),
    .Y(net6687));
 BUFx3_ASAP7_75t_R place6688 (.A(net6689),
    .Y(net6688));
 BUFx6f_ASAP7_75t_R place6689 (.A(net6690),
    .Y(net6689));
 BUFx6f_ASAP7_75t_R place6690 (.A(net129),
    .Y(net6690));
 DFFHQNx1_ASAP7_75t_R \sa00_sr[0]$_DFF_P_  (.CLK(clknet_leaf_16_clk),
    .D(_00032_),
    .QN(_00575_));
 DFFHQNx1_ASAP7_75t_R \sa00_sr[1]$_DFF_P_  (.CLK(clknet_leaf_17_clk),
    .D(_00033_),
    .QN(_00576_));
 DFFHQNx1_ASAP7_75t_R \sa00_sr[2]$_DFF_P_  (.CLK(clknet_leaf_23_clk),
    .D(_00034_),
    .QN(_00577_));
 DFFHQNx1_ASAP7_75t_R \sa00_sr[3]$_DFF_P_  (.CLK(clknet_leaf_22_clk),
    .D(_00035_),
    .QN(_00578_));
 DFFHQNx1_ASAP7_75t_R \sa00_sr[4]$_DFF_P_  (.CLK(clknet_leaf_22_clk),
    .D(_00036_),
    .QN(_00579_));
 DFFHQNx1_ASAP7_75t_R \sa00_sr[5]$_DFF_P_  (.CLK(clknet_leaf_17_clk),
    .D(_00037_),
    .QN(_00580_));
 DFFHQNx1_ASAP7_75t_R \sa00_sr[6]$_DFF_P_  (.CLK(clknet_leaf_22_clk),
    .D(_00038_),
    .QN(_00581_));
 DFFHQNx1_ASAP7_75t_R \sa00_sr[7]$_DFF_P_  (.CLK(clknet_leaf_22_clk),
    .D(_00039_),
    .QN(_00582_));
 DFFHQNx1_ASAP7_75t_R \sa01_sr[0]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .D(_00040_),
    .QN(_00583_));
 DFFHQNx1_ASAP7_75t_R \sa01_sr[1]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .D(_00041_),
    .QN(_00584_));
 DFFHQNx1_ASAP7_75t_R \sa01_sr[2]$_DFF_P_  (.CLK(clknet_leaf_24_clk),
    .D(_00042_),
    .QN(_00585_));
 DFFHQNx1_ASAP7_75t_R \sa01_sr[3]$_DFF_P_  (.CLK(clknet_leaf_25_clk),
    .D(_00043_),
    .QN(_00586_));
 DFFHQNx1_ASAP7_75t_R \sa01_sr[4]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .D(_00044_),
    .QN(_00587_));
 DFFHQNx1_ASAP7_75t_R \sa01_sr[5]$_DFF_P_  (.CLK(clknet_leaf_25_clk),
    .D(_00045_),
    .QN(_00588_));
 DFFHQNx1_ASAP7_75t_R \sa01_sr[6]$_DFF_P_  (.CLK(clknet_leaf_24_clk),
    .D(_00046_),
    .QN(_00589_));
 DFFHQNx1_ASAP7_75t_R \sa01_sr[7]$_DFF_P_  (.CLK(clknet_leaf_24_clk),
    .D(_00047_),
    .QN(_00590_));
 DFFHQNx1_ASAP7_75t_R \sa02_sr[0]$_DFF_P_  (.CLK(clknet_leaf_10_clk),
    .D(_00048_),
    .QN(_00591_));
 DFFHQNx1_ASAP7_75t_R \sa02_sr[1]$_DFF_P_  (.CLK(clknet_leaf_8_clk),
    .D(_00049_),
    .QN(_00592_));
 DFFHQNx1_ASAP7_75t_R \sa02_sr[2]$_DFF_P_  (.CLK(clknet_leaf_9_clk),
    .D(_00050_),
    .QN(_00593_));
 DFFHQNx1_ASAP7_75t_R \sa02_sr[3]$_DFF_P_  (.CLK(clknet_leaf_9_clk),
    .D(_00051_),
    .QN(_00594_));
 DFFHQNx1_ASAP7_75t_R \sa02_sr[4]$_DFF_P_  (.CLK(clknet_leaf_9_clk),
    .D(_00052_),
    .QN(_00595_));
 DFFHQNx1_ASAP7_75t_R \sa02_sr[5]$_DFF_P_  (.CLK(clknet_leaf_9_clk),
    .D(_00053_),
    .QN(_00596_));
 DFFHQNx1_ASAP7_75t_R \sa02_sr[6]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .D(_00054_),
    .QN(_00597_));
 DFFHQNx1_ASAP7_75t_R \sa02_sr[7]$_DFF_P_  (.CLK(clknet_leaf_8_clk),
    .D(_00055_),
    .QN(_00598_));
 DFFHQNx1_ASAP7_75t_R \sa03_sr[0]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .D(_00056_),
    .QN(_00599_));
 DFFHQNx1_ASAP7_75t_R \sa03_sr[1]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .D(_00057_),
    .QN(_00600_));
 DFFHQNx1_ASAP7_75t_R \sa03_sr[2]$_DFF_P_  (.CLK(clknet_leaf_34_clk),
    .D(_00058_),
    .QN(_00601_));
 DFFHQNx1_ASAP7_75t_R \sa03_sr[3]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .D(_00059_),
    .QN(_00602_));
 DFFHQNx1_ASAP7_75t_R \sa03_sr[4]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .D(_00060_),
    .QN(_00603_));
 DFFHQNx1_ASAP7_75t_R \sa03_sr[5]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .D(_00061_),
    .QN(_00604_));
 DFFHQNx1_ASAP7_75t_R \sa03_sr[6]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .D(_00062_),
    .QN(_00605_));
 DFFHQNx1_ASAP7_75t_R \sa03_sr[7]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .D(_00063_),
    .QN(_00606_));
 DFFHQNx1_ASAP7_75t_R \sa10_sr[0]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .D(_00072_),
    .QN(_00607_));
 DFFHQNx1_ASAP7_75t_R \sa10_sr[1]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .D(_00073_),
    .QN(_00608_));
 DFFHQNx1_ASAP7_75t_R \sa10_sr[2]$_DFF_P_  (.CLK(clknet_leaf_25_clk),
    .D(_00074_),
    .QN(_00609_));
 DFFHQNx1_ASAP7_75t_R \sa10_sr[3]$_DFF_P_  (.CLK(clknet_leaf_26_clk),
    .D(_00075_),
    .QN(_00610_));
 DFFHQNx1_ASAP7_75t_R \sa10_sr[4]$_DFF_P_  (.CLK(clknet_leaf_26_clk),
    .D(_00076_),
    .QN(_00611_));
 DFFHQNx1_ASAP7_75t_R \sa10_sr[5]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .D(_00077_),
    .QN(_00612_));
 DFFHQNx1_ASAP7_75t_R \sa10_sr[6]$_DFF_P_  (.CLK(clknet_leaf_25_clk),
    .D(_00078_),
    .QN(_00613_));
 DFFHQNx1_ASAP7_75t_R \sa10_sr[7]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .D(_00079_),
    .QN(_00614_));
 DFFHQNx1_ASAP7_75t_R \sa11_sr[0]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .D(_00080_),
    .QN(_00615_));
 DFFHQNx1_ASAP7_75t_R \sa11_sr[1]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .D(_00081_),
    .QN(_00616_));
 DFFHQNx1_ASAP7_75t_R \sa11_sr[2]$_DFF_P_  (.CLK(clknet_leaf_27_clk),
    .D(_00082_),
    .QN(_00617_));
 DFFHQNx1_ASAP7_75t_R \sa11_sr[3]$_DFF_P_  (.CLK(clknet_leaf_27_clk),
    .D(_00083_),
    .QN(_00618_));
 DFFHQNx1_ASAP7_75t_R \sa11_sr[4]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .D(_00084_),
    .QN(_00619_));
 DFFHQNx1_ASAP7_75t_R \sa11_sr[5]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .D(_00085_),
    .QN(_00620_));
 DFFHQNx1_ASAP7_75t_R \sa11_sr[6]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .D(_00086_),
    .QN(_00621_));
 DFFHQNx1_ASAP7_75t_R \sa11_sr[7]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .D(_00087_),
    .QN(_00622_));
 DFFHQNx1_ASAP7_75t_R \sa12_sr[0]$_DFF_P_  (.CLK(clknet_leaf_9_clk),
    .D(_00088_),
    .QN(_00623_));
 DFFHQNx1_ASAP7_75t_R \sa12_sr[1]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .D(_00089_),
    .QN(_00624_));
 DFFHQNx1_ASAP7_75t_R \sa12_sr[2]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .D(_00090_),
    .QN(_00625_));
 DFFHQNx1_ASAP7_75t_R \sa12_sr[3]$_DFF_P_  (.CLK(clknet_leaf_2_clk),
    .D(_00091_),
    .QN(_00626_));
 DFFHQNx1_ASAP7_75t_R \sa12_sr[4]$_DFF_P_  (.CLK(clknet_leaf_30_clk),
    .D(_00092_),
    .QN(_00627_));
 DFFHQNx1_ASAP7_75t_R \sa12_sr[5]$_DFF_P_  (.CLK(clknet_leaf_31_clk),
    .D(_00093_),
    .QN(_00628_));
 DFFHQNx1_ASAP7_75t_R \sa12_sr[6]$_DFF_P_  (.CLK(clknet_leaf_31_clk),
    .D(_00094_),
    .QN(_00629_));
 DFFHQNx1_ASAP7_75t_R \sa12_sr[7]$_DFF_P_  (.CLK(clknet_leaf_10_clk),
    .D(_00095_),
    .QN(_00630_));
 DFFHQNx1_ASAP7_75t_R \sa13_sr[0]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .D(_00064_),
    .QN(_00631_));
 DFFHQNx1_ASAP7_75t_R \sa13_sr[1]$_DFF_P_  (.CLK(clknet_leaf_30_clk),
    .D(_00065_),
    .QN(_00632_));
 DFFHQNx1_ASAP7_75t_R \sa13_sr[2]$_DFF_P_  (.CLK(clknet_leaf_30_clk),
    .D(_00066_),
    .QN(_00633_));
 DFFHQNx1_ASAP7_75t_R \sa13_sr[3]$_DFF_P_  (.CLK(clknet_leaf_30_clk),
    .D(_00067_),
    .QN(_00634_));
 DFFHQNx1_ASAP7_75t_R \sa13_sr[4]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .D(_00068_),
    .QN(_00635_));
 DFFHQNx1_ASAP7_75t_R \sa13_sr[5]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .D(_00069_),
    .QN(_00636_));
 DFFHQNx1_ASAP7_75t_R \sa13_sr[6]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .D(_00070_),
    .QN(_00637_));
 DFFHQNx1_ASAP7_75t_R \sa13_sr[7]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .D(_00071_),
    .QN(_00638_));
 DFFHQNx1_ASAP7_75t_R \sa20_sr[0]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .D(_00112_),
    .QN(_00639_));
 DFFHQNx1_ASAP7_75t_R \sa20_sr[1]$_DFF_P_  (.CLK(clknet_leaf_12_clk),
    .D(_00113_),
    .QN(_00640_));
 DFFHQNx1_ASAP7_75t_R \sa20_sr[2]$_DFF_P_  (.CLK(clknet_leaf_15_clk),
    .D(_00114_),
    .QN(_00641_));
 DFFHQNx1_ASAP7_75t_R \sa20_sr[3]$_DFF_P_  (.CLK(clknet_leaf_12_clk),
    .D(_00115_),
    .QN(_00642_));
 DFFHQNx1_ASAP7_75t_R \sa20_sr[4]$_DFF_P_  (.CLK(clknet_leaf_12_clk),
    .D(_00116_),
    .QN(_00643_));
 DFFHQNx1_ASAP7_75t_R \sa20_sr[5]$_DFF_P_  (.CLK(clknet_leaf_12_clk),
    .D(_00117_),
    .QN(_00644_));
 DFFHQNx1_ASAP7_75t_R \sa20_sr[6]$_DFF_P_  (.CLK(clknet_leaf_15_clk),
    .D(_00118_),
    .QN(_00645_));
 DFFHQNx1_ASAP7_75t_R \sa20_sr[7]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .D(_00119_),
    .QN(_00646_));
 DFFHQNx1_ASAP7_75t_R \sa21_sr[0]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .D(_00120_),
    .QN(_00647_));
 DFFHQNx1_ASAP7_75t_R \sa21_sr[1]$_DFF_P_  (.CLK(clknet_leaf_19_clk),
    .D(_00121_),
    .QN(_00648_));
 DFFHQNx1_ASAP7_75t_R \sa21_sr[2]$_DFF_P_  (.CLK(clknet_leaf_19_clk),
    .D(_00122_),
    .QN(_00649_));
 DFFHQNx1_ASAP7_75t_R \sa21_sr[3]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .D(_00123_),
    .QN(_00650_));
 DFFHQNx1_ASAP7_75t_R \sa21_sr[4]$_DFF_P_  (.CLK(clknet_leaf_19_clk),
    .D(_00124_),
    .QN(_00651_));
 DFFHQNx1_ASAP7_75t_R \sa21_sr[5]$_DFF_P_  (.CLK(clknet_leaf_11_clk),
    .D(_00125_),
    .QN(_00652_));
 DFFHQNx1_ASAP7_75t_R \sa21_sr[6]$_DFF_P_  (.CLK(clknet_leaf_19_clk),
    .D(_00126_),
    .QN(_00653_));
 DFFHQNx1_ASAP7_75t_R \sa21_sr[7]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .D(_00127_),
    .QN(_00654_));
 DFFHQNx1_ASAP7_75t_R \sa22_sr[0]$_DFF_P_  (.CLK(clknet_leaf_12_clk),
    .D(_00096_),
    .QN(_00655_));
 DFFHQNx2_ASAP7_75t_R \sa22_sr[1]$_DFF_P_  (.CLK(clknet_leaf_11_clk),
    .D(_00097_),
    .QN(_00656_));
 DFFHQNx1_ASAP7_75t_R \sa22_sr[2]$_DFF_P_  (.CLK(clknet_leaf_15_clk),
    .D(_00098_),
    .QN(_00657_));
 DFFHQNx1_ASAP7_75t_R \sa22_sr[3]$_DFF_P_  (.CLK(clknet_leaf_15_clk),
    .D(_00099_),
    .QN(_00658_));
 DFFHQNx1_ASAP7_75t_R \sa22_sr[4]$_DFF_P_  (.CLK(clknet_leaf_12_clk),
    .D(_00100_),
    .QN(_00659_));
 DFFHQNx1_ASAP7_75t_R \sa22_sr[5]$_DFF_P_  (.CLK(clknet_leaf_12_clk),
    .D(_00101_),
    .QN(_00660_));
 DFFHQNx1_ASAP7_75t_R \sa22_sr[6]$_DFF_P_  (.CLK(clknet_leaf_12_clk),
    .D(_00102_),
    .QN(_00661_));
 DFFHQNx1_ASAP7_75t_R \sa22_sr[7]$_DFF_P_  (.CLK(clknet_leaf_11_clk),
    .D(_00103_),
    .QN(_00662_));
 DFFHQNx1_ASAP7_75t_R \sa23_sr[0]$_DFF_P_  (.CLK(clknet_leaf_19_clk),
    .D(_00104_),
    .QN(_00663_));
 DFFHQNx2_ASAP7_75t_R \sa23_sr[1]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .D(_00105_),
    .QN(_00664_));
 DFFHQNx1_ASAP7_75t_R \sa23_sr[2]$_DFF_P_  (.CLK(clknet_leaf_19_clk),
    .D(_00106_),
    .QN(_00665_));
 DFFHQNx1_ASAP7_75t_R \sa23_sr[3]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .D(_00107_),
    .QN(_00666_));
 DFFHQNx1_ASAP7_75t_R \sa23_sr[4]$_DFF_P_  (.CLK(clknet_leaf_19_clk),
    .D(_00108_),
    .QN(_00667_));
 DFFHQNx1_ASAP7_75t_R \sa23_sr[5]$_DFF_P_  (.CLK(clknet_leaf_19_clk),
    .D(_00109_),
    .QN(_00668_));
 DFFHQNx1_ASAP7_75t_R \sa23_sr[6]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .D(_00110_),
    .QN(_00669_));
 DFFHQNx1_ASAP7_75t_R \sa23_sr[7]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .D(_00111_),
    .QN(_00670_));
 DFFHQNx1_ASAP7_75t_R \sa30_sr[0]$_DFF_P_  (.CLK(clknet_leaf_11_clk),
    .D(_00152_),
    .QN(_00671_));
 DFFHQNx1_ASAP7_75t_R \sa30_sr[1]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .D(_00153_),
    .QN(_00672_));
 DFFHQNx1_ASAP7_75t_R \sa30_sr[2]$_DFF_P_  (.CLK(clknet_leaf_10_clk),
    .D(_00154_),
    .QN(_00673_));
 DFFHQNx1_ASAP7_75t_R \sa30_sr[3]$_DFF_P_  (.CLK(clknet_leaf_10_clk),
    .D(_00155_),
    .QN(_00674_));
 DFFHQNx1_ASAP7_75t_R \sa30_sr[4]$_DFF_P_  (.CLK(clknet_leaf_11_clk),
    .D(_00156_),
    .QN(_00675_));
 DFFHQNx1_ASAP7_75t_R \sa30_sr[5]$_DFF_P_  (.CLK(clknet_leaf_11_clk),
    .D(_00157_),
    .QN(_00676_));
 DFFHQNx1_ASAP7_75t_R \sa30_sr[6]$_DFF_P_  (.CLK(clknet_leaf_2_clk),
    .D(_00158_),
    .QN(_00677_));
 DFFHQNx1_ASAP7_75t_R \sa30_sr[7]$_DFF_P_  (.CLK(clknet_leaf_10_clk),
    .D(_00159_),
    .QN(_00678_));
 DFFHQNx1_ASAP7_75t_R \sa31_sr[0]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .D(_00128_),
    .QN(_00679_));
 DFFHQNx1_ASAP7_75t_R \sa31_sr[1]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .D(_00129_),
    .QN(_00680_));
 DFFHQNx1_ASAP7_75t_R \sa31_sr[2]$_DFF_P_  (.CLK(clknet_leaf_17_clk),
    .D(_00130_),
    .QN(_00681_));
 DFFHQNx1_ASAP7_75t_R \sa31_sr[3]$_DFF_P_  (.CLK(clknet_leaf_17_clk),
    .D(_00131_),
    .QN(_00682_));
 DFFHQNx1_ASAP7_75t_R \sa31_sr[4]$_DFF_P_  (.CLK(clknet_leaf_17_clk),
    .D(_00132_),
    .QN(_00683_));
 DFFHQNx1_ASAP7_75t_R \sa31_sr[5]$_DFF_P_  (.CLK(clknet_leaf_17_clk),
    .D(_00133_),
    .QN(_00684_));
 DFFHQNx1_ASAP7_75t_R \sa31_sr[6]$_DFF_P_  (.CLK(clknet_leaf_16_clk),
    .D(_00134_),
    .QN(_00685_));
 DFFHQNx1_ASAP7_75t_R \sa31_sr[7]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .D(_00135_),
    .QN(_00686_));
 DFFHQNx1_ASAP7_75t_R \sa32_sr[0]$_DFF_P_  (.CLK(clknet_leaf_12_clk),
    .D(_00136_),
    .QN(_00687_));
 DFFHQNx1_ASAP7_75t_R \sa32_sr[1]$_DFF_P_  (.CLK(clknet_leaf_12_clk),
    .D(_00137_),
    .QN(_00688_));
 DFFHQNx1_ASAP7_75t_R \sa32_sr[2]$_DFF_P_  (.CLK(clknet_leaf_11_clk),
    .D(_00138_),
    .QN(_00689_));
 DFFHQNx1_ASAP7_75t_R \sa32_sr[3]$_DFF_P_  (.CLK(clknet_leaf_11_clk),
    .D(_00139_),
    .QN(_00690_));
 DFFHQNx1_ASAP7_75t_R \sa32_sr[4]$_DFF_P_  (.CLK(clknet_leaf_11_clk),
    .D(_00140_),
    .QN(_00691_));
 DFFHQNx1_ASAP7_75t_R \sa32_sr[5]$_DFF_P_  (.CLK(clknet_leaf_11_clk),
    .D(_00141_),
    .QN(_00692_));
 DFFHQNx1_ASAP7_75t_R \sa32_sr[6]$_DFF_P_  (.CLK(clknet_leaf_11_clk),
    .D(_00142_),
    .QN(_00693_));
 DFFHQNx1_ASAP7_75t_R \sa32_sr[7]$_DFF_P_  (.CLK(clknet_leaf_11_clk),
    .D(_00143_),
    .QN(_00694_));
 DFFHQNx1_ASAP7_75t_R \sa33_sr[0]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .D(_00144_),
    .QN(_00695_));
 DFFHQNx1_ASAP7_75t_R \sa33_sr[1]$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .D(_00145_),
    .QN(_00696_));
 DFFHQNx1_ASAP7_75t_R \sa33_sr[2]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .D(_00146_),
    .QN(_00697_));
 DFFHQNx1_ASAP7_75t_R \sa33_sr[3]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .D(_00147_),
    .QN(_00698_));
 DFFHQNx1_ASAP7_75t_R \sa33_sr[4]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .D(_00148_),
    .QN(_00699_));
 DFFHQNx1_ASAP7_75t_R \sa33_sr[5]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .D(_00149_),
    .QN(_00700_));
 DFFHQNx1_ASAP7_75t_R \sa33_sr[6]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .D(_00150_),
    .QN(_00701_));
 DFFHQNx1_ASAP7_75t_R \sa33_sr[7]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .D(_00151_),
    .QN(_00569_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[0]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .D(_01409_),
    .QN(_00409_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[100]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_01410_),
    .QN(_00568_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[101]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_01411_),
    .QN(_00567_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[102]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_01412_),
    .QN(_00566_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[103]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_01413_),
    .QN(_00565_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[104]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_01414_),
    .QN(_00469_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[105]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .D(_01415_),
    .QN(_00468_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[106]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .D(_01416_),
    .QN(_00470_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[107]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_01417_),
    .QN(_00564_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[108]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_01418_),
    .QN(_00563_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[109]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_01419_),
    .QN(_00562_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[10]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .D(_01420_),
    .QN(_00479_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[110]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_01421_),
    .QN(_00561_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[111]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_01422_),
    .QN(_00560_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[112]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .D(_01423_),
    .QN(_00457_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[113]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .D(_01424_),
    .QN(_00456_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[114]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .D(_01425_),
    .QN(_00458_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[115]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .D(_01426_),
    .QN(_00559_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[116]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .D(_01427_),
    .QN(_00558_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[117]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .D(_01428_),
    .QN(_00557_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[118]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .D(_01429_),
    .QN(_00556_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[119]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .D(_01430_),
    .QN(_00555_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[11]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .D(_01431_),
    .QN(_00554_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[120]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .D(_01432_),
    .QN(_00445_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[121]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .D(_01433_),
    .QN(_00444_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[122]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .D(_01434_),
    .QN(_00446_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[123]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_01435_),
    .QN(_00553_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[124]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_01436_),
    .QN(_00552_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[125]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .D(_01437_),
    .QN(_00551_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[126]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .D(_01438_),
    .QN(_00550_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[127]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_01439_),
    .QN(_00549_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[12]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .D(_01440_),
    .QN(_00548_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[13]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .D(_01441_),
    .QN(_00547_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[14]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .D(_01442_),
    .QN(_00546_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[15]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .D(_01443_),
    .QN(_00545_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[16]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .D(_01444_),
    .QN(_00466_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[17]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .D(_01445_),
    .QN(_00465_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[18]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .D(_01446_),
    .QN(_00467_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[19]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .D(_01447_),
    .QN(_00544_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[1]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .D(_01448_),
    .QN(_00408_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[20]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .D(_01449_),
    .QN(_00543_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[21]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .D(_01450_),
    .QN(_00542_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[22]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .D(_01451_),
    .QN(_00541_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[23]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .D(_01452_),
    .QN(_00540_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[24]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .D(_01453_),
    .QN(_00454_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[25]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .D(_01454_),
    .QN(_00453_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[26]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .D(_01455_),
    .QN(_00455_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[27]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .D(_01456_),
    .QN(_00539_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[28]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .D(_01457_),
    .QN(_00538_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[29]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .D(_01458_),
    .QN(_00537_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[2]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .D(_01459_),
    .QN(_00410_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[30]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .D(_01460_),
    .QN(_00536_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[31]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .D(_01461_),
    .QN(_00535_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[32]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .D(_01462_),
    .QN(_00406_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[33]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .D(_01463_),
    .QN(_00405_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[34]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .D(_01464_),
    .QN(_00407_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[35]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .D(_01465_),
    .QN(_00534_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[36]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .D(_01466_),
    .QN(_00533_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[37]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .D(_01467_),
    .QN(_00532_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[38]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .D(_01468_),
    .QN(_00531_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[39]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .D(_01469_),
    .QN(_00530_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[3]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .D(_01470_),
    .QN(_00529_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[40]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_01471_),
    .QN(_00475_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[41]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_01472_),
    .QN(_00474_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[42]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_01473_),
    .QN(_00476_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[43]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_01474_),
    .QN(_00528_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[44]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_01475_),
    .QN(_00527_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[45]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_01476_),
    .QN(_00526_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[46]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_01477_),
    .QN(_00525_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[47]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_01478_),
    .QN(_00524_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[48]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .D(_01479_),
    .QN(_00463_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[49]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .D(_01480_),
    .QN(_00462_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[4]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .D(_01481_),
    .QN(_00523_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[50]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .D(_01482_),
    .QN(_00464_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[51]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .D(_01483_),
    .QN(_00522_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[52]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .D(_01484_),
    .QN(_00521_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[53]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .D(_01485_),
    .QN(_00520_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[54]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_01486_),
    .QN(_00519_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[55]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .D(_01487_),
    .QN(_00518_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[56]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .D(_01488_),
    .QN(_00451_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[57]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .D(_01489_),
    .QN(_00450_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[58]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_01490_),
    .QN(_00452_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[59]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .D(_01491_),
    .QN(_00517_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[5]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .D(_01492_),
    .QN(_00516_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[60]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_01493_),
    .QN(_00515_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[61]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_01494_),
    .QN(_00514_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[62]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_01495_),
    .QN(_00513_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[63]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .D(_01496_),
    .QN(_00512_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[64]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .D(_01497_),
    .QN(_00484_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[65]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .D(_01498_),
    .QN(_00483_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[66]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_01499_),
    .QN(_00485_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[67]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .D(_01500_),
    .QN(_00511_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[68]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .D(_01501_),
    .QN(_00510_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[69]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .D(_01502_),
    .QN(_00509_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[6]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_01503_),
    .QN(_00508_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[70]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .D(_01504_),
    .QN(_00507_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[71]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .D(_01505_),
    .QN(_00506_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[72]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .D(_01506_),
    .QN(_00472_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[73]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .D(_01507_),
    .QN(_00471_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[74]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .D(_01508_),
    .QN(_00473_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[75]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .D(_01509_),
    .QN(_00505_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[76]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .D(_01510_),
    .QN(_00504_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[77]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .D(_01511_),
    .QN(_00503_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[78]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .D(_01512_),
    .QN(_00502_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[79]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .D(_01513_),
    .QN(_00501_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[7]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .D(_01514_),
    .QN(_00500_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[80]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .D(_01515_),
    .QN(_00460_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[81]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .D(_01516_),
    .QN(_00459_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[82]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .D(_01517_),
    .QN(_00461_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[83]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .D(_01518_),
    .QN(_00499_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[84]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .D(_01519_),
    .QN(_00498_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[85]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .D(_01520_),
    .QN(_00497_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[86]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .D(_01521_),
    .QN(_00496_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[87]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .D(_01522_),
    .QN(_00495_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[88]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .D(_01523_),
    .QN(_00448_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[89]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .D(_01524_),
    .QN(_00447_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[8]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_01525_),
    .QN(_00478_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[90]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .D(_01526_),
    .QN(_00449_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[91]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .D(_01527_),
    .QN(_00494_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[92]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .D(_01528_),
    .QN(_00493_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[93]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .D(_01529_),
    .QN(_00492_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[94]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .D(_01530_),
    .QN(_00491_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[95]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .D(_01531_),
    .QN(_00490_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[96]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_01532_),
    .QN(_00481_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[97]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_01533_),
    .QN(_00480_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[98]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .D(_01534_),
    .QN(_00482_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[99]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .D(_01535_),
    .QN(_00489_));
 DFFHQNx1_ASAP7_75t_R \text_in_r[9]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .D(_01536_),
    .QN(_00477_));
 DFFHQNx1_ASAP7_75t_R \text_out[0]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .D(_00265_),
    .QN(_00702_));
 DFFHQNx1_ASAP7_75t_R \text_out[100]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .D(_00165_),
    .QN(_00703_));
 DFFHQNx1_ASAP7_75t_R \text_out[101]$_DFF_P_  (.CLK(clknet_leaf_16_clk),
    .D(_00166_),
    .QN(_00704_));
 DFFHQNx1_ASAP7_75t_R \text_out[102]$_DFF_P_  (.CLK(clknet_leaf_12_clk),
    .D(_00167_),
    .QN(_00705_));
 DFFHQNx1_ASAP7_75t_R \text_out[103]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .D(_00168_),
    .QN(_00706_));
 DFFHQNx1_ASAP7_75t_R \text_out[104]$_DFF_P_  (.CLK(clknet_leaf_15_clk),
    .D(_00169_),
    .QN(_00707_));
 DFFHQNx1_ASAP7_75t_R \text_out[105]$_DFF_P_  (.CLK(clknet_leaf_15_clk),
    .D(_00170_),
    .QN(_00708_));
 DFFHQNx1_ASAP7_75t_R \text_out[106]$_DFF_P_  (.CLK(clknet_leaf_15_clk),
    .D(_00171_),
    .QN(_00709_));
 DFFHQNx1_ASAP7_75t_R \text_out[107]$_DFF_P_  (.CLK(clknet_leaf_15_clk),
    .D(_00172_),
    .QN(_00710_));
 DFFHQNx1_ASAP7_75t_R \text_out[108]$_DFF_P_  (.CLK(clknet_leaf_17_clk),
    .D(_00173_),
    .QN(_00711_));
 DFFHQNx1_ASAP7_75t_R \text_out[109]$_DFF_P_  (.CLK(clknet_leaf_17_clk),
    .D(_00174_),
    .QN(_00712_));
 DFFHQNx1_ASAP7_75t_R \text_out[10]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .D(_00195_),
    .QN(_00713_));
 DFFHQNx1_ASAP7_75t_R \text_out[110]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .D(_00175_),
    .QN(_00714_));
 DFFHQNx1_ASAP7_75t_R \text_out[111]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .D(_00176_),
    .QN(_00715_));
 DFFHQNx1_ASAP7_75t_R \text_out[112]$_DFF_P_  (.CLK(clknet_leaf_26_clk),
    .D(_00177_),
    .QN(_00716_));
 DFFHQNx1_ASAP7_75t_R \text_out[113]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .D(_00178_),
    .QN(_00717_));
 DFFHQNx1_ASAP7_75t_R \text_out[114]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .D(_00179_),
    .QN(_00718_));
 DFFHQNx1_ASAP7_75t_R \text_out[115]$_DFF_P_  (.CLK(clknet_leaf_22_clk),
    .D(_00180_),
    .QN(_00719_));
 DFFHQNx1_ASAP7_75t_R \text_out[116]$_DFF_P_  (.CLK(clknet_leaf_22_clk),
    .D(_00181_),
    .QN(_00720_));
 DFFHQNx1_ASAP7_75t_R \text_out[117]$_DFF_P_  (.CLK(clknet_leaf_22_clk),
    .D(_00182_),
    .QN(_00721_));
 DFFHQNx1_ASAP7_75t_R \text_out[118]$_DFF_P_  (.CLK(clknet_leaf_22_clk),
    .D(_00183_),
    .QN(_00722_));
 DFFHQNx1_ASAP7_75t_R \text_out[119]$_DFF_P_  (.CLK(clknet_leaf_16_clk),
    .D(_00184_),
    .QN(_00723_));
 DFFHQNx1_ASAP7_75t_R \text_out[11]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .D(_00196_),
    .QN(_00724_));
 DFFHQNx1_ASAP7_75t_R \text_out[120]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .D(_00185_),
    .QN(_00725_));
 DFFHQNx1_ASAP7_75t_R \text_out[121]$_DFF_P_  (.CLK(clknet_leaf_22_clk),
    .D(_00186_),
    .QN(_00726_));
 DFFHQNx1_ASAP7_75t_R \text_out[122]$_DFF_P_  (.CLK(clknet_leaf_24_clk),
    .D(_00187_),
    .QN(_00727_));
 DFFHQNx1_ASAP7_75t_R \text_out[123]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .D(_00188_),
    .QN(_00728_));
 DFFHQNx1_ASAP7_75t_R \text_out[124]$_DFF_P_  (.CLK(clknet_leaf_25_clk),
    .D(_00189_),
    .QN(_00729_));
 DFFHQNx1_ASAP7_75t_R \text_out[125]$_DFF_P_  (.CLK(clknet_leaf_24_clk),
    .D(_00190_),
    .QN(_00730_));
 DFFHQNx1_ASAP7_75t_R \text_out[126]$_DFF_P_  (.CLK(clknet_leaf_26_clk),
    .D(_00191_),
    .QN(_00731_));
 DFFHQNx1_ASAP7_75t_R \text_out[127]$_DFF_P_  (.CLK(clknet_leaf_22_clk),
    .D(_00192_),
    .QN(_00732_));
 DFFHQNx1_ASAP7_75t_R \text_out[12]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .D(_00197_),
    .QN(_00733_));
 DFFHQNx1_ASAP7_75t_R \text_out[13]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .D(_00198_),
    .QN(_00734_));
 DFFHQNx1_ASAP7_75t_R \text_out[14]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .D(_00199_),
    .QN(_00735_));
 DFFHQNx1_ASAP7_75t_R \text_out[15]$_DFF_P_  (.CLK(clknet_leaf_34_clk),
    .D(_00200_),
    .QN(_00736_));
 DFFHQNx1_ASAP7_75t_R \text_out[16]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .D(_00201_),
    .QN(_00737_));
 DFFHQNx1_ASAP7_75t_R \text_out[17]$_DFF_P_  (.CLK(clknet_leaf_30_clk),
    .D(_00202_),
    .QN(_00738_));
 DFFHQNx1_ASAP7_75t_R \text_out[18]$_DFF_P_  (.CLK(clknet_leaf_33_clk),
    .D(_00203_),
    .QN(_00739_));
 DFFHQNx1_ASAP7_75t_R \text_out[19]$_DFF_P_  (.CLK(clknet_leaf_30_clk),
    .D(_00204_),
    .QN(_00740_));
 DFFHQNx1_ASAP7_75t_R \text_out[1]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .D(_00266_),
    .QN(_00741_));
 DFFHQNx1_ASAP7_75t_R \text_out[20]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .D(_00205_),
    .QN(_00742_));
 DFFHQNx1_ASAP7_75t_R \text_out[21]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .D(_00206_),
    .QN(_00743_));
 DFFHQNx1_ASAP7_75t_R \text_out[22]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .D(_00207_),
    .QN(_00744_));
 DFFHQNx1_ASAP7_75t_R \text_out[23]$_DFF_P_  (.CLK(clknet_leaf_32_clk),
    .D(_00208_),
    .QN(_00745_));
 DFFHQNx1_ASAP7_75t_R \text_out[24]$_DFF_P_  (.CLK(clknet_leaf_33_clk),
    .D(_00209_),
    .QN(_00746_));
 DFFHQNx1_ASAP7_75t_R \text_out[25]$_DFF_P_  (.CLK(clknet_leaf_34_clk),
    .D(_00210_),
    .QN(_00747_));
 DFFHQNx1_ASAP7_75t_R \text_out[26]$_DFF_P_  (.CLK(clknet_leaf_33_clk),
    .D(_00211_),
    .QN(_00748_));
 DFFHQNx1_ASAP7_75t_R \text_out[27]$_DFF_P_  (.CLK(clknet_leaf_33_clk),
    .D(_00212_),
    .QN(_00749_));
 DFFHQNx1_ASAP7_75t_R \text_out[28]$_DFF_P_  (.CLK(clknet_leaf_34_clk),
    .D(_00213_),
    .QN(_00750_));
 DFFHQNx1_ASAP7_75t_R \text_out[29]$_DFF_P_  (.CLK(clknet_leaf_34_clk),
    .D(_00214_),
    .QN(_00751_));
 DFFHQNx1_ASAP7_75t_R \text_out[2]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .D(_00267_),
    .QN(_00752_));
 DFFHQNx1_ASAP7_75t_R \text_out[30]$_DFF_P_  (.CLK(clknet_leaf_34_clk),
    .D(_00215_),
    .QN(_00753_));
 DFFHQNx1_ASAP7_75t_R \text_out[31]$_DFF_P_  (.CLK(clknet_leaf_34_clk),
    .D(_00216_),
    .QN(_00754_));
 DFFHQNx1_ASAP7_75t_R \text_out[32]$_DFF_P_  (.CLK(clknet_leaf_8_clk),
    .D(_00217_),
    .QN(_00755_));
 DFFHQNx1_ASAP7_75t_R \text_out[33]$_DFF_P_  (.CLK(clknet_leaf_8_clk),
    .D(_00218_),
    .QN(_00756_));
 DFFHQNx1_ASAP7_75t_R \text_out[34]$_DFF_P_  (.CLK(clknet_leaf_8_clk),
    .D(_00219_),
    .QN(_00757_));
 DFFHQNx1_ASAP7_75t_R \text_out[35]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .D(_00220_),
    .QN(_00758_));
 DFFHQNx1_ASAP7_75t_R \text_out[36]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .D(_00221_),
    .QN(_00759_));
 DFFHQNx1_ASAP7_75t_R \text_out[37]$_DFF_P_  (.CLK(clknet_leaf_8_clk),
    .D(_00222_),
    .QN(_00760_));
 DFFHQNx1_ASAP7_75t_R \text_out[38]$_DFF_P_  (.CLK(clknet_leaf_8_clk),
    .D(_00223_),
    .QN(_00761_));
 DFFHQNx1_ASAP7_75t_R \text_out[39]$_DFF_P_  (.CLK(clknet_leaf_8_clk),
    .D(_00224_),
    .QN(_00762_));
 DFFHQNx1_ASAP7_75t_R \text_out[3]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .D(_00268_),
    .QN(_00763_));
 DFFHQNx1_ASAP7_75t_R \text_out[40]$_DFF_P_  (.CLK(clknet_leaf_14_clk),
    .D(_00225_),
    .QN(_00764_));
 DFFHQNx1_ASAP7_75t_R \text_out[41]$_DFF_P_  (.CLK(clknet_leaf_14_clk),
    .D(_00226_),
    .QN(_00765_));
 DFFHQNx1_ASAP7_75t_R \text_out[42]$_DFF_P_  (.CLK(clknet_leaf_13_clk),
    .D(_00227_),
    .QN(_00766_));
 DFFHQNx1_ASAP7_75t_R \text_out[43]$_DFF_P_  (.CLK(clknet_leaf_13_clk),
    .D(_00228_),
    .QN(_00767_));
 DFFHQNx1_ASAP7_75t_R \text_out[44]$_DFF_P_  (.CLK(clknet_leaf_14_clk),
    .D(_00229_),
    .QN(_00768_));
 DFFHQNx1_ASAP7_75t_R \text_out[45]$_DFF_P_  (.CLK(clknet_leaf_14_clk),
    .D(_00230_),
    .QN(_00769_));
 DFFHQNx1_ASAP7_75t_R \text_out[46]$_DFF_P_  (.CLK(clknet_leaf_14_clk),
    .D(_00231_),
    .QN(_00770_));
 DFFHQNx1_ASAP7_75t_R \text_out[47]$_DFF_P_  (.CLK(clknet_leaf_14_clk),
    .D(_00232_),
    .QN(_00771_));
 DFFHQNx1_ASAP7_75t_R \text_out[48]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .D(_00233_),
    .QN(_00772_));
 DFFHQNx1_ASAP7_75t_R \text_out[49]$_DFF_P_  (.CLK(clknet_leaf_27_clk),
    .D(_00234_),
    .QN(_00773_));
 DFFHQNx1_ASAP7_75t_R \text_out[4]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .D(_00269_),
    .QN(_00774_));
 DFFHQNx1_ASAP7_75t_R \text_out[50]$_DFF_P_  (.CLK(clknet_leaf_26_clk),
    .D(_00235_),
    .QN(_00775_));
 DFFHQNx1_ASAP7_75t_R \text_out[51]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .D(_00236_),
    .QN(_00776_));
 DFFHQNx1_ASAP7_75t_R \text_out[52]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .D(_00237_),
    .QN(_00777_));
 DFFHQNx1_ASAP7_75t_R \text_out[53]$_DFF_P_  (.CLK(clknet_leaf_30_clk),
    .D(_00238_),
    .QN(_00778_));
 DFFHQNx1_ASAP7_75t_R \text_out[54]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .D(_00239_),
    .QN(_00779_));
 DFFHQNx1_ASAP7_75t_R \text_out[55]$_DFF_P_  (.CLK(clknet_leaf_19_clk),
    .D(_00240_),
    .QN(_00780_));
 DFFHQNx1_ASAP7_75t_R \text_out[56]$_DFF_P_  (.CLK(clknet_leaf_8_clk),
    .D(_00241_),
    .QN(_00781_));
 DFFHQNx1_ASAP7_75t_R \text_out[57]$_DFF_P_  (.CLK(clknet_leaf_13_clk),
    .D(_00242_),
    .QN(_00782_));
 DFFHQNx1_ASAP7_75t_R \text_out[58]$_DFF_P_  (.CLK(clknet_leaf_13_clk),
    .D(_00243_),
    .QN(_00783_));
 DFFHQNx1_ASAP7_75t_R \text_out[59]$_DFF_P_  (.CLK(clknet_leaf_13_clk),
    .D(_00244_),
    .QN(_00784_));
 DFFHQNx1_ASAP7_75t_R \text_out[5]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .D(_00270_),
    .QN(_00785_));
 DFFHQNx1_ASAP7_75t_R \text_out[60]$_DFF_P_  (.CLK(clknet_leaf_13_clk),
    .D(_00245_),
    .QN(_00786_));
 DFFHQNx1_ASAP7_75t_R \text_out[61]$_DFF_P_  (.CLK(clknet_leaf_19_clk),
    .D(_00246_),
    .QN(_00787_));
 DFFHQNx1_ASAP7_75t_R \text_out[62]$_DFF_P_  (.CLK(clknet_leaf_13_clk),
    .D(_00247_),
    .QN(_00788_));
 DFFHQNx1_ASAP7_75t_R \text_out[63]$_DFF_P_  (.CLK(clknet_leaf_13_clk),
    .D(_00248_),
    .QN(_00789_));
 DFFHQNx1_ASAP7_75t_R \text_out[64]$_DFF_P_  (.CLK(clknet_leaf_16_clk),
    .D(_00249_),
    .QN(_00790_));
 DFFHQNx1_ASAP7_75t_R \text_out[65]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .D(_00250_),
    .QN(_00791_));
 DFFHQNx1_ASAP7_75t_R \text_out[66]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .D(_00251_),
    .QN(_00792_));
 DFFHQNx1_ASAP7_75t_R \text_out[67]$_DFF_P_  (.CLK(clknet_leaf_16_clk),
    .D(_00252_),
    .QN(_00793_));
 DFFHQNx1_ASAP7_75t_R \text_out[68]$_DFF_P_  (.CLK(clknet_leaf_17_clk),
    .D(_00253_),
    .QN(_00794_));
 DFFHQNx1_ASAP7_75t_R \text_out[69]$_DFF_P_  (.CLK(clknet_leaf_22_clk),
    .D(_00254_),
    .QN(_00795_));
 DFFHQNx1_ASAP7_75t_R \text_out[6]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .D(_00271_),
    .QN(_00796_));
 DFFHQNx1_ASAP7_75t_R \text_out[70]$_DFF_P_  (.CLK(clknet_leaf_16_clk),
    .D(_00255_),
    .QN(_00797_));
 DFFHQNx1_ASAP7_75t_R \text_out[71]$_DFF_P_  (.CLK(clknet_leaf_17_clk),
    .D(_00256_),
    .QN(_00798_));
 DFFHQNx1_ASAP7_75t_R \text_out[72]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .D(_00257_),
    .QN(_00799_));
 DFFHQNx1_ASAP7_75t_R \text_out[73]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .D(_00258_),
    .QN(_00800_));
 DFFHQNx1_ASAP7_75t_R \text_out[74]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .D(_00259_),
    .QN(_00801_));
 DFFHQNx1_ASAP7_75t_R \text_out[75]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .D(_00260_),
    .QN(_00802_));
 DFFHQNx1_ASAP7_75t_R \text_out[76]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .D(_00261_),
    .QN(_00803_));
 DFFHQNx1_ASAP7_75t_R \text_out[77]$_DFF_P_  (.CLK(clknet_leaf_22_clk),
    .D(_00262_),
    .QN(_00804_));
 DFFHQNx1_ASAP7_75t_R \text_out[78]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .D(_00263_),
    .QN(_00805_));
 DFFHQNx1_ASAP7_75t_R \text_out[79]$_DFF_P_  (.CLK(clknet_leaf_22_clk),
    .D(_00264_),
    .QN(_00806_));
 DFFHQNx1_ASAP7_75t_R \text_out[7]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .D(_00272_),
    .QN(_00807_));
 DFFHQNx1_ASAP7_75t_R \text_out[80]$_DFF_P_  (.CLK(clknet_leaf_26_clk),
    .D(_00273_),
    .QN(_00808_));
 DFFHQNx1_ASAP7_75t_R \text_out[81]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .D(_00274_),
    .QN(_00809_));
 DFFHQNx1_ASAP7_75t_R \text_out[82]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .D(_00275_),
    .QN(_00810_));
 DFFHQNx1_ASAP7_75t_R \text_out[83]$_DFF_P_  (.CLK(clknet_leaf_26_clk),
    .D(_00276_),
    .QN(_00811_));
 DFFHQNx1_ASAP7_75t_R \text_out[84]$_DFF_P_  (.CLK(clknet_leaf_22_clk),
    .D(_00277_),
    .QN(_00812_));
 DFFHQNx1_ASAP7_75t_R \text_out[85]$_DFF_P_  (.CLK(clknet_leaf_24_clk),
    .D(_00278_),
    .QN(_00813_));
 DFFHQNx1_ASAP7_75t_R \text_out[86]$_DFF_P_  (.CLK(clknet_leaf_22_clk),
    .D(_00279_),
    .QN(_00814_));
 DFFHQNx1_ASAP7_75t_R \text_out[87]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .D(_00280_),
    .QN(_00815_));
 DFFHQNx1_ASAP7_75t_R \text_out[88]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .D(_00281_),
    .QN(_00816_));
 DFFHQNx1_ASAP7_75t_R \text_out[89]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .D(_00282_),
    .QN(_00817_));
 DFFHQNx1_ASAP7_75t_R \text_out[8]$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .D(_00193_),
    .QN(_00818_));
 DFFHQNx1_ASAP7_75t_R \text_out[90]$_DFF_P_  (.CLK(clknet_leaf_24_clk),
    .D(_00283_),
    .QN(_00819_));
 DFFHQNx1_ASAP7_75t_R \text_out[91]$_DFF_P_  (.CLK(clknet_leaf_25_clk),
    .D(_00284_),
    .QN(_00820_));
 DFFHQNx1_ASAP7_75t_R \text_out[92]$_DFF_P_  (.CLK(clknet_leaf_25_clk),
    .D(_00285_),
    .QN(_00821_));
 DFFHQNx1_ASAP7_75t_R \text_out[93]$_DFF_P_  (.CLK(clknet_leaf_24_clk),
    .D(_00286_),
    .QN(_00822_));
 DFFHQNx1_ASAP7_75t_R \text_out[94]$_DFF_P_  (.CLK(clknet_leaf_24_clk),
    .D(_00287_),
    .QN(_00823_));
 DFFHQNx1_ASAP7_75t_R \text_out[95]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .D(_00288_),
    .QN(_00824_));
 DFFHQNx1_ASAP7_75t_R \text_out[96]$_DFF_P_  (.CLK(clknet_leaf_19_clk),
    .D(_00161_),
    .QN(_00825_));
 DFFHQNx1_ASAP7_75t_R \text_out[97]$_DFF_P_  (.CLK(clknet_leaf_16_clk),
    .D(_00162_),
    .QN(_00826_));
 DFFHQNx1_ASAP7_75t_R \text_out[98]$_DFF_P_  (.CLK(clknet_leaf_15_clk),
    .D(_00163_),
    .QN(_00827_));
 DFFHQNx1_ASAP7_75t_R \text_out[99]$_DFF_P_  (.CLK(clknet_leaf_11_clk),
    .D(_00164_),
    .QN(_00828_));
 DFFHQNx1_ASAP7_75t_R \text_out[9]$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .D(_00194_),
    .QN(_00488_));
 DFFHQNx1_ASAP7_75t_R \u0.r0.out[24]$_SDFF_PP1_  (.CLK(clknet_leaf_31_clk),
    .D(_01537_),
    .QN(_00413_));
 DFFHQNx1_ASAP7_75t_R \u0.r0.out[25]$_SDFF_PP0_  (.CLK(clknet_leaf_29_clk),
    .D(_01538_),
    .QN(_00414_));
 DFFHQNx1_ASAP7_75t_R \u0.r0.out[26]$_SDFF_PP0_  (.CLK(clknet_leaf_30_clk),
    .D(_01539_),
    .QN(_00415_));
 DFFHQNx1_ASAP7_75t_R \u0.r0.out[27]$_SDFF_PP0_  (.CLK(clknet_leaf_31_clk),
    .D(_01540_),
    .QN(_00416_));
 DFFHQNx1_ASAP7_75t_R \u0.r0.out[28]$_SDFF_PP0_  (.CLK(clknet_leaf_31_clk),
    .D(_01541_),
    .QN(_00417_));
 DFFHQNx1_ASAP7_75t_R \u0.r0.out[29]$_SDFF_PP0_  (.CLK(clknet_leaf_31_clk),
    .D(_01542_),
    .QN(_00418_));
 DFFHQNx1_ASAP7_75t_R \u0.r0.out[30]$_SDFF_PP0_  (.CLK(clknet_leaf_27_clk),
    .D(_01543_),
    .QN(_00419_));
 DFFHQNx1_ASAP7_75t_R \u0.r0.out[31]$_SDFF_PP0_  (.CLK(clknet_leaf_31_clk),
    .D(_01544_),
    .QN(_00420_));
 DFFHQNx1_ASAP7_75t_R \u0.r0.rcnt[0]$_SDFF_PP0_  (.CLK(clknet_leaf_31_clk),
    .D(_01545_),
    .QN(\u0.r0.rcnt_next[0] ));
 DFFHQNx1_ASAP7_75t_R \u0.r0.rcnt[1]$_SDFF_PP0_  (.CLK(clknet_leaf_31_clk),
    .D(_01546_),
    .QN(_00965_));
 DFFHQNx1_ASAP7_75t_R \u0.r0.rcnt[2]$_SDFF_PP0_  (.CLK(clknet_leaf_31_clk),
    .D(_01547_),
    .QN(_00487_));
 DFFHQNx1_ASAP7_75t_R \u0.r0.rcnt[3]$_SDFF_PP0_  (.CLK(clknet_leaf_31_clk),
    .D(_01548_),
    .QN(_00829_));
 DFFHQNx1_ASAP7_75t_R \u0.u0.d[0]$_DFF_P_  (.CLK(clknet_leaf_32_clk),
    .D(_00000_),
    .QN(_00830_));
 DFFHQNx1_ASAP7_75t_R \u0.u0.d[1]$_DFF_P_  (.CLK(clknet_leaf_31_clk),
    .D(_00001_),
    .QN(_00831_));
 DFFHQNx1_ASAP7_75t_R \u0.u0.d[2]$_DFF_P_  (.CLK(clknet_leaf_31_clk),
    .D(_00002_),
    .QN(_00832_));
 DFFHQNx1_ASAP7_75t_R \u0.u0.d[3]$_DFF_P_  (.CLK(clknet_leaf_32_clk),
    .D(_00003_),
    .QN(_00833_));
 DFFHQNx1_ASAP7_75t_R \u0.u0.d[4]$_DFF_P_  (.CLK(clknet_leaf_32_clk),
    .D(_00004_),
    .QN(_00834_));
 DFFHQNx1_ASAP7_75t_R \u0.u0.d[5]$_DFF_P_  (.CLK(clknet_leaf_32_clk),
    .D(_00005_),
    .QN(_00835_));
 DFFHQNx1_ASAP7_75t_R \u0.u0.d[6]$_DFF_P_  (.CLK(clknet_leaf_27_clk),
    .D(_00006_),
    .QN(_00836_));
 DFFHQNx1_ASAP7_75t_R \u0.u0.d[7]$_DFF_P_  (.CLK(clknet_leaf_27_clk),
    .D(_00007_),
    .QN(_00837_));
 DFFHQNx1_ASAP7_75t_R \u0.u1.d[0]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .D(_00008_),
    .QN(_00437_));
 DFFHQNx1_ASAP7_75t_R \u0.u1.d[1]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .D(_00009_),
    .QN(_00438_));
 DFFHQNx1_ASAP7_75t_R \u0.u1.d[2]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .D(_00010_),
    .QN(_00412_));
 DFFHQNx1_ASAP7_75t_R \u0.u1.d[3]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .D(_00011_),
    .QN(_00439_));
 DFFHQNx1_ASAP7_75t_R \u0.u1.d[4]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .D(_00012_),
    .QN(_00440_));
 DFFHQNx1_ASAP7_75t_R \u0.u1.d[5]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .D(_00013_),
    .QN(_00441_));
 DFFHQNx1_ASAP7_75t_R \u0.u1.d[6]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .D(_00014_),
    .QN(_00442_));
 DFFHQNx1_ASAP7_75t_R \u0.u1.d[7]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .D(_00015_),
    .QN(_00443_));
 DFFHQNx1_ASAP7_75t_R \u0.u2.d[0]$_DFF_P_  (.CLK(clknet_leaf_10_clk),
    .D(_00016_),
    .QN(_00429_));
 DFFHQNx1_ASAP7_75t_R \u0.u2.d[1]$_DFF_P_  (.CLK(clknet_leaf_10_clk),
    .D(_00017_),
    .QN(_00430_));
 DFFHQNx1_ASAP7_75t_R \u0.u2.d[2]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .D(_00018_),
    .QN(_00431_));
 DFFHQNx1_ASAP7_75t_R \u0.u2.d[3]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .D(_00019_),
    .QN(_00432_));
 DFFHQNx1_ASAP7_75t_R \u0.u2.d[4]$_DFF_P_  (.CLK(clknet_leaf_10_clk),
    .D(_00020_),
    .QN(_00433_));
 DFFHQNx1_ASAP7_75t_R \u0.u2.d[5]$_DFF_P_  (.CLK(clknet_leaf_10_clk),
    .D(_00021_),
    .QN(_00434_));
 DFFHQNx1_ASAP7_75t_R \u0.u2.d[6]$_DFF_P_  (.CLK(clknet_leaf_10_clk),
    .D(_00022_),
    .QN(_00435_));
 DFFHQNx1_ASAP7_75t_R \u0.u2.d[7]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .D(_00023_),
    .QN(_00436_));
 DFFHQNx1_ASAP7_75t_R \u0.u3.d[0]$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .D(_00024_),
    .QN(_00421_));
 DFFHQNx1_ASAP7_75t_R \u0.u3.d[1]$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .D(_00025_),
    .QN(_00422_));
 DFFHQNx1_ASAP7_75t_R \u0.u3.d[2]$_DFF_P_  (.CLK(clknet_leaf_34_clk),
    .D(_00026_),
    .QN(_00423_));
 DFFHQNx1_ASAP7_75t_R \u0.u3.d[3]$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .D(_00027_),
    .QN(_00424_));
 DFFHQNx1_ASAP7_75t_R \u0.u3.d[4]$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .D(_00028_),
    .QN(_00425_));
 DFFHQNx1_ASAP7_75t_R \u0.u3.d[5]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .D(_00029_),
    .QN(_00426_));
 DFFHQNx1_ASAP7_75t_R \u0.u3.d[6]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .D(_00030_),
    .QN(_00427_));
 DFFHQNx1_ASAP7_75t_R \u0.u3.d[7]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .D(_00031_),
    .QN(_00428_));
 DFFHQNx1_ASAP7_75t_R \u0.w[0][0]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .D(_00289_),
    .QN(_00838_));
 DFFHQNx1_ASAP7_75t_R \u0.w[0][10]$_DFF_P_  (.CLK(clknet_leaf_9_clk),
    .D(_00290_),
    .QN(_00839_));
 DFFHQNx1_ASAP7_75t_R \u0.w[0][11]$_DFF_P_  (.CLK(clknet_leaf_13_clk),
    .D(_00291_),
    .QN(_00840_));
 DFFHQNx1_ASAP7_75t_R \u0.w[0][12]$_DFF_P_  (.CLK(clknet_leaf_9_clk),
    .D(_00292_),
    .QN(_00841_));
 DFFHQNx1_ASAP7_75t_R \u0.w[0][13]$_DFF_P_  (.CLK(clknet_leaf_10_clk),
    .D(_00293_),
    .QN(_00842_));
 DFFHQNx1_ASAP7_75t_R \u0.w[0][14]$_DFF_P_  (.CLK(clknet_leaf_9_clk),
    .D(_00294_),
    .QN(_00843_));
 DFFHQNx1_ASAP7_75t_R \u0.w[0][15]$_DFF_P_  (.CLK(clknet_leaf_11_clk),
    .D(_00295_),
    .QN(_00844_));
 DFFHQNx1_ASAP7_75t_R \u0.w[0][16]$_DFF_P_  (.CLK(clknet_leaf_27_clk),
    .D(_00296_),
    .QN(_00845_));
 DFFHQNx1_ASAP7_75t_R \u0.w[0][17]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .D(_00297_),
    .QN(_00846_));
 DFFHQNx1_ASAP7_75t_R \u0.w[0][18]$_DFF_P_  (.CLK(clknet_leaf_2_clk),
    .D(_00298_),
    .QN(_00847_));
 DFFHQNx1_ASAP7_75t_R \u0.w[0][19]$_DFF_P_  (.CLK(clknet_leaf_27_clk),
    .D(_00299_),
    .QN(_00848_));
 DFFHQNx2_ASAP7_75t_R \u0.w[0][1]$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .D(_00300_),
    .QN(_00849_));
 DFFHQNx1_ASAP7_75t_R \u0.w[0][20]$_DFF_P_  (.CLK(clknet_leaf_22_clk),
    .D(_00301_),
    .QN(_00850_));
 DFFHQNx1_ASAP7_75t_R \u0.w[0][21]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .D(_00302_),
    .QN(_00851_));
 DFFHQNx1_ASAP7_75t_R \u0.w[0][22]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .D(_00303_),
    .QN(_00852_));
 DFFHQNx1_ASAP7_75t_R \u0.w[0][23]$_DFF_P_  (.CLK(clknet_leaf_26_clk),
    .D(_00304_),
    .QN(_00853_));
 DFFHQNx2_ASAP7_75t_R \u0.w[0][24]$_DFF_P_  (.CLK(clknet_leaf_32_clk),
    .D(_00305_),
    .QN(_00854_));
 DFFHQNx1_ASAP7_75t_R \u0.w[0][25]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .D(_00306_),
    .QN(_00855_));
 DFFHQNx1_ASAP7_75t_R \u0.w[0][26]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .D(_00307_),
    .QN(_00856_));
 DFFHQNx1_ASAP7_75t_R \u0.w[0][27]$_DFF_P_  (.CLK(clknet_leaf_31_clk),
    .D(_00308_),
    .QN(_00857_));
 DFFHQNx1_ASAP7_75t_R \u0.w[0][28]$_DFF_P_  (.CLK(clknet_leaf_32_clk),
    .D(_00309_),
    .QN(_00858_));
 DFFHQNx1_ASAP7_75t_R \u0.w[0][29]$_DFF_P_  (.CLK(clknet_leaf_31_clk),
    .D(_00310_),
    .QN(_00859_));
 DFFHQNx1_ASAP7_75t_R \u0.w[0][2]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .D(_00311_),
    .QN(_00860_));
 DFFHQNx1_ASAP7_75t_R \u0.w[0][30]$_DFF_P_  (.CLK(clknet_leaf_27_clk),
    .D(_00312_),
    .QN(_00861_));
 DFFHQNx1_ASAP7_75t_R \u0.w[0][31]$_DFF_P_  (.CLK(clknet_leaf_27_clk),
    .D(_00313_),
    .QN(_00862_));
 DFFHQNx1_ASAP7_75t_R \u0.w[0][3]$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .D(_00314_),
    .QN(_00863_));
 DFFHQNx1_ASAP7_75t_R \u0.w[0][4]$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .D(_00315_),
    .QN(_00864_));
 DFFHQNx1_ASAP7_75t_R \u0.w[0][5]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .D(_00316_),
    .QN(_00865_));
 DFFHQNx1_ASAP7_75t_R \u0.w[0][6]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .D(_00317_),
    .QN(_00866_));
 DFFHQNx1_ASAP7_75t_R \u0.w[0][7]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .D(_00318_),
    .QN(_00867_));
 DFFHQNx1_ASAP7_75t_R \u0.w[0][8]$_DFF_P_  (.CLK(clknet_leaf_9_clk),
    .D(_00319_),
    .QN(_00868_));
 DFFHQNx1_ASAP7_75t_R \u0.w[0][9]$_DFF_P_  (.CLK(clknet_leaf_11_clk),
    .D(_00320_),
    .QN(_00869_));
 DFFHQNx1_ASAP7_75t_R \u0.w[1][0]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .D(_00321_),
    .QN(_00870_));
 DFFHQNx1_ASAP7_75t_R \u0.w[1][10]$_DFF_P_  (.CLK(clknet_leaf_9_clk),
    .D(_00322_),
    .QN(_00871_));
 DFFHQNx1_ASAP7_75t_R \u0.w[1][11]$_DFF_P_  (.CLK(clknet_leaf_13_clk),
    .D(_00323_),
    .QN(_00872_));
 DFFHQNx1_ASAP7_75t_R \u0.w[1][12]$_DFF_P_  (.CLK(clknet_leaf_9_clk),
    .D(_00324_),
    .QN(_00873_));
 DFFHQNx1_ASAP7_75t_R \u0.w[1][13]$_DFF_P_  (.CLK(clknet_leaf_2_clk),
    .D(_00325_),
    .QN(_00874_));
 DFFHQNx1_ASAP7_75t_R \u0.w[1][14]$_DFF_P_  (.CLK(clknet_leaf_2_clk),
    .D(_00326_),
    .QN(_00875_));
 DFFHQNx1_ASAP7_75t_R \u0.w[1][15]$_DFF_P_  (.CLK(clknet_leaf_19_clk),
    .D(_00327_),
    .QN(_00876_));
 DFFHQNx1_ASAP7_75t_R \u0.w[1][16]$_DFF_P_  (.CLK(clknet_leaf_27_clk),
    .D(_00328_),
    .QN(_00877_));
 DFFHQNx1_ASAP7_75t_R \u0.w[1][17]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .D(_00329_),
    .QN(_00878_));
 DFFHQNx1_ASAP7_75t_R \u0.w[1][18]$_DFF_P_  (.CLK(clknet_leaf_31_clk),
    .D(_00330_),
    .QN(_00879_));
 DFFHQNx1_ASAP7_75t_R \u0.w[1][19]$_DFF_P_  (.CLK(clknet_leaf_27_clk),
    .D(_00331_),
    .QN(_00880_));
 DFFHQNx1_ASAP7_75t_R \u0.w[1][1]$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .D(_00332_),
    .QN(_00881_));
 DFFHQNx1_ASAP7_75t_R \u0.w[1][20]$_DFF_P_  (.CLK(clknet_leaf_22_clk),
    .D(_00333_),
    .QN(_00882_));
 DFFHQNx1_ASAP7_75t_R \u0.w[1][21]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .D(_00334_),
    .QN(_00883_));
 DFFHQNx1_ASAP7_75t_R \u0.w[1][22]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .D(_00335_),
    .QN(_00884_));
 DFFHQNx1_ASAP7_75t_R \u0.w[1][23]$_DFF_P_  (.CLK(clknet_leaf_26_clk),
    .D(_00336_),
    .QN(_00885_));
 DFFHQNx1_ASAP7_75t_R \u0.w[1][24]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .D(_00337_),
    .QN(_00886_));
 DFFHQNx1_ASAP7_75t_R \u0.w[1][25]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .D(_00338_),
    .QN(_00887_));
 DFFHQNx1_ASAP7_75t_R \u0.w[1][26]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .D(_00339_),
    .QN(_00888_));
 DFFHQNx1_ASAP7_75t_R \u0.w[1][27]$_DFF_P_  (.CLK(clknet_leaf_31_clk),
    .D(_00340_),
    .QN(_00889_));
 DFFHQNx1_ASAP7_75t_R \u0.w[1][28]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .D(_00341_),
    .QN(_00890_));
 DFFHQNx1_ASAP7_75t_R \u0.w[1][29]$_DFF_P_  (.CLK(clknet_leaf_31_clk),
    .D(_00342_),
    .QN(_00891_));
 DFFHQNx1_ASAP7_75t_R \u0.w[1][2]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .D(_00343_),
    .QN(_00892_));
 DFFHQNx1_ASAP7_75t_R \u0.w[1][30]$_DFF_P_  (.CLK(clknet_leaf_27_clk),
    .D(_00344_),
    .QN(_00893_));
 DFFHQNx1_ASAP7_75t_R \u0.w[1][31]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .D(_00345_),
    .QN(_00894_));
 DFFHQNx1_ASAP7_75t_R \u0.w[1][3]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .D(_00346_),
    .QN(_00895_));
 DFFHQNx1_ASAP7_75t_R \u0.w[1][4]$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .D(_00347_),
    .QN(_00896_));
 DFFHQNx1_ASAP7_75t_R \u0.w[1][5]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .D(_00348_),
    .QN(_00897_));
 DFFHQNx1_ASAP7_75t_R \u0.w[1][6]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .D(_00349_),
    .QN(_00898_));
 DFFHQNx1_ASAP7_75t_R \u0.w[1][7]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .D(_00350_),
    .QN(_00899_));
 DFFHQNx1_ASAP7_75t_R \u0.w[1][8]$_DFF_P_  (.CLK(clknet_leaf_10_clk),
    .D(_00351_),
    .QN(_00900_));
 DFFHQNx1_ASAP7_75t_R \u0.w[1][9]$_DFF_P_  (.CLK(clknet_leaf_19_clk),
    .D(_00352_),
    .QN(_00901_));
 DFFHQNx1_ASAP7_75t_R \u0.w[2][0]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .D(_00353_),
    .QN(_00902_));
 DFFHQNx1_ASAP7_75t_R \u0.w[2][10]$_DFF_P_  (.CLK(clknet_leaf_9_clk),
    .D(_00354_),
    .QN(_00903_));
 DFFHQNx1_ASAP7_75t_R \u0.w[2][11]$_DFF_P_  (.CLK(clknet_leaf_9_clk),
    .D(_00355_),
    .QN(_00904_));
 DFFHQNx1_ASAP7_75t_R \u0.w[2][12]$_DFF_P_  (.CLK(clknet_leaf_10_clk),
    .D(_00356_),
    .QN(_00905_));
 DFFHQNx1_ASAP7_75t_R \u0.w[2][13]$_DFF_P_  (.CLK(clknet_leaf_2_clk),
    .D(_00357_),
    .QN(_00906_));
 DFFHQNx1_ASAP7_75t_R \u0.w[2][14]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .D(_00358_),
    .QN(_00907_));
 DFFHQNx1_ASAP7_75t_R \u0.w[2][15]$_DFF_P_  (.CLK(clknet_leaf_19_clk),
    .D(_00359_),
    .QN(_00908_));
 DFFHQNx1_ASAP7_75t_R \u0.w[2][16]$_DFF_P_  (.CLK(clknet_leaf_31_clk),
    .D(_00360_),
    .QN(_00909_));
 DFFHQNx1_ASAP7_75t_R \u0.w[2][17]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .D(_00361_),
    .QN(_00910_));
 DFFHQNx1_ASAP7_75t_R \u0.w[2][18]$_DFF_P_  (.CLK(clknet_leaf_31_clk),
    .D(_00362_),
    .QN(_00911_));
 DFFHQNx1_ASAP7_75t_R \u0.w[2][19]$_DFF_P_  (.CLK(clknet_leaf_27_clk),
    .D(_00363_),
    .QN(_00912_));
 DFFHQNx1_ASAP7_75t_R \u0.w[2][1]$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .D(_00364_),
    .QN(_00913_));
 DFFHQNx1_ASAP7_75t_R \u0.w[2][20]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .D(_00365_),
    .QN(_00914_));
 DFFHQNx1_ASAP7_75t_R \u0.w[2][21]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .D(_00366_),
    .QN(_00915_));
 DFFHQNx1_ASAP7_75t_R \u0.w[2][22]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .D(_00367_),
    .QN(_00916_));
 DFFHQNx1_ASAP7_75t_R \u0.w[2][23]$_DFF_P_  (.CLK(clknet_leaf_26_clk),
    .D(_00368_),
    .QN(_00917_));
 DFFHQNx1_ASAP7_75t_R \u0.w[2][24]$_DFF_P_  (.CLK(clknet_leaf_30_clk),
    .D(_00369_),
    .QN(_00918_));
 DFFHQNx1_ASAP7_75t_R \u0.w[2][25]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .D(_00370_),
    .QN(_00919_));
 DFFHQNx1_ASAP7_75t_R \u0.w[2][26]$_DFF_P_  (.CLK(clknet_leaf_30_clk),
    .D(_00371_),
    .QN(_00920_));
 DFFHQNx1_ASAP7_75t_R \u0.w[2][27]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .D(_00372_),
    .QN(_00921_));
 DFFHQNx1_ASAP7_75t_R \u0.w[2][28]$_DFF_P_  (.CLK(clknet_leaf_2_clk),
    .D(_00373_),
    .QN(_00922_));
 DFFHQNx1_ASAP7_75t_R \u0.w[2][29]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .D(_00374_),
    .QN(_00923_));
 DFFHQNx1_ASAP7_75t_R \u0.w[2][2]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .D(_00375_),
    .QN(_00924_));
 DFFHQNx1_ASAP7_75t_R \u0.w[2][30]$_DFF_P_  (.CLK(clknet_leaf_31_clk),
    .D(_00376_),
    .QN(_00925_));
 DFFHQNx1_ASAP7_75t_R \u0.w[2][31]$_DFF_P_  (.CLK(clknet_leaf_2_clk),
    .D(_00377_),
    .QN(_00926_));
 DFFHQNx1_ASAP7_75t_R \u0.w[2][3]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .D(_00378_),
    .QN(_00927_));
 DFFHQNx1_ASAP7_75t_R \u0.w[2][4]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .D(_00379_),
    .QN(_00928_));
 DFFHQNx1_ASAP7_75t_R \u0.w[2][5]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .D(_00380_),
    .QN(_00929_));
 DFFHQNx1_ASAP7_75t_R \u0.w[2][6]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .D(_00381_),
    .QN(_00930_));
 DFFHQNx1_ASAP7_75t_R \u0.w[2][7]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .D(_00382_),
    .QN(_00931_));
 DFFHQNx1_ASAP7_75t_R \u0.w[2][8]$_DFF_P_  (.CLK(clknet_leaf_9_clk),
    .D(_00383_),
    .QN(_00932_));
 DFFHQNx1_ASAP7_75t_R \u0.w[2][9]$_DFF_P_  (.CLK(clknet_leaf_11_clk),
    .D(_00384_),
    .QN(_00933_));
 DFFHQNx1_ASAP7_75t_R \u0.w[3][0]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .D(net6296),
    .QN(_00934_));
 DFFHQNx1_ASAP7_75t_R \u0.w[3][10]$_DFF_P_  (.CLK(clknet_leaf_2_clk),
    .D(_08962_),
    .QN(_00935_));
 DFFHQNx1_ASAP7_75t_R \u0.w[3][11]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .D(net5945),
    .QN(_00936_));
 DFFHQNx1_ASAP7_75t_R \u0.w[3][12]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .D(net6304),
    .QN(_00937_));
 DFFHQNx1_ASAP7_75t_R \u0.w[3][13]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .D(net6303),
    .QN(_00938_));
 DFFHQNx1_ASAP7_75t_R \u0.w[3][14]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .D(net5943),
    .QN(_00939_));
 DFFHQNx1_ASAP7_75t_R \u0.w[3][15]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .D(net5942),
    .QN(_00940_));
 DFFHQNx1_ASAP7_75t_R \u0.w[3][16]$_DFF_P_  (.CLK(clknet_leaf_30_clk),
    .D(net5981),
    .QN(_00941_));
 DFFHQNx1_ASAP7_75t_R \u0.w[3][17]$_DFF_P_  (.CLK(clknet_leaf_30_clk),
    .D(net5983),
    .QN(_00942_));
 DFFHQNx1_ASAP7_75t_R \u0.w[3][18]$_DFF_P_  (.CLK(clknet_leaf_30_clk),
    .D(net6338),
    .QN(_00943_));
 DFFHQNx1_ASAP7_75t_R \u0.w[3][19]$_DFF_P_  (.CLK(clknet_leaf_30_clk),
    .D(net6374),
    .QN(_00944_));
 DFFHQNx1_ASAP7_75t_R \u0.w[3][1]$_DFF_P_  (.CLK(clknet_leaf_2_clk),
    .D(net6323),
    .QN(_00945_));
 DFFHQNx1_ASAP7_75t_R \u0.w[3][20]$_DFF_P_  (.CLK(clknet_leaf_30_clk),
    .D(net6336),
    .QN(_00946_));
 DFFHQNx1_ASAP7_75t_R \u0.w[3][21]$_DFF_P_  (.CLK(clknet_leaf_31_clk),
    .D(net6333),
    .QN(_00947_));
 DFFHQNx1_ASAP7_75t_R \u0.w[3][22]$_DFF_P_  (.CLK(clknet_leaf_27_clk),
    .D(net6332),
    .QN(_00948_));
 DFFHQNx1_ASAP7_75t_R \u0.w[3][23]$_DFF_P_  (.CLK(clknet_leaf_27_clk),
    .D(_08097_),
    .QN(_00949_));
 DFFHQNx1_ASAP7_75t_R \u0.w[3][24]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .D(net6287),
    .QN(_00950_));
 DFFHQNx1_ASAP7_75t_R \u0.w[3][25]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .D(net6299),
    .QN(_00951_));
 DFFHQNx1_ASAP7_75t_R \u0.w[3][26]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .D(net6289),
    .QN(_00952_));
 DFFHQNx1_ASAP7_75t_R \u0.w[3][27]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .D(net5934),
    .QN(_00953_));
 DFFHQNx1_ASAP7_75t_R \u0.w[3][28]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .D(net6297),
    .QN(_00954_));
 DFFHQNx1_ASAP7_75t_R \u0.w[3][29]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .D(net5558),
    .QN(_00955_));
 DFFHQNx1_ASAP7_75t_R \u0.w[3][2]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .D(net5963),
    .QN(_00956_));
 DFFHQNx1_ASAP7_75t_R \u0.w[3][30]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .D(net5932),
    .QN(_00957_));
 DFFHQNx1_ASAP7_75t_R \u0.w[3][31]$_DFF_P_  (.CLK(clknet_leaf_34_clk),
    .D(net5557),
    .QN(_00958_));
 DFFHQNx1_ASAP7_75t_R \u0.w[3][3]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .D(net5961),
    .QN(_00959_));
 DFFHQNx1_ASAP7_75t_R \u0.w[3][4]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .D(net6318),
    .QN(_00960_));
 DFFHQNx1_ASAP7_75t_R \u0.w[3][5]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .D(net6313),
    .QN(_00961_));
 DFFHQNx1_ASAP7_75t_R \u0.w[3][6]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .D(net5954),
    .QN(_00962_));
 DFFHQNx1_ASAP7_75t_R \u0.w[3][7]$_DFF_P_  (.CLK(clknet_leaf_2_clk),
    .D(net5953),
    .QN(_00963_));
 DFFHQNx1_ASAP7_75t_R \u0.w[3][8]$_DFF_P_  (.CLK(clknet_leaf_2_clk),
    .D(net6311),
    .QN(_00964_));
 DFFHQNx1_ASAP7_75t_R \u0.w[3][9]$_DFF_P_  (.CLK(clknet_leaf_2_clk),
    .D(net5931),
    .QN(_00486_));
endmodule
